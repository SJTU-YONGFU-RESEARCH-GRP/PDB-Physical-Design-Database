module dynamic_node_top_wrap (clk,
    reset_in,
    thanksIn_P,
    validIn_E,
    validIn_N,
    validIn_P,
    validIn_S,
    validIn_W,
    validOut_E,
    validOut_N,
    validOut_P,
    validOut_S,
    validOut_W,
    yummyIn_E,
    yummyIn_N,
    yummyIn_P,
    yummyIn_S,
    yummyIn_W,
    yummyOut_E,
    yummyOut_N,
    yummyOut_P,
    yummyOut_S,
    yummyOut_W,
    dataIn_E,
    dataIn_N,
    dataIn_P,
    dataIn_S,
    dataIn_W,
    dataOut_E,
    dataOut_N,
    dataOut_P,
    dataOut_S,
    dataOut_W,
    myChipID,
    myLocX,
    myLocY);
 input clk;
 input reset_in;
 output thanksIn_P;
 input validIn_E;
 input validIn_N;
 input validIn_P;
 input validIn_S;
 input validIn_W;
 output validOut_E;
 output validOut_N;
 output validOut_P;
 output validOut_S;
 output validOut_W;
 input yummyIn_E;
 input yummyIn_N;
 input yummyIn_P;
 input yummyIn_S;
 input yummyIn_W;
 output yummyOut_E;
 output yummyOut_N;
 output yummyOut_P;
 output yummyOut_S;
 output yummyOut_W;
 input [63:0] dataIn_E;
 input [63:0] dataIn_N;
 input [63:0] dataIn_P;
 input [63:0] dataIn_S;
 input [63:0] dataIn_W;
 output [63:0] dataOut_E;
 output [63:0] dataOut_N;
 output [63:0] dataOut_P;
 output [63:0] dataOut_S;
 output [63:0] dataOut_W;
 input [13:0] myChipID;
 input [7:0] myLocX;
 input [7:0] myLocY;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire net2;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire net4;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire net6;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire net1;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire net752;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire net7;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire net3;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire net770;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire net756;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire net760;
 wire _05699_;
 wire _05700_;
 wire net761;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire net691;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire net5;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire \dynamic_node_top.REG_reset_fin.q ;
 wire \dynamic_node_top.east_input.NIB.elements_in_array_f[0] ;
 wire \dynamic_node_top.east_input.NIB.elements_in_array_f[1] ;
 wire \dynamic_node_top.east_input.NIB.elements_in_array_f[2] ;
 wire \dynamic_node_top.east_input.NIB.elements_in_array_next[0] ;
 wire \dynamic_node_top.east_input.NIB.head_ptr_f[0] ;
 wire \dynamic_node_top.east_input.NIB.head_ptr_f[1] ;
 wire \dynamic_node_top.east_input.NIB.head_ptr_next[0] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][0] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][10] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][11] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][12] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][13] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][14] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][15] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][16] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][17] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][18] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][19] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][1] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][20] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][21] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][22] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][23] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][24] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][25] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][26] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][27] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][28] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][29] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][2] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][30] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][31] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][32] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][33] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][34] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][35] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][36] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][37] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][38] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][39] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][3] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][40] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][41] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][42] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][43] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][44] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][45] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][46] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][47] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][48] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][49] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][4] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][50] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][51] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][52] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][53] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][54] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][55] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][56] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][57] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][58] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][59] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][5] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][60] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][61] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][62] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][63] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][6] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][7] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][8] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[0][9] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][0] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][10] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][11] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][12] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][13] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][14] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][15] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][16] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][17] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][18] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][19] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][1] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][20] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][21] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][22] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][23] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][24] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][25] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][26] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][27] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][28] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][29] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][2] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][30] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][31] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][32] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][33] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][34] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][35] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][36] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][37] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][38] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][39] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][3] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][40] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][41] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][42] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][43] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][44] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][45] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][46] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][47] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][48] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][49] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][4] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][50] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][51] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][52] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][53] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][54] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][55] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][56] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][57] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][58] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][59] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][5] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][60] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][61] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][62] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][63] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][6] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][7] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][8] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[1][9] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][0] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][10] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][11] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][12] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][13] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][14] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][15] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][16] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][17] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][18] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][19] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][1] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][20] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][21] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][22] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][23] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][24] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][25] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][26] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][27] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][28] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][29] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][2] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][30] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][31] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][32] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][33] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][34] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][35] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][36] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][37] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][38] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][39] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][3] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][40] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][41] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][42] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][43] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][44] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][45] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][46] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][47] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][48] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][49] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][4] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][50] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][51] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][52] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][53] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][54] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][55] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][56] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][57] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][58] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][59] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][5] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][60] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][61] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][62] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][63] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][6] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][7] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][8] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[2][9] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][0] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][10] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][11] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][12] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][13] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][14] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][15] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][16] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][17] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][18] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][19] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][1] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][20] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][21] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][22] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][23] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][24] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][25] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][26] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][27] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][28] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][29] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][2] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][30] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][31] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][32] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][33] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][34] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][35] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][36] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][37] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][38] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][39] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][3] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][40] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][41] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][42] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][43] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][44] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][45] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][46] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][47] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][48] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][49] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][4] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][50] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][51] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][52] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][53] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][54] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][55] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][56] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][57] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][58] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][59] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][5] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][60] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][61] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][62] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][63] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][6] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][7] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][8] ;
 wire \dynamic_node_top.east_input.NIB.storage_data_f[3][9] ;
 wire \dynamic_node_top.east_input.NIB.tail_ptr_f[0] ;
 wire \dynamic_node_top.east_input.NIB.tail_ptr_f[1] ;
 wire \dynamic_node_top.east_input.NIB.tail_ptr_next[0] ;
 wire \dynamic_node_top.east_input.NIB.tail_ptr_next[1] ;
 wire \dynamic_node_top.east_input.NIB.thanks_in ;
 wire \dynamic_node_top.east_input.control.count_f[0] ;
 wire \dynamic_node_top.east_input.control.count_f[1] ;
 wire \dynamic_node_top.east_input.control.count_f[2] ;
 wire \dynamic_node_top.east_input.control.count_f[3] ;
 wire \dynamic_node_top.east_input.control.count_f[4] ;
 wire \dynamic_node_top.east_input.control.count_f[5] ;
 wire \dynamic_node_top.east_input.control.count_f[6] ;
 wire \dynamic_node_top.east_input.control.count_f[7] ;
 wire \dynamic_node_top.east_input.control.count_one_f ;
 wire \dynamic_node_top.east_input.control.header_last_temp ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[0] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[10] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[11] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[12] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[13] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[1] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[2] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[3] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[4] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[5] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[6] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[7] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[8] ;
 wire \dynamic_node_top.east_input.control.my_chip_id_in[9] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[0] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[1] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[2] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[3] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[4] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[5] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[6] ;
 wire \dynamic_node_top.east_input.control.my_loc_x_in[7] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[0] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[1] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[2] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[3] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[4] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[5] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[6] ;
 wire \dynamic_node_top.east_input.control.my_loc_y_in[7] ;
 wire \dynamic_node_top.east_input.control.tail_last_f ;
 wire \dynamic_node_top.east_output.control.current_route_f[0] ;
 wire \dynamic_node_top.east_output.control.current_route_f[1] ;
 wire \dynamic_node_top.east_output.control.current_route_f[2] ;
 wire \dynamic_node_top.east_output.control.current_route_f[3] ;
 wire \dynamic_node_top.east_output.control.current_route_f[4] ;
 wire \dynamic_node_top.east_output.control.planned_f ;
 wire \dynamic_node_top.east_output.space.count_f[0] ;
 wire \dynamic_node_top.east_output.space.count_f[1] ;
 wire \dynamic_node_top.east_output.space.count_f[2] ;
 wire \dynamic_node_top.east_output.space.is_one_f ;
 wire \dynamic_node_top.east_output.space.is_two_or_more_f ;
 wire \dynamic_node_top.east_output.space.valid_f ;
 wire \dynamic_node_top.east_output.space.yummy_f ;
 wire \dynamic_node_top.north_input.NIB.elements_in_array_f[0] ;
 wire \dynamic_node_top.north_input.NIB.elements_in_array_f[1] ;
 wire \dynamic_node_top.north_input.NIB.elements_in_array_f[2] ;
 wire \dynamic_node_top.north_input.NIB.elements_in_array_next[0] ;
 wire \dynamic_node_top.north_input.NIB.head_ptr_f[0] ;
 wire \dynamic_node_top.north_input.NIB.head_ptr_f[1] ;
 wire \dynamic_node_top.north_input.NIB.head_ptr_next[0] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][0] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][10] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][11] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][12] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][13] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][14] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][15] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][16] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][17] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][18] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][19] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][1] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][20] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][21] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][22] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][23] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][24] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][25] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][26] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][27] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][28] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][29] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][2] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][30] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][31] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][32] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][33] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][34] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][35] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][36] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][37] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][38] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][39] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][3] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][40] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][41] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][42] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][43] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][44] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][45] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][46] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][47] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][48] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][49] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][4] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][50] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][51] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][52] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][53] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][54] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][55] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][56] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][57] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][58] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][59] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][5] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][60] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][61] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][62] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][63] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][6] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][7] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][8] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[0][9] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][0] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][10] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][11] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][12] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][13] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][14] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][15] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][16] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][17] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][18] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][19] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][1] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][20] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][21] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][22] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][23] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][24] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][25] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][26] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][27] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][28] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][29] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][2] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][30] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][31] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][32] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][33] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][34] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][35] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][36] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][37] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][38] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][39] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][3] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][40] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][41] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][42] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][43] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][44] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][45] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][46] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][47] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][48] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][49] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][4] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][50] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][51] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][52] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][53] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][54] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][55] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][56] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][57] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][58] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][59] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][5] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][60] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][61] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][62] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][63] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][6] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][7] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][8] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[1][9] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][0] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][10] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][11] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][12] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][13] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][14] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][15] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][16] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][17] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][18] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][19] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][1] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][20] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][21] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][22] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][23] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][24] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][25] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][26] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][27] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][28] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][29] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][2] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][30] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][31] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][32] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][33] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][34] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][35] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][36] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][37] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][38] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][39] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][3] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][40] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][41] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][42] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][43] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][44] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][45] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][46] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][47] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][48] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][49] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][4] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][50] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][51] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][52] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][53] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][54] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][55] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][56] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][57] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][58] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][59] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][5] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][60] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][61] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][62] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][63] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][6] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][7] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][8] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[2][9] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][0] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][10] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][11] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][12] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][13] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][14] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][15] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][16] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][17] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][18] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][19] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][1] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][20] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][21] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][22] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][23] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][24] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][25] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][26] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][27] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][28] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][29] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][2] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][30] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][31] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][32] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][33] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][34] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][35] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][36] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][37] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][38] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][39] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][3] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][40] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][41] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][42] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][43] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][44] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][45] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][46] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][47] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][48] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][49] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][4] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][50] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][51] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][52] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][53] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][54] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][55] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][56] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][57] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][58] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][59] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][5] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][60] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][61] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][62] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][63] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][6] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][7] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][8] ;
 wire \dynamic_node_top.north_input.NIB.storage_data_f[3][9] ;
 wire \dynamic_node_top.north_input.NIB.tail_ptr_f[0] ;
 wire \dynamic_node_top.north_input.NIB.tail_ptr_f[1] ;
 wire \dynamic_node_top.north_input.NIB.tail_ptr_next[0] ;
 wire \dynamic_node_top.north_input.NIB.tail_ptr_next[1] ;
 wire \dynamic_node_top.north_input.NIB.thanks_in ;
 wire \dynamic_node_top.north_input.control.count_f[0] ;
 wire \dynamic_node_top.north_input.control.count_f[1] ;
 wire \dynamic_node_top.north_input.control.count_f[2] ;
 wire \dynamic_node_top.north_input.control.count_f[3] ;
 wire \dynamic_node_top.north_input.control.count_f[4] ;
 wire \dynamic_node_top.north_input.control.count_f[5] ;
 wire \dynamic_node_top.north_input.control.count_f[6] ;
 wire \dynamic_node_top.north_input.control.count_f[7] ;
 wire \dynamic_node_top.north_input.control.count_one_f ;
 wire \dynamic_node_top.north_input.control.header_last_temp ;
 wire \dynamic_node_top.north_input.control.tail_last_f ;
 wire \dynamic_node_top.north_output.control.current_route_f[0] ;
 wire \dynamic_node_top.north_output.control.current_route_f[1] ;
 wire \dynamic_node_top.north_output.control.current_route_f[2] ;
 wire \dynamic_node_top.north_output.control.current_route_f[3] ;
 wire \dynamic_node_top.north_output.control.current_route_f[4] ;
 wire \dynamic_node_top.north_output.control.planned_f ;
 wire \dynamic_node_top.north_output.space.count_f[0] ;
 wire \dynamic_node_top.north_output.space.count_f[1] ;
 wire \dynamic_node_top.north_output.space.count_f[2] ;
 wire \dynamic_node_top.north_output.space.is_one_f ;
 wire \dynamic_node_top.north_output.space.is_two_or_more_f ;
 wire \dynamic_node_top.north_output.space.valid_f ;
 wire \dynamic_node_top.north_output.space.yummy_f ;
 wire \dynamic_node_top.proc_input.NIB.elements_in_array_f[0] ;
 wire \dynamic_node_top.proc_input.NIB.elements_in_array_f[1] ;
 wire \dynamic_node_top.proc_input.NIB.elements_in_array_f[2] ;
 wire \dynamic_node_top.proc_input.NIB.elements_in_array_f[3] ;
 wire \dynamic_node_top.proc_input.NIB.elements_in_array_f[4] ;
 wire \dynamic_node_top.proc_input.NIB.elements_in_array_next[0] ;
 wire \dynamic_node_top.proc_input.NIB.head_ptr_f[0] ;
 wire \dynamic_node_top.proc_input.NIB.head_ptr_f[1] ;
 wire \dynamic_node_top.proc_input.NIB.head_ptr_f[2] ;
 wire \dynamic_node_top.proc_input.NIB.head_ptr_f[3] ;
 wire \dynamic_node_top.proc_input.NIB.head_ptr_next[0] ;
 wire \dynamic_node_top.proc_input.NIB.head_ptr_next[1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[0][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[10][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[11][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[12][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[13][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[14][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[15][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[1][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[2][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[3][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[4][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[5][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[6][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[7][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[8][9] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][0] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][10] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][11] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][12] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][13] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][14] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][15] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][16] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][17] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][18] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][19] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][1] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][20] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][21] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][22] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][23] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][24] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][25] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][26] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][27] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][28] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][29] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][2] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][30] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][31] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][32] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][33] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][34] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][35] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][36] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][37] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][38] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][39] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][3] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][40] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][41] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][42] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][43] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][44] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][45] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][46] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][47] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][48] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][49] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][4] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][50] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][51] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][52] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][53] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][54] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][55] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][56] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][57] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][58] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][59] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][5] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][60] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][61] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][62] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][63] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][6] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][7] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][8] ;
 wire \dynamic_node_top.proc_input.NIB.storage_data_f[9][9] ;
 wire \dynamic_node_top.proc_input.NIB.tail_ptr_f[0] ;
 wire \dynamic_node_top.proc_input.NIB.tail_ptr_f[1] ;
 wire \dynamic_node_top.proc_input.NIB.tail_ptr_f[2] ;
 wire \dynamic_node_top.proc_input.NIB.tail_ptr_f[3] ;
 wire \dynamic_node_top.proc_input.NIB.tail_ptr_next[0] ;
 wire \dynamic_node_top.proc_input.NIB.tail_ptr_next[1] ;
 wire \dynamic_node_top.proc_input.control.count_f[0] ;
 wire \dynamic_node_top.proc_input.control.count_f[1] ;
 wire \dynamic_node_top.proc_input.control.count_f[2] ;
 wire \dynamic_node_top.proc_input.control.count_f[3] ;
 wire \dynamic_node_top.proc_input.control.count_f[4] ;
 wire \dynamic_node_top.proc_input.control.count_f[5] ;
 wire \dynamic_node_top.proc_input.control.count_f[6] ;
 wire \dynamic_node_top.proc_input.control.count_f[7] ;
 wire \dynamic_node_top.proc_input.control.count_one_f ;
 wire \dynamic_node_top.proc_input.control.header_last_temp ;
 wire \dynamic_node_top.proc_input.control.tail_last_f ;
 wire \dynamic_node_top.proc_output.control.current_route_f[0] ;
 wire \dynamic_node_top.proc_output.control.current_route_f[1] ;
 wire \dynamic_node_top.proc_output.control.current_route_f[2] ;
 wire \dynamic_node_top.proc_output.control.current_route_f[3] ;
 wire \dynamic_node_top.proc_output.control.current_route_f[4] ;
 wire \dynamic_node_top.proc_output.control.planned_f ;
 wire \dynamic_node_top.proc_output.space.count_f[0] ;
 wire \dynamic_node_top.proc_output.space.count_f[1] ;
 wire \dynamic_node_top.proc_output.space.count_f[2] ;
 wire \dynamic_node_top.proc_output.space.is_one_f ;
 wire \dynamic_node_top.proc_output.space.is_two_or_more_f ;
 wire \dynamic_node_top.proc_output.space.valid_f ;
 wire \dynamic_node_top.proc_output.space.yummy_f ;
 wire \dynamic_node_top.south_input.NIB.elements_in_array_f[0] ;
 wire \dynamic_node_top.south_input.NIB.elements_in_array_f[1] ;
 wire \dynamic_node_top.south_input.NIB.elements_in_array_f[2] ;
 wire \dynamic_node_top.south_input.NIB.elements_in_array_next[0] ;
 wire \dynamic_node_top.south_input.NIB.head_ptr_f[0] ;
 wire \dynamic_node_top.south_input.NIB.head_ptr_f[1] ;
 wire \dynamic_node_top.south_input.NIB.head_ptr_next[0] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][0] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][10] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][11] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][12] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][13] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][14] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][15] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][16] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][17] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][18] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][19] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][1] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][20] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][21] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][22] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][23] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][24] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][25] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][26] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][27] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][28] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][29] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][2] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][30] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][31] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][32] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][33] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][34] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][35] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][36] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][37] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][38] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][39] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][3] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][40] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][41] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][42] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][43] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][44] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][45] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][46] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][47] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][48] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][49] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][4] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][50] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][51] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][52] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][53] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][54] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][55] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][56] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][57] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][58] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][59] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][5] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][60] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][61] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][62] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][63] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][6] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][7] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][8] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[0][9] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][0] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][10] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][11] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][12] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][13] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][14] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][15] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][16] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][17] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][18] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][19] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][1] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][20] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][21] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][22] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][23] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][24] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][25] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][26] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][27] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][28] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][29] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][2] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][30] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][31] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][32] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][33] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][34] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][35] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][36] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][37] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][38] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][39] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][3] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][40] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][41] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][42] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][43] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][44] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][45] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][46] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][47] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][48] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][49] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][4] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][50] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][51] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][52] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][53] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][54] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][55] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][56] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][57] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][58] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][59] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][5] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][60] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][61] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][62] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][63] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][6] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][7] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][8] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[1][9] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][0] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][10] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][11] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][12] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][13] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][14] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][15] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][16] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][17] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][18] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][19] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][1] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][20] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][21] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][22] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][23] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][24] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][25] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][26] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][27] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][28] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][29] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][2] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][30] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][31] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][32] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][33] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][34] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][35] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][36] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][37] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][38] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][39] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][3] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][40] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][41] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][42] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][43] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][44] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][45] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][46] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][47] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][48] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][49] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][4] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][50] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][51] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][52] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][53] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][54] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][55] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][56] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][57] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][58] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][59] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][5] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][60] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][61] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][62] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][63] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][6] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][7] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][8] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[2][9] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][0] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][10] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][11] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][12] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][13] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][14] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][15] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][16] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][17] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][18] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][19] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][1] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][20] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][21] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][22] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][23] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][24] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][25] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][26] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][27] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][28] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][29] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][2] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][30] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][31] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][32] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][33] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][34] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][35] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][36] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][37] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][38] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][39] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][3] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][40] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][41] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][42] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][43] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][44] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][45] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][46] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][47] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][48] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][49] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][4] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][50] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][51] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][52] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][53] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][54] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][55] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][56] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][57] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][58] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][59] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][5] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][60] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][61] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][62] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][63] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][6] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][7] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][8] ;
 wire \dynamic_node_top.south_input.NIB.storage_data_f[3][9] ;
 wire \dynamic_node_top.south_input.NIB.tail_ptr_f[0] ;
 wire \dynamic_node_top.south_input.NIB.tail_ptr_f[1] ;
 wire \dynamic_node_top.south_input.NIB.tail_ptr_next[0] ;
 wire \dynamic_node_top.south_input.NIB.tail_ptr_next[1] ;
 wire \dynamic_node_top.south_input.NIB.thanks_in ;
 wire \dynamic_node_top.south_input.control.count_f[0] ;
 wire \dynamic_node_top.south_input.control.count_f[1] ;
 wire \dynamic_node_top.south_input.control.count_f[2] ;
 wire \dynamic_node_top.south_input.control.count_f[3] ;
 wire \dynamic_node_top.south_input.control.count_f[4] ;
 wire \dynamic_node_top.south_input.control.count_f[5] ;
 wire \dynamic_node_top.south_input.control.count_f[6] ;
 wire \dynamic_node_top.south_input.control.count_f[7] ;
 wire \dynamic_node_top.south_input.control.count_one_f ;
 wire \dynamic_node_top.south_input.control.header_last_temp ;
 wire \dynamic_node_top.south_input.control.tail_last_f ;
 wire \dynamic_node_top.south_output.control.current_route_f[0] ;
 wire \dynamic_node_top.south_output.control.current_route_f[1] ;
 wire \dynamic_node_top.south_output.control.current_route_f[2] ;
 wire \dynamic_node_top.south_output.control.current_route_f[3] ;
 wire \dynamic_node_top.south_output.control.current_route_f[4] ;
 wire \dynamic_node_top.south_output.control.planned_f ;
 wire \dynamic_node_top.south_output.space.count_f[0] ;
 wire \dynamic_node_top.south_output.space.count_f[1] ;
 wire \dynamic_node_top.south_output.space.count_f[2] ;
 wire \dynamic_node_top.south_output.space.is_one_f ;
 wire \dynamic_node_top.south_output.space.is_two_or_more_f ;
 wire \dynamic_node_top.south_output.space.valid_f ;
 wire \dynamic_node_top.south_output.space.yummy_f ;
 wire \dynamic_node_top.west_input.NIB.elements_in_array_f[0] ;
 wire \dynamic_node_top.west_input.NIB.elements_in_array_f[1] ;
 wire \dynamic_node_top.west_input.NIB.elements_in_array_f[2] ;
 wire \dynamic_node_top.west_input.NIB.elements_in_array_next[0] ;
 wire \dynamic_node_top.west_input.NIB.head_ptr_f[0] ;
 wire \dynamic_node_top.west_input.NIB.head_ptr_f[1] ;
 wire \dynamic_node_top.west_input.NIB.head_ptr_next[0] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][0] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][10] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][11] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][12] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][13] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][14] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][15] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][16] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][17] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][18] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][19] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][1] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][20] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][21] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][22] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][23] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][24] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][25] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][26] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][27] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][28] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][29] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][2] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][30] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][31] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][32] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][33] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][34] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][35] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][36] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][37] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][38] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][39] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][3] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][40] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][41] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][42] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][43] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][44] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][45] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][46] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][47] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][48] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][49] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][4] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][50] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][51] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][52] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][53] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][54] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][55] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][56] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][57] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][58] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][59] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][5] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][60] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][61] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][62] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][63] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][6] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][7] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][8] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[0][9] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][0] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][10] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][11] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][12] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][13] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][14] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][15] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][16] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][17] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][18] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][19] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][1] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][20] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][21] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][22] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][23] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][24] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][25] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][26] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][27] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][28] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][29] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][2] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][30] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][31] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][32] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][33] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][34] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][35] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][36] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][37] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][38] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][39] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][3] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][40] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][41] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][42] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][43] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][44] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][45] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][46] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][47] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][48] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][49] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][4] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][50] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][51] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][52] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][53] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][54] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][55] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][56] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][57] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][58] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][59] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][5] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][60] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][61] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][62] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][63] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][6] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][7] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][8] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[1][9] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][0] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][10] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][11] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][12] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][13] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][14] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][15] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][16] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][17] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][18] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][19] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][1] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][20] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][21] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][22] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][23] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][24] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][25] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][26] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][27] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][28] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][29] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][2] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][30] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][31] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][32] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][33] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][34] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][35] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][36] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][37] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][38] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][39] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][3] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][40] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][41] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][42] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][43] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][44] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][45] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][46] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][47] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][48] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][49] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][4] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][50] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][51] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][52] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][53] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][54] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][55] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][56] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][57] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][58] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][59] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][5] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][60] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][61] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][62] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][63] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][6] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][7] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][8] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[2][9] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][0] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][10] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][11] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][12] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][13] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][14] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][15] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][16] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][17] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][18] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][19] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][1] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][20] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][21] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][22] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][23] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][24] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][25] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][26] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][27] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][28] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][29] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][2] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][30] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][31] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][32] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][33] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][34] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][35] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][36] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][37] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][38] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][39] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][3] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][40] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][41] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][42] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][43] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][44] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][45] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][46] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][47] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][48] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][49] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][4] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][50] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][51] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][52] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][53] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][54] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][55] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][56] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][57] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][58] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][59] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][5] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][60] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][61] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][62] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][63] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][6] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][7] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][8] ;
 wire \dynamic_node_top.west_input.NIB.storage_data_f[3][9] ;
 wire \dynamic_node_top.west_input.NIB.tail_ptr_f[0] ;
 wire \dynamic_node_top.west_input.NIB.tail_ptr_f[1] ;
 wire \dynamic_node_top.west_input.NIB.tail_ptr_next[0] ;
 wire \dynamic_node_top.west_input.NIB.tail_ptr_next[1] ;
 wire \dynamic_node_top.west_input.NIB.thanks_in ;
 wire \dynamic_node_top.west_input.control.count_f[0] ;
 wire \dynamic_node_top.west_input.control.count_f[1] ;
 wire \dynamic_node_top.west_input.control.count_f[2] ;
 wire \dynamic_node_top.west_input.control.count_f[3] ;
 wire \dynamic_node_top.west_input.control.count_f[4] ;
 wire \dynamic_node_top.west_input.control.count_f[5] ;
 wire \dynamic_node_top.west_input.control.count_f[6] ;
 wire \dynamic_node_top.west_input.control.count_f[7] ;
 wire \dynamic_node_top.west_input.control.count_one_f ;
 wire \dynamic_node_top.west_input.control.header_last_temp ;
 wire \dynamic_node_top.west_input.control.tail_last_f ;
 wire \dynamic_node_top.west_output.control.current_route_f[0] ;
 wire \dynamic_node_top.west_output.control.current_route_f[1] ;
 wire \dynamic_node_top.west_output.control.current_route_f[2] ;
 wire \dynamic_node_top.west_output.control.current_route_f[3] ;
 wire \dynamic_node_top.west_output.control.current_route_f[4] ;
 wire \dynamic_node_top.west_output.control.planned_f ;
 wire \dynamic_node_top.west_output.space.count_f[0] ;
 wire \dynamic_node_top.west_output.space.count_f[1] ;
 wire \dynamic_node_top.west_output.space.count_f[2] ;
 wire \dynamic_node_top.west_output.space.is_one_f ;
 wire \dynamic_node_top.west_output.space.is_two_or_more_f ;
 wire \dynamic_node_top.west_output.space.valid_f ;
 wire \dynamic_node_top.west_output.space.yummy_f ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net758;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net765;
 wire net764;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net744;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net742;
 wire net743;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net753;
 wire net754;
 wire net757;
 wire net771;

 BUF_X8 _10617_ (.A(_00013_),
    .Z(_05124_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 BUF_X4 _10619_ (.A(_05124_),
    .Z(_05126_));
 BUF_X8 _10620_ (.A(_05126_),
    .Z(_05127_));
 BUF_X8 _10621_ (.A(_00014_),
    .Z(_05128_));
 BUF_X16 _10622_ (.A(_05128_),
    .Z(_05129_));
 BUF_X32 _10623_ (.A(_05129_),
    .Z(_05130_));
 BUF_X2 clone2 (.A(net658),
    .Z(net2));
 BUF_X32 _10625_ (.A(_05130_),
    .Z(_05132_));
 MUX2_X1 _10626_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][42] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][42] ),
    .S(_05132_),
    .Z(_05133_));
 INV_X1 _10627_ (.A(_05133_),
    .ZN(_05134_));
 NAND2_X1 _10628_ (.A1(_05127_),
    .A2(_05134_),
    .ZN(_05135_));
 BUF_X32 _10629_ (.A(_05130_),
    .Z(_05136_));
 MUX2_X1 _10630_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][42] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][42] ),
    .S(net745),
    .Z(_05137_));
 OAI21_X4 _10631_ (.A(_05135_),
    .B1(_05137_),
    .B2(_05127_),
    .ZN(_05138_));
 INV_X1 _10632_ (.A(_05138_),
    .ZN(_10179_));
 MUX2_X1 _10633_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][34] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][34] ),
    .S(net745),
    .Z(_05139_));
 MUX2_X1 _10634_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][34] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][34] ),
    .S(net745),
    .Z(_05140_));
 MUX2_X2 _10635_ (.A(_05139_),
    .B(_05140_),
    .S(_05126_),
    .Z(_10225_));
 BUF_X8 _10636_ (.A(_00016_),
    .Z(_05141_));
 BUF_X16 _10637_ (.A(_05141_),
    .Z(_05142_));
 BUF_X32 _10638_ (.A(_05142_),
    .Z(_05143_));
 BUF_X32 _10639_ (.A(_05143_),
    .Z(_05144_));
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 BUF_X32 _10641_ (.A(_05144_),
    .Z(_05146_));
 BUF_X32 _10642_ (.A(_05146_),
    .Z(_05147_));
 MUX2_X1 _10643_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][42] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][42] ),
    .S(_05147_),
    .Z(_05148_));
 MUX2_X1 _10644_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][42] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][42] ),
    .S(_05147_),
    .Z(_05149_));
 CLKBUF_X3 _10645_ (.A(_00015_),
    .Z(_05150_));
 BUF_X4 _10646_ (.A(_05150_),
    .Z(_05151_));
 CLKBUF_X3 _10647_ (.A(_05151_),
    .Z(_05152_));
 BUF_X4 _10648_ (.A(_05152_),
    .Z(_05153_));
 MUX2_X2 _10649_ (.A(_05148_),
    .B(_05149_),
    .S(_05153_),
    .Z(_10249_));
 MUX2_X1 _10650_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][34] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][34] ),
    .S(net739),
    .Z(_05154_));
 MUX2_X1 _10651_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][34] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][34] ),
    .S(net739),
    .Z(_05155_));
 MUX2_X2 _10652_ (.A(_05154_),
    .B(_05155_),
    .S(_05152_),
    .Z(_10252_));
 BUF_X4 _10653_ (.A(_00045_),
    .Z(_05156_));
 INV_X2 _10654_ (.A(_05156_),
    .ZN(_05157_));
 CLKBUF_X3 _10655_ (.A(\dynamic_node_top.east_output.control.current_route_f[3] ),
    .Z(_05158_));
 CLKBUF_X3 _10656_ (.A(\dynamic_node_top.east_output.control.current_route_f[1] ),
    .Z(_05159_));
 NOR4_X4 _10657_ (.A1(\dynamic_node_top.east_output.control.current_route_f[4] ),
    .A2(\dynamic_node_top.east_output.control.current_route_f[2] ),
    .A3(_05158_),
    .A4(_05159_),
    .ZN(_05160_));
 INV_X1 _10658_ (.A(_05160_),
    .ZN(_05161_));
 NOR2_X1 _10659_ (.A1(_05157_),
    .A2(_05161_),
    .ZN(_05162_));
 BUF_X8 _10660_ (.A(_05162_),
    .Z(_05163_));
 INV_X1 _10661_ (.A(\dynamic_node_top.east_output.space.is_one_f ),
    .ZN(_05164_));
 NOR2_X1 _10662_ (.A1(_05164_),
    .A2(\dynamic_node_top.east_output.space.valid_f ),
    .ZN(_05165_));
 NOR3_X2 _10663_ (.A1(\dynamic_node_top.east_output.space.is_two_or_more_f ),
    .A2(\dynamic_node_top.east_output.space.yummy_f ),
    .A3(_05165_),
    .ZN(_05166_));
 CLKBUF_X3 _10664_ (.A(\dynamic_node_top.east_output.control.current_route_f[2] ),
    .Z(_05167_));
 OR3_X4 _10665_ (.A1(\dynamic_node_top.north_input.NIB.elements_in_array_f[1] ),
    .A2(\dynamic_node_top.north_input.NIB.elements_in_array_f[0] ),
    .A3(\dynamic_node_top.north_input.NIB.elements_in_array_f[2] ),
    .ZN(_05168_));
 OR3_X1 _10666_ (.A1(\dynamic_node_top.south_input.NIB.elements_in_array_f[1] ),
    .A2(\dynamic_node_top.south_input.NIB.elements_in_array_f[0] ),
    .A3(\dynamic_node_top.south_input.NIB.elements_in_array_f[2] ),
    .ZN(_05169_));
 CLKBUF_X3 _10667_ (.A(_05169_),
    .Z(_05170_));
 CLKBUF_X3 _10668_ (.A(\dynamic_node_top.east_output.control.current_route_f[4] ),
    .Z(_05171_));
 AOI22_X1 _10669_ (.A1(_05167_),
    .A2(_05168_),
    .B1(_05170_),
    .B2(_05171_),
    .ZN(_05172_));
 BUF_X2 _10670_ (.A(\dynamic_node_top.east_output.control.current_route_f[0] ),
    .Z(_05173_));
 OR3_X1 _10671_ (.A1(\dynamic_node_top.west_input.NIB.elements_in_array_f[1] ),
    .A2(\dynamic_node_top.west_input.NIB.elements_in_array_f[0] ),
    .A3(\dynamic_node_top.west_input.NIB.elements_in_array_f[2] ),
    .ZN(_05174_));
 CLKBUF_X3 _10672_ (.A(_05174_),
    .Z(_05175_));
 OR3_X1 _10673_ (.A1(\dynamic_node_top.east_input.NIB.elements_in_array_f[1] ),
    .A2(\dynamic_node_top.east_input.NIB.elements_in_array_f[0] ),
    .A3(\dynamic_node_top.east_input.NIB.elements_in_array_f[2] ),
    .ZN(_05176_));
 BUF_X4 _10674_ (.A(_05176_),
    .Z(_05177_));
 INV_X1 _10675_ (.A(_00044_),
    .ZN(_05178_));
 AOI22_X1 _10676_ (.A1(_05173_),
    .A2(_05175_),
    .B1(_05177_),
    .B2(_05178_),
    .ZN(_05179_));
 NAND2_X1 _10677_ (.A1(_05172_),
    .A2(_05179_),
    .ZN(_05180_));
 OR4_X2 _10678_ (.A1(\dynamic_node_top.proc_input.NIB.elements_in_array_f[0] ),
    .A2(\dynamic_node_top.proc_input.NIB.elements_in_array_f[3] ),
    .A3(\dynamic_node_top.proc_input.NIB.elements_in_array_f[2] ),
    .A4(\dynamic_node_top.proc_input.NIB.elements_in_array_f[4] ),
    .ZN(_05181_));
 OR2_X4 _10679_ (.A1(\dynamic_node_top.proc_input.NIB.elements_in_array_f[1] ),
    .A2(_05181_),
    .ZN(_05182_));
 AOI21_X2 _10680_ (.A(_05180_),
    .B1(_05182_),
    .B2(_05158_),
    .ZN(_05183_));
 NOR3_X4 _10681_ (.A1(_05163_),
    .A2(_05166_),
    .A3(_05183_),
    .ZN(_05184_));
 NAND2_X4 _10682_ (.A1(\dynamic_node_top.west_input.control.header_last_temp ),
    .A2(_05175_),
    .ZN(_05185_));
 BUF_X4 _10683_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[1] ),
    .Z(_05186_));
 MUX2_X1 _10684_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][51] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][51] ),
    .S(_05142_),
    .Z(_05187_));
 MUX2_X1 _10685_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][51] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][51] ),
    .S(_05142_),
    .Z(_05188_));
 MUX2_X2 _10686_ (.A(_05187_),
    .B(_05188_),
    .S(_05150_),
    .Z(_05189_));
 XNOR2_X1 _10687_ (.A(_05186_),
    .B(_05189_),
    .ZN(_05190_));
 BUF_X4 _10688_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[10] ),
    .Z(_05191_));
 MUX2_X1 _10689_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][60] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][60] ),
    .S(_05142_),
    .Z(_05192_));
 MUX2_X1 _10690_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][60] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][60] ),
    .S(_05142_),
    .Z(_05193_));
 MUX2_X2 _10691_ (.A(_05192_),
    .B(_05193_),
    .S(_05150_),
    .Z(_05194_));
 XNOR2_X1 _10692_ (.A(_05191_),
    .B(_05194_),
    .ZN(_05195_));
 NAND2_X2 _10693_ (.A1(_05190_),
    .A2(_05195_),
    .ZN(_05196_));
 BUF_X4 _10694_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[12] ),
    .Z(_05197_));
 MUX2_X1 _10695_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][62] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][62] ),
    .S(net736),
    .Z(_05198_));
 MUX2_X1 _10696_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][62] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][62] ),
    .S(net736),
    .Z(_05199_));
 INV_X2 _10697_ (.A(_05150_),
    .ZN(_05200_));
 BUF_X4 _10698_ (.A(_05200_),
    .Z(_05201_));
 MUX2_X1 _10699_ (.A(_05198_),
    .B(_05199_),
    .S(_05201_),
    .Z(_05202_));
 XNOR2_X2 _10700_ (.A(_05197_),
    .B(_05202_),
    .ZN(_05203_));
 BUF_X4 _10701_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[6] ),
    .Z(_05204_));
 MUX2_X1 _10702_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][56] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][56] ),
    .S(net736),
    .Z(_05205_));
 MUX2_X1 _10703_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][56] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][56] ),
    .S(net736),
    .Z(_05206_));
 MUX2_X1 _10704_ (.A(_05205_),
    .B(_05206_),
    .S(_05201_),
    .Z(_05207_));
 XNOR2_X2 _10705_ (.A(_05204_),
    .B(_05207_),
    .ZN(_05208_));
 BUF_X4 _10706_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[5] ),
    .Z(_05209_));
 MUX2_X1 _10707_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][55] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][55] ),
    .S(net736),
    .Z(_05210_));
 CLKBUF_X3 _10708_ (.A(net672),
    .Z(_05211_));
 MUX2_X1 _10709_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][55] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][55] ),
    .S(_05211_),
    .Z(_05212_));
 MUX2_X1 _10710_ (.A(_05210_),
    .B(_05212_),
    .S(_05201_),
    .Z(_05213_));
 XNOR2_X2 _10711_ (.A(_05209_),
    .B(_05213_),
    .ZN(_05214_));
 BUF_X4 _10712_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[8] ),
    .Z(_05215_));
 MUX2_X1 _10713_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][58] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][58] ),
    .S(_05211_),
    .Z(_05216_));
 MUX2_X1 _10714_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][58] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][58] ),
    .S(_05211_),
    .Z(_05217_));
 MUX2_X1 _10715_ (.A(_05216_),
    .B(_05217_),
    .S(_05201_),
    .Z(_05218_));
 XNOR2_X2 _10716_ (.A(_05215_),
    .B(_05218_),
    .ZN(_05219_));
 NAND4_X4 _10717_ (.A1(_05203_),
    .A2(_05208_),
    .A3(_05214_),
    .A4(_05219_),
    .ZN(_05220_));
 BUF_X4 _10718_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[13] ),
    .Z(_05221_));
 MUX2_X1 _10719_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][63] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][63] ),
    .S(_05211_),
    .Z(_05222_));
 MUX2_X1 _10720_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][63] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][63] ),
    .S(_05211_),
    .Z(_05223_));
 MUX2_X1 _10721_ (.A(_05222_),
    .B(_05223_),
    .S(_05201_),
    .Z(_05224_));
 XNOR2_X1 _10722_ (.A(_05221_),
    .B(_05224_),
    .ZN(_05225_));
 BUF_X4 _10723_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[9] ),
    .Z(_05226_));
 MUX2_X1 _10724_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][59] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][59] ),
    .S(_05211_),
    .Z(_05227_));
 MUX2_X1 _10725_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][59] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][59] ),
    .S(_05211_),
    .Z(_05228_));
 MUX2_X1 _10726_ (.A(_05227_),
    .B(_05228_),
    .S(_05201_),
    .Z(_05229_));
 XNOR2_X1 _10727_ (.A(_05226_),
    .B(_05229_),
    .ZN(_05230_));
 BUF_X4 _10728_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[7] ),
    .Z(_05231_));
 MUX2_X1 _10729_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][57] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][57] ),
    .S(_05211_),
    .Z(_05232_));
 MUX2_X1 _10730_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][57] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][57] ),
    .S(_05141_),
    .Z(_05233_));
 MUX2_X1 _10731_ (.A(_05232_),
    .B(_05233_),
    .S(_05200_),
    .Z(_05234_));
 XNOR2_X1 _10732_ (.A(_05231_),
    .B(_05234_),
    .ZN(_05235_));
 BUF_X4 _10733_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[11] ),
    .Z(_05236_));
 MUX2_X1 _10734_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][61] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][61] ),
    .S(net735),
    .Z(_05237_));
 MUX2_X1 _10735_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][61] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][61] ),
    .S(net735),
    .Z(_05238_));
 MUX2_X1 _10736_ (.A(_05237_),
    .B(_05238_),
    .S(_05200_),
    .Z(_05239_));
 XNOR2_X1 _10737_ (.A(_05236_),
    .B(_05239_),
    .ZN(_05240_));
 NAND4_X2 _10738_ (.A1(_05225_),
    .A2(_05230_),
    .A3(_05235_),
    .A4(_05240_),
    .ZN(_05241_));
 BUF_X4 _10739_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[3] ),
    .Z(_05242_));
 MUX2_X1 _10740_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][53] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][53] ),
    .S(_05211_),
    .Z(_05243_));
 MUX2_X1 _10741_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][53] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][53] ),
    .S(_05211_),
    .Z(_05244_));
 MUX2_X1 _10742_ (.A(_05243_),
    .B(_05244_),
    .S(_05201_),
    .Z(_05245_));
 XNOR2_X1 _10743_ (.A(_05242_),
    .B(_05245_),
    .ZN(_05246_));
 BUF_X4 _10744_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[0] ),
    .Z(_05247_));
 MUX2_X1 _10745_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][50] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][50] ),
    .S(net735),
    .Z(_05248_));
 MUX2_X1 _10746_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][50] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][50] ),
    .S(net735),
    .Z(_05249_));
 MUX2_X1 _10747_ (.A(_05248_),
    .B(_05249_),
    .S(_05200_),
    .Z(_05250_));
 XNOR2_X1 _10748_ (.A(_05247_),
    .B(_05250_),
    .ZN(_05251_));
 BUF_X4 _10749_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[4] ),
    .Z(_05252_));
 MUX2_X1 _10750_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][54] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][54] ),
    .S(_05141_),
    .Z(_05253_));
 MUX2_X1 _10751_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][54] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][54] ),
    .S(net735),
    .Z(_05254_));
 MUX2_X1 _10752_ (.A(_05253_),
    .B(_05254_),
    .S(_05200_),
    .Z(_05255_));
 XNOR2_X1 _10753_ (.A(_05252_),
    .B(_05255_),
    .ZN(_05256_));
 BUF_X4 _10754_ (.A(\dynamic_node_top.east_input.control.my_chip_id_in[2] ),
    .Z(_05257_));
 MUX2_X1 _10755_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][52] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][52] ),
    .S(_05141_),
    .Z(_05258_));
 MUX2_X1 _10756_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][52] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][52] ),
    .S(_05141_),
    .Z(_05259_));
 MUX2_X1 _10757_ (.A(_05258_),
    .B(_05259_),
    .S(_05200_),
    .Z(_05260_));
 XNOR2_X1 _10758_ (.A(_05257_),
    .B(_05260_),
    .ZN(_05261_));
 NAND4_X2 _10759_ (.A1(_05246_),
    .A2(_05251_),
    .A3(_05256_),
    .A4(_05261_),
    .ZN(_05262_));
 NOR4_X4 _10760_ (.A1(_05196_),
    .A2(_05220_),
    .A3(_05241_),
    .A4(_05262_),
    .ZN(_05263_));
 NAND4_X4 _10761_ (.A1(_10230_),
    .A2(_10233_),
    .A3(_10236_),
    .A4(_10239_),
    .ZN(_05264_));
 NAND4_X1 _10762_ (.A1(_10242_),
    .A2(_10245_),
    .A3(_10248_),
    .A4(_10251_),
    .ZN(_05265_));
 NOR2_X4 _10763_ (.A1(net734),
    .A2(_05265_),
    .ZN(_05266_));
 AND4_X2 _10764_ (.A1(_10275_),
    .A2(_10272_),
    .A3(_10254_),
    .A4(_10257_),
    .ZN(_05267_));
 AND2_X2 _10765_ (.A1(_10269_),
    .A2(_10266_),
    .ZN(_05268_));
 AND4_X4 _10766_ (.A1(_10260_),
    .A2(_10263_),
    .A3(_05267_),
    .A4(_05268_),
    .ZN(_05269_));
 NAND2_X4 _10767_ (.A1(_05266_),
    .A2(_05269_),
    .ZN(_05270_));
 MUX2_X1 _10768_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][30] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][30] ),
    .S(net739),
    .Z(_05271_));
 MUX2_X1 _10769_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][30] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][30] ),
    .S(net739),
    .Z(_05272_));
 MUX2_X2 _10770_ (.A(_05271_),
    .B(_05272_),
    .S(_05151_),
    .Z(_05273_));
 INV_X2 _10771_ (.A(_05273_),
    .ZN(_05274_));
 MUX2_X1 _10772_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][32] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][32] ),
    .S(net738),
    .Z(_05275_));
 MUX2_X1 _10773_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][32] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][32] ),
    .S(net738),
    .Z(_05276_));
 MUX2_X2 _10774_ (.A(_05275_),
    .B(_05276_),
    .S(_05152_),
    .Z(_05277_));
 MUX2_X1 _10775_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][31] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][31] ),
    .S(net739),
    .Z(_05278_));
 OR2_X1 _10776_ (.A1(_05152_),
    .A2(_05278_),
    .ZN(_05279_));
 MUX2_X1 _10777_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][31] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][31] ),
    .S(net738),
    .Z(_05280_));
 OAI21_X2 _10778_ (.A(_05279_),
    .B1(_05280_),
    .B2(_05201_),
    .ZN(_05281_));
 NAND3_X2 _10779_ (.A1(_05274_),
    .A2(_05277_),
    .A3(_05281_),
    .ZN(_05282_));
 NOR2_X4 _10780_ (.A1(_05270_),
    .A2(_05282_),
    .ZN(_05283_));
 INV_X1 _10781_ (.A(_05264_),
    .ZN(_05284_));
 INV_X1 _10782_ (.A(_10241_),
    .ZN(_05285_));
 INV_X1 _10783_ (.A(_10247_),
    .ZN(_05286_));
 INV_X1 _10784_ (.A(_10248_),
    .ZN(_05287_));
 OAI21_X2 _10785_ (.A(_05286_),
    .B1(_05287_),
    .B2(_10250_),
    .ZN(_05288_));
 AOI21_X2 _10786_ (.A(_10244_),
    .B1(_05288_),
    .B2(_10245_),
    .ZN(_05289_));
 INV_X1 _10787_ (.A(_10242_),
    .ZN(_05290_));
 OAI21_X2 _10788_ (.A(_05285_),
    .B1(_05289_),
    .B2(_05290_),
    .ZN(_05291_));
 INV_X1 _10789_ (.A(_10232_),
    .ZN(_05292_));
 AOI21_X1 _10790_ (.A(_10235_),
    .B1(_10236_),
    .B2(_10238_),
    .ZN(_05293_));
 INV_X1 _10791_ (.A(_10233_),
    .ZN(_05294_));
 OAI21_X1 _10792_ (.A(_05292_),
    .B1(_05293_),
    .B2(_05294_),
    .ZN(_05295_));
 AOI221_X2 _10793_ (.A(_10229_),
    .B1(_05284_),
    .B2(_05291_),
    .C1(_05295_),
    .C2(net635),
    .ZN(_05296_));
 OAI21_X4 _10794_ (.A(_05263_),
    .B1(_05283_),
    .B2(net770),
    .ZN(_05297_));
 NOR4_X4 _10795_ (.A1(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .A2(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .A3(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .A4(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .ZN(_05298_));
 NOR4_X4 _10796_ (.A1(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .A2(\dynamic_node_top.east_input.control.my_loc_x_in[0] ),
    .A3(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .A4(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .ZN(_05299_));
 AND2_X2 _10797_ (.A1(_05298_),
    .A2(_05299_),
    .ZN(_05300_));
 NOR4_X4 _10798_ (.A1(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .A2(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .A3(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .A4(\dynamic_node_top.east_input.control.my_loc_y_in[0] ),
    .ZN(_05301_));
 NOR4_X4 _10799_ (.A1(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .A2(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .A3(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .A4(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .ZN(_05302_));
 AND2_X2 _10800_ (.A1(_05301_),
    .A2(_05302_),
    .ZN(_05303_));
 NAND2_X4 _10801_ (.A1(_05300_),
    .A2(_05303_),
    .ZN(_05304_));
 OR3_X2 _10802_ (.A1(_05282_),
    .A2(_05263_),
    .A3(_05304_),
    .ZN(_05305_));
 AOI21_X4 _10803_ (.A(_05185_),
    .B1(_05297_),
    .B2(_05305_),
    .ZN(_05306_));
 INV_X2 _10804_ (.A(_00046_),
    .ZN(_05307_));
 OAI21_X4 _10805_ (.A(_05184_),
    .B1(_05306_),
    .B2(_05307_),
    .ZN(_05308_));
 INV_X2 _10806_ (.A(_05308_),
    .ZN(net621));
 BUF_X8 _10807_ (.A(_00008_),
    .Z(_05309_));
 BUF_X32 _10808_ (.A(_05309_),
    .Z(_05310_));
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 BUF_X16 _10810_ (.A(_05310_),
    .Z(_05312_));
 MUX2_X1 _10811_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][42] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][42] ),
    .S(_05312_),
    .Z(_05313_));
 BUF_X32 _10812_ (.A(_05310_),
    .Z(_05314_));
 BUF_X32 _10813_ (.A(_05314_),
    .Z(_05315_));
 MUX2_X1 _10814_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][42] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][42] ),
    .S(_05315_),
    .Z(_05316_));
 BUF_X8 _10815_ (.A(_00007_),
    .Z(_05317_));
 AOI21_X2 clone1 (.A(_05345_),
    .B1(_05454_),
    .B2(_05452_),
    .ZN(net1));
 BUF_X8 _10817_ (.A(_05317_),
    .Z(_05319_));
 BUF_X4 _10818_ (.A(_05319_),
    .Z(_05320_));
 BUF_X8 _10819_ (.A(_05320_),
    .Z(_05321_));
 MUX2_X2 _10820_ (.A(_05313_),
    .B(_05316_),
    .S(_05321_),
    .Z(_10276_));
 MUX2_X1 _10821_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][34] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][34] ),
    .S(_05314_),
    .Z(_05322_));
 OR2_X1 _10822_ (.A1(_05320_),
    .A2(_05322_),
    .ZN(_05323_));
 MUX2_X1 _10823_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][34] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][34] ),
    .S(_05312_),
    .Z(_05324_));
 INV_X2 _10824_ (.A(_05317_),
    .ZN(_05325_));
 BUF_X8 _10825_ (.A(_05325_),
    .Z(_05326_));
 OAI21_X4 _10826_ (.A(_05323_),
    .B1(_05324_),
    .B2(_05326_),
    .ZN(_05327_));
 INV_X1 _10827_ (.A(_05327_),
    .ZN(_10321_));
 BUF_X4 _10828_ (.A(_00048_),
    .Z(_05328_));
 CLKBUF_X3 _10829_ (.A(\dynamic_node_top.south_output.control.current_route_f[4] ),
    .Z(_05329_));
 CLKBUF_X3 _10830_ (.A(\dynamic_node_top.south_output.control.current_route_f[2] ),
    .Z(_05330_));
 CLKBUF_X3 _10831_ (.A(\dynamic_node_top.south_output.control.current_route_f[3] ),
    .Z(_05331_));
 CLKBUF_X3 _10832_ (.A(\dynamic_node_top.south_output.control.current_route_f[1] ),
    .Z(_05332_));
 NOR4_X4 _10833_ (.A1(_05329_),
    .A2(_05330_),
    .A3(_05331_),
    .A4(_05332_),
    .ZN(_05333_));
 AND2_X1 _10834_ (.A1(_05328_),
    .A2(_05333_),
    .ZN(_05334_));
 INV_X1 _10835_ (.A(\dynamic_node_top.south_output.space.is_one_f ),
    .ZN(_05335_));
 NOR2_X1 _10836_ (.A1(_05335_),
    .A2(\dynamic_node_top.south_output.space.valid_f ),
    .ZN(_05336_));
 NOR3_X2 _10837_ (.A1(\dynamic_node_top.south_output.space.is_two_or_more_f ),
    .A2(\dynamic_node_top.south_output.space.yummy_f ),
    .A3(_05336_),
    .ZN(_05337_));
 BUF_X2 _10838_ (.A(\dynamic_node_top.south_output.control.current_route_f[0] ),
    .Z(_05338_));
 AOI22_X1 _10839_ (.A1(_05338_),
    .A2(_05168_),
    .B1(_05177_),
    .B2(_05331_),
    .ZN(_05339_));
 INV_X1 _10840_ (.A(_00047_),
    .ZN(_05340_));
 AOI22_X1 _10841_ (.A1(_05340_),
    .A2(_05170_),
    .B1(_05175_),
    .B2(_05330_),
    .ZN(_05341_));
 NAND2_X1 _10842_ (.A1(_05339_),
    .A2(_05341_),
    .ZN(_05342_));
 AOI21_X1 _10843_ (.A(_05342_),
    .B1(_05182_),
    .B2(_05329_),
    .ZN(_05343_));
 NOR3_X2 _10844_ (.A1(_05334_),
    .A2(_05337_),
    .A3(_05343_),
    .ZN(_05344_));
 INV_X1 _10845_ (.A(_05344_),
    .ZN(_05345_));
 NAND2_X1 _10846_ (.A1(\dynamic_node_top.north_input.control.header_last_temp ),
    .A2(_05168_),
    .ZN(_05346_));
 AND4_X2 _10847_ (.A1(_10281_),
    .A2(_10284_),
    .A3(_10287_),
    .A4(_10290_),
    .ZN(_05347_));
 AND2_X2 _10848_ (.A1(_10296_),
    .A2(_10299_),
    .ZN(_05348_));
 NAND4_X4 _10849_ (.A1(_10278_),
    .A2(_10293_),
    .A3(_05347_),
    .A4(_05348_),
    .ZN(_05349_));
 NOR2_X2 _10850_ (.A1(_05349_),
    .A2(_05346_),
    .ZN(_05350_));
 AND4_X4 _10851_ (.A1(_10308_),
    .A2(_10305_),
    .A3(_10302_),
    .A4(_10311_),
    .ZN(_05351_));
 AOI21_X1 _10852_ (.A(_10313_),
    .B1(_10316_),
    .B2(net681),
    .ZN(_05352_));
 NAND2_X1 _10853_ (.A1(net681),
    .A2(_10317_),
    .ZN(_05353_));
 INV_X1 _10854_ (.A(_10322_),
    .ZN(_05354_));
 AOI21_X1 _10855_ (.A(_10319_),
    .B1(_05354_),
    .B2(_10320_),
    .ZN(_05355_));
 OAI21_X1 _10856_ (.A(_05352_),
    .B1(_05353_),
    .B2(_05355_),
    .ZN(_05356_));
 INV_X1 _10857_ (.A(_10304_),
    .ZN(_05357_));
 AOI21_X1 _10858_ (.A(_10307_),
    .B1(net633),
    .B2(_10310_),
    .ZN(_05358_));
 INV_X1 _10859_ (.A(_10305_),
    .ZN(_05359_));
 OAI21_X1 _10860_ (.A(_05357_),
    .B1(_05358_),
    .B2(_05359_),
    .ZN(_05360_));
 AOI221_X2 _10861_ (.A(_10301_),
    .B1(_05351_),
    .B2(_05356_),
    .C1(_05360_),
    .C2(net691),
    .ZN(_05361_));
 CLKBUF_X3 _10862_ (.A(net728),
    .Z(_05362_));
 MUX2_X1 _10863_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][30] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][30] ),
    .S(_05362_),
    .Z(_05363_));
 OR2_X1 _10864_ (.A1(_05320_),
    .A2(_05363_),
    .ZN(_05364_));
 MUX2_X1 _10865_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][30] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][30] ),
    .S(net726),
    .Z(_05365_));
 OAI21_X2 _10866_ (.A(_05364_),
    .B1(_05365_),
    .B2(_05325_),
    .ZN(_05366_));
 MUX2_X1 _10867_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][32] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][32] ),
    .S(net728),
    .Z(_05367_));
 MUX2_X1 _10868_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][32] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][32] ),
    .S(net726),
    .Z(_05368_));
 MUX2_X1 _10869_ (.A(_05367_),
    .B(_05368_),
    .S(_05319_),
    .Z(_05369_));
 BUF_X4 _10870_ (.A(_05369_),
    .Z(_05370_));
 MUX2_X1 _10871_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][31] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][31] ),
    .S(net728),
    .Z(_05371_));
 NOR2_X2 _10872_ (.A1(_05319_),
    .A2(_05371_),
    .ZN(_05372_));
 MUX2_X1 _10873_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][31] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][31] ),
    .S(net728),
    .Z(_05373_));
 NOR2_X1 _10874_ (.A1(_05325_),
    .A2(_05373_),
    .ZN(_05374_));
 OR2_X1 _10875_ (.A1(_05372_),
    .A2(_05374_),
    .ZN(_05375_));
 CLKBUF_X3 _10876_ (.A(_05375_),
    .Z(_05376_));
 AND2_X2 _10877_ (.A1(_10314_),
    .A2(_10317_),
    .ZN(_05377_));
 AND2_X2 _10878_ (.A1(_10323_),
    .A2(_10320_),
    .ZN(_05378_));
 NAND3_X4 _10879_ (.A1(_05351_),
    .A2(_05377_),
    .A3(_05378_),
    .ZN(_05379_));
 NOR4_X4 _10880_ (.A1(_05379_),
    .A2(_05370_),
    .A3(_05376_),
    .A4(_05366_),
    .ZN(_05380_));
 OAI21_X1 _10881_ (.A(_05350_),
    .B1(_05380_),
    .B2(_05361_),
    .ZN(_05381_));
 NAND2_X4 _10882_ (.A1(_05298_),
    .A2(_05299_),
    .ZN(_05382_));
 NAND2_X4 _10883_ (.A1(_05301_),
    .A2(_05302_),
    .ZN(_05383_));
 NOR2_X2 _10884_ (.A1(_05382_),
    .A2(_05383_),
    .ZN(_05384_));
 AND2_X1 _10885_ (.A1(\dynamic_node_top.north_input.control.header_last_temp ),
    .A2(_05168_),
    .ZN(_05385_));
 BUF_X4 _10886_ (.A(_05385_),
    .Z(_05386_));
 NOR3_X1 _10887_ (.A1(_05366_),
    .A2(_05370_),
    .A3(_05376_),
    .ZN(_05387_));
 NAND3_X1 _10888_ (.A1(_05384_),
    .A2(_05386_),
    .A3(_05387_),
    .ZN(_05388_));
 BUF_X4 _10889_ (.A(net678),
    .Z(_05389_));
 MUX2_X1 _10890_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][59] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][59] ),
    .S(_05389_),
    .Z(_05390_));
 MUX2_X1 _10891_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][59] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][59] ),
    .S(_05389_),
    .Z(_05391_));
 MUX2_X1 _10892_ (.A(_05390_),
    .B(_05391_),
    .S(_05317_),
    .Z(_05392_));
 XNOR2_X2 _10893_ (.A(_05226_),
    .B(_05392_),
    .ZN(_05393_));
 MUX2_X1 _10894_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][58] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][58] ),
    .S(_05389_),
    .Z(_05394_));
 MUX2_X1 _10895_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][58] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][58] ),
    .S(_05389_),
    .Z(_05395_));
 MUX2_X1 _10896_ (.A(_05394_),
    .B(_05395_),
    .S(_05317_),
    .Z(_05396_));
 XNOR2_X2 _10897_ (.A(_05215_),
    .B(_05396_),
    .ZN(_05397_));
 MUX2_X1 _10898_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][56] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][56] ),
    .S(_05389_),
    .Z(_05398_));
 MUX2_X1 _10899_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][56] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][56] ),
    .S(_05389_),
    .Z(_05399_));
 MUX2_X1 _10900_ (.A(_05398_),
    .B(_05399_),
    .S(_05317_),
    .Z(_05400_));
 XNOR2_X2 _10901_ (.A(_05204_),
    .B(_05400_),
    .ZN(_05401_));
 MUX2_X1 _10902_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][63] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][63] ),
    .S(_05389_),
    .Z(_05402_));
 MUX2_X1 _10903_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][63] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][63] ),
    .S(_05389_),
    .Z(_05403_));
 MUX2_X1 _10904_ (.A(_05402_),
    .B(_05403_),
    .S(_05317_),
    .Z(_05404_));
 XNOR2_X2 _10905_ (.A(_05221_),
    .B(_05404_),
    .ZN(_05405_));
 NAND4_X4 _10906_ (.A1(_05393_),
    .A2(_05397_),
    .A3(_05401_),
    .A4(_05405_),
    .ZN(_05406_));
 MUX2_X1 _10907_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][54] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][54] ),
    .S(_05389_),
    .Z(_05407_));
 CLKBUF_X3 _10908_ (.A(net662),
    .Z(_05408_));
 MUX2_X1 _10909_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][54] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][54] ),
    .S(_05408_),
    .Z(_05409_));
 MUX2_X1 _10910_ (.A(_05407_),
    .B(_05409_),
    .S(_05317_),
    .Z(_05410_));
 XNOR2_X2 _10911_ (.A(_05252_),
    .B(_05410_),
    .ZN(_05411_));
 MUX2_X1 _10912_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][51] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][51] ),
    .S(_05408_),
    .Z(_05412_));
 MUX2_X1 _10913_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][51] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][51] ),
    .S(_05408_),
    .Z(_05413_));
 MUX2_X1 _10914_ (.A(_05412_),
    .B(_05413_),
    .S(_05317_),
    .Z(_05414_));
 XNOR2_X2 _10915_ (.A(_05186_),
    .B(_05414_),
    .ZN(_05415_));
 MUX2_X1 _10916_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][52] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][52] ),
    .S(_05408_),
    .Z(_05416_));
 MUX2_X1 _10917_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][52] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][52] ),
    .S(_05408_),
    .Z(_05417_));
 MUX2_X1 _10918_ (.A(_05416_),
    .B(_05417_),
    .S(_05317_),
    .Z(_05418_));
 XNOR2_X2 _10919_ (.A(_05257_),
    .B(_05418_),
    .ZN(_05419_));
 MUX2_X1 _10920_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][55] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][55] ),
    .S(_05408_),
    .Z(_05420_));
 MUX2_X1 _10921_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][55] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][55] ),
    .S(_05408_),
    .Z(_05421_));
 MUX2_X1 _10922_ (.A(_05420_),
    .B(_05421_),
    .S(_05317_),
    .Z(_05422_));
 XNOR2_X2 _10923_ (.A(_05209_),
    .B(_05422_),
    .ZN(_05423_));
 NAND4_X4 _10924_ (.A1(_05411_),
    .A2(_05415_),
    .A3(_05419_),
    .A4(_05423_),
    .ZN(_05424_));
 MUX2_X1 _10925_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][60] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][60] ),
    .S(net2),
    .Z(_05425_));
 MUX2_X1 _10926_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][60] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][60] ),
    .S(net2),
    .Z(_05426_));
 MUX2_X2 _10927_ (.A(_05425_),
    .B(_05426_),
    .S(_05317_),
    .Z(_05427_));
 XNOR2_X2 _10928_ (.A(_05191_),
    .B(_05427_),
    .ZN(_05428_));
 MUX2_X1 _10929_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][50] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][50] ),
    .S(net2),
    .Z(_05429_));
 MUX2_X1 _10930_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][50] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][50] ),
    .S(net677),
    .Z(_05430_));
 MUX2_X1 _10931_ (.A(_05429_),
    .B(_05430_),
    .S(_05317_),
    .Z(_05431_));
 XNOR2_X2 _10932_ (.A(_05247_),
    .B(_05431_),
    .ZN(_05432_));
 MUX2_X1 _10933_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][62] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][62] ),
    .S(net2),
    .Z(_05433_));
 MUX2_X1 _10934_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][62] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][62] ),
    .S(net677),
    .Z(_05434_));
 MUX2_X1 _10935_ (.A(_05433_),
    .B(_05434_),
    .S(_05317_),
    .Z(_05435_));
 XNOR2_X2 _10936_ (.A(_05197_),
    .B(_05435_),
    .ZN(_05436_));
 MUX2_X1 _10937_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][61] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][61] ),
    .S(net2),
    .Z(_05437_));
 MUX2_X1 _10938_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][61] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][61] ),
    .S(net677),
    .Z(_05438_));
 MUX2_X1 _10939_ (.A(_05437_),
    .B(_05438_),
    .S(_05317_),
    .Z(_05439_));
 XNOR2_X2 _10940_ (.A(_05236_),
    .B(_05439_),
    .ZN(_05440_));
 NAND4_X4 _10941_ (.A1(_05428_),
    .A2(_05432_),
    .A3(_05436_),
    .A4(_05440_),
    .ZN(_05441_));
 MUX2_X1 _10942_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][57] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][57] ),
    .S(_05389_),
    .Z(_05442_));
 MUX2_X1 _10943_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][57] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][57] ),
    .S(_05408_),
    .Z(_05443_));
 MUX2_X1 _10944_ (.A(_05442_),
    .B(_05443_),
    .S(_05317_),
    .Z(_05444_));
 XNOR2_X1 _10945_ (.A(_05231_),
    .B(_05444_),
    .ZN(_05445_));
 MUX2_X1 _10946_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][53] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][53] ),
    .S(_05408_),
    .Z(_05446_));
 MUX2_X1 _10947_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][53] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][53] ),
    .S(_05408_),
    .Z(_05447_));
 MUX2_X1 _10948_ (.A(_05446_),
    .B(_05447_),
    .S(_05317_),
    .Z(_05448_));
 XNOR2_X1 _10949_ (.A(_05242_),
    .B(_05448_),
    .ZN(_05449_));
 NAND2_X2 _10950_ (.A1(_05445_),
    .A2(_05449_),
    .ZN(_05450_));
 OR4_X4 _10951_ (.A1(_05406_),
    .A2(_05424_),
    .A3(_05441_),
    .A4(_05450_),
    .ZN(_05451_));
 MUX2_X2 _10952_ (.A(_05381_),
    .B(_05388_),
    .S(_05451_),
    .Z(_05452_));
 BUF_X1 rebuffer100 (.A(_07420_),
    .Z(net752));
 BUF_X2 _10954_ (.A(_00049_),
    .Z(_05454_));
 AOI21_X4 _10955_ (.A(_05345_),
    .B1(_05454_),
    .B2(_05452_),
    .ZN(net624));
 BUF_X8 _10956_ (.A(_00006_),
    .Z(_05455_));
 BUF_X32 _10957_ (.A(_05455_),
    .Z(_05456_));
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 BUF_X32 _10959_ (.A(_05456_),
    .Z(_05458_));
 BUF_X32 _10960_ (.A(_05458_),
    .Z(_05459_));
 MUX2_X1 _10961_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][42] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][42] ),
    .S(_05459_),
    .Z(_05460_));
 MUX2_X1 _10962_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][42] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][42] ),
    .S(_05459_),
    .Z(_05461_));
 BUF_X4 _10963_ (.A(_00005_),
    .Z(_05462_));
 BUF_X8 _10964_ (.A(_05462_),
    .Z(_05463_));
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 BUF_X2 _10966_ (.A(_05463_),
    .Z(_05465_));
 MUX2_X2 _10967_ (.A(_05460_),
    .B(_05461_),
    .S(_05465_),
    .Z(_10345_));
 MUX2_X1 _10968_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][34] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][34] ),
    .S(net721),
    .Z(_05466_));
 MUX2_X1 _10969_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][34] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][34] ),
    .S(net721),
    .Z(_05467_));
 CLKBUF_X3 _10970_ (.A(_05463_),
    .Z(_05468_));
 MUX2_X2 _10971_ (.A(_05466_),
    .B(_05467_),
    .S(_05468_),
    .Z(_10348_));
 INV_X4 _10972_ (.A(_00051_),
    .ZN(_05469_));
 BUF_X4 _10973_ (.A(\dynamic_node_top.west_output.control.current_route_f[3] ),
    .Z(_05470_));
 BUF_X2 _10974_ (.A(\dynamic_node_top.west_output.control.current_route_f[1] ),
    .Z(_05471_));
 NOR4_X4 _10975_ (.A1(\dynamic_node_top.west_output.control.current_route_f[4] ),
    .A2(\dynamic_node_top.west_output.control.current_route_f[2] ),
    .A3(_05470_),
    .A4(_05471_),
    .ZN(_05472_));
 INV_X1 _10976_ (.A(_05472_),
    .ZN(_05473_));
 NOR2_X2 _10977_ (.A1(_05469_),
    .A2(_05473_),
    .ZN(_05474_));
 INV_X1 _10978_ (.A(\dynamic_node_top.west_output.space.is_one_f ),
    .ZN(_05475_));
 NOR2_X1 _10979_ (.A1(_05475_),
    .A2(\dynamic_node_top.west_output.space.valid_f ),
    .ZN(_05476_));
 NOR3_X2 _10980_ (.A1(\dynamic_node_top.west_output.space.is_two_or_more_f ),
    .A2(\dynamic_node_top.west_output.space.yummy_f ),
    .A3(_05476_),
    .ZN(_05477_));
 CLKBUF_X3 _10981_ (.A(\dynamic_node_top.west_output.control.current_route_f[4] ),
    .Z(_05478_));
 INV_X1 _10982_ (.A(_00050_),
    .ZN(_05479_));
 AOI22_X1 _10983_ (.A1(_05478_),
    .A2(_05168_),
    .B1(_05175_),
    .B2(_05479_),
    .ZN(_05480_));
 CLKBUF_X3 _10984_ (.A(\dynamic_node_top.west_output.control.current_route_f[0] ),
    .Z(_05481_));
 AOI22_X1 _10985_ (.A1(_05470_),
    .A2(_05170_),
    .B1(_05177_),
    .B2(_05481_),
    .ZN(_05482_));
 NAND2_X1 _10986_ (.A1(_05480_),
    .A2(_05482_),
    .ZN(_05483_));
 CLKBUF_X3 _10987_ (.A(\dynamic_node_top.west_output.control.current_route_f[2] ),
    .Z(_05484_));
 AOI21_X1 _10988_ (.A(_05483_),
    .B1(_05182_),
    .B2(_05484_),
    .ZN(_05485_));
 NOR3_X1 _10989_ (.A1(_05474_),
    .A2(_05477_),
    .A3(_05485_),
    .ZN(_05486_));
 INV_X1 _10990_ (.A(_05486_),
    .ZN(_05487_));
 BUF_X2 _10991_ (.A(\dynamic_node_top.east_input.control.header_last_temp ),
    .Z(_05488_));
 NAND2_X4 _10992_ (.A1(_05488_),
    .A2(_05177_),
    .ZN(_05489_));
 MUX2_X1 _10993_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][30] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][30] ),
    .S(net700),
    .Z(_05490_));
 MUX2_X2 _10994_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][30] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][30] ),
    .S(net701),
    .Z(_05491_));
 MUX2_X2 _10995_ (.A(_05490_),
    .B(_05491_),
    .S(_05462_),
    .Z(_05492_));
 MUX2_X1 _10996_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][31] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][31] ),
    .S(net711),
    .Z(_05493_));
 NOR2_X2 _10997_ (.A1(_05463_),
    .A2(_05493_),
    .ZN(_05494_));
 INV_X4 _10998_ (.A(_05462_),
    .ZN(_05495_));
 MUX2_X1 _10999_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][31] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][31] ),
    .S(net711),
    .Z(_05496_));
 NOR2_X4 _11000_ (.A1(_05495_),
    .A2(_05496_),
    .ZN(_05497_));
 MUX2_X1 _11001_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][32] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][32] ),
    .S(net700),
    .Z(_05498_));
 MUX2_X2 _11002_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][32] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][32] ),
    .S(net700),
    .Z(_05499_));
 MUX2_X2 _11003_ (.A(_05498_),
    .B(_05499_),
    .S(_05462_),
    .Z(_05500_));
 NOR4_X2 _11004_ (.A1(_05492_),
    .A2(_05494_),
    .A3(_05497_),
    .A4(_05500_),
    .ZN(_05501_));
 AOI21_X1 _11005_ (.A(_05382_),
    .B1(_05303_),
    .B2(_05501_),
    .ZN(_05502_));
 OR2_X1 _11006_ (.A1(_05489_),
    .A2(_05502_),
    .ZN(_05503_));
 NAND2_X1 _11007_ (.A1(_10326_),
    .A2(_10329_),
    .ZN(_05504_));
 AOI21_X2 _11008_ (.A(_10325_),
    .B1(_10328_),
    .B2(net638),
    .ZN(_05505_));
 AND2_X1 _11009_ (.A1(_05504_),
    .A2(_05505_),
    .ZN(_05506_));
 NAND4_X2 _11010_ (.A1(_10335_),
    .A2(_10332_),
    .A3(_10344_),
    .A4(_10347_),
    .ZN(_05507_));
 NAND2_X1 _11011_ (.A1(_10338_),
    .A2(_10341_),
    .ZN(_05508_));
 OR3_X4 _11012_ (.A1(_05507_),
    .A2(_05504_),
    .A3(_05508_),
    .ZN(_05509_));
 NAND2_X1 _11013_ (.A1(_10368_),
    .A2(_10350_),
    .ZN(_05510_));
 NAND2_X2 _11014_ (.A1(_10371_),
    .A2(_10362_),
    .ZN(_05511_));
 NAND4_X2 _11015_ (.A1(_10365_),
    .A2(_10356_),
    .A3(_10359_),
    .A4(_10353_),
    .ZN(_05512_));
 NOR3_X4 _11016_ (.A1(_05512_),
    .A2(_05511_),
    .A3(_05510_),
    .ZN(_05513_));
 AOI21_X2 _11017_ (.A(net682),
    .B1(_05501_),
    .B2(_05513_),
    .ZN(_05514_));
 NAND2_X4 _11018_ (.A1(_05509_),
    .A2(_05505_),
    .ZN(_05515_));
 INV_X1 _11019_ (.A(_10331_),
    .ZN(_05516_));
 OAI21_X1 _11020_ (.A(net660),
    .B1(net637),
    .B2(_10334_),
    .ZN(_05517_));
 NAND2_X1 _11021_ (.A1(_05516_),
    .A2(_05517_),
    .ZN(_05518_));
 OR3_X1 _11022_ (.A1(_10331_),
    .A2(_10334_),
    .A3(_10337_),
    .ZN(_05519_));
 AOI21_X1 _11023_ (.A(_05519_),
    .B1(_10340_),
    .B2(net724),
    .ZN(_05520_));
 INV_X1 _11024_ (.A(_10346_),
    .ZN(_05521_));
 AOI21_X1 _11025_ (.A(_10343_),
    .B1(_05521_),
    .B2(net716),
    .ZN(_05522_));
 OAI21_X2 _11026_ (.A(_05520_),
    .B1(_05522_),
    .B2(_05508_),
    .ZN(_05523_));
 AOI21_X4 _11027_ (.A(_05515_),
    .B1(_05518_),
    .B2(_05523_),
    .ZN(_05524_));
 OR4_X4 _11028_ (.A1(_05489_),
    .A2(_05524_),
    .A3(_05514_),
    .A4(_05506_),
    .ZN(_05525_));
 MUX2_X1 _11029_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][58] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][58] ),
    .S(net711),
    .Z(_05526_));
 MUX2_X1 _11030_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][58] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][58] ),
    .S(net717),
    .Z(_05527_));
 MUX2_X1 _11031_ (.A(_05526_),
    .B(_05527_),
    .S(_05463_),
    .Z(_05528_));
 XNOR2_X1 _11032_ (.A(_05215_),
    .B(_05528_),
    .ZN(_05529_));
 MUX2_X1 _11033_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][51] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][51] ),
    .S(net717),
    .Z(_05530_));
 MUX2_X1 _11034_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][51] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][51] ),
    .S(net717),
    .Z(_05531_));
 CLKBUF_X3 _11035_ (.A(_05462_),
    .Z(_05532_));
 MUX2_X1 _11036_ (.A(_05530_),
    .B(_05531_),
    .S(_05532_),
    .Z(_05533_));
 XNOR2_X1 _11037_ (.A(_05186_),
    .B(_05533_),
    .ZN(_05534_));
 MUX2_X1 _11038_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][57] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][57] ),
    .S(net717),
    .Z(_05535_));
 BUF_X4 _11039_ (.A(net699),
    .Z(_05536_));
 MUX2_X1 _11040_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][57] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][57] ),
    .S(_05536_),
    .Z(_05537_));
 MUX2_X1 _11041_ (.A(_05535_),
    .B(_05537_),
    .S(_05532_),
    .Z(_05538_));
 XNOR2_X1 _11042_ (.A(_05231_),
    .B(_05538_),
    .ZN(_05539_));
 MUX2_X1 _11043_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][62] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][62] ),
    .S(_05536_),
    .Z(_05540_));
 MUX2_X2 _11044_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][62] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][62] ),
    .S(_05536_),
    .Z(_05541_));
 MUX2_X1 _11045_ (.A(_05540_),
    .B(_05541_),
    .S(_05532_),
    .Z(_05542_));
 XNOR2_X1 _11046_ (.A(_05197_),
    .B(_05542_),
    .ZN(_05543_));
 NAND4_X2 _11047_ (.A1(_05529_),
    .A2(_05534_),
    .A3(_05539_),
    .A4(_05543_),
    .ZN(_05544_));
 MUX2_X1 _11048_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][56] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][56] ),
    .S(_05536_),
    .Z(_05545_));
 MUX2_X1 _11049_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][56] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][56] ),
    .S(_05536_),
    .Z(_05546_));
 MUX2_X1 _11050_ (.A(_05545_),
    .B(_05546_),
    .S(_05532_),
    .Z(_05547_));
 XNOR2_X1 _11051_ (.A(_05204_),
    .B(_05547_),
    .ZN(_05548_));
 MUX2_X1 _11052_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][50] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][50] ),
    .S(_05536_),
    .Z(_05549_));
 BUF_X4 rebuffer120 (.A(_05296_),
    .Z(net770));
 MUX2_X1 _11054_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][50] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][50] ),
    .S(net708),
    .Z(_05551_));
 MUX2_X1 _11055_ (.A(_05549_),
    .B(_05551_),
    .S(_05532_),
    .Z(_05552_));
 XNOR2_X1 _11056_ (.A(_05247_),
    .B(_05552_),
    .ZN(_05553_));
 MUX2_X1 _11057_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][60] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][60] ),
    .S(net698),
    .Z(_05554_));
 MUX2_X1 _11058_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][60] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][60] ),
    .S(net708),
    .Z(_05555_));
 MUX2_X2 _11059_ (.A(_05554_),
    .B(_05555_),
    .S(_05462_),
    .Z(_05556_));
 XNOR2_X1 _11060_ (.A(_05191_),
    .B(_05556_),
    .ZN(_05557_));
 MUX2_X1 _11061_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][54] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][54] ),
    .S(net708),
    .Z(_05558_));
 MUX2_X1 _11062_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][54] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][54] ),
    .S(net708),
    .Z(_05559_));
 MUX2_X1 _11063_ (.A(_05558_),
    .B(_05559_),
    .S(_05532_),
    .Z(_05560_));
 XNOR2_X1 _11064_ (.A(_05252_),
    .B(_05560_),
    .ZN(_05561_));
 NAND4_X2 _11065_ (.A1(_05548_),
    .A2(_05553_),
    .A3(_05557_),
    .A4(_05561_),
    .ZN(_05562_));
 MUX2_X1 _11066_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][61] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][61] ),
    .S(net708),
    .Z(_05563_));
 MUX2_X1 _11067_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][61] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][61] ),
    .S(net708),
    .Z(_05564_));
 MUX2_X1 _11068_ (.A(_05563_),
    .B(_05564_),
    .S(_05532_),
    .Z(_05565_));
 XNOR2_X1 _11069_ (.A(_05236_),
    .B(_05565_),
    .ZN(_05566_));
 MUX2_X1 _11070_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][59] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][59] ),
    .S(net708),
    .Z(_05567_));
 MUX2_X1 _11071_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][59] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][59] ),
    .S(net708),
    .Z(_05568_));
 MUX2_X1 _11072_ (.A(_05567_),
    .B(_05568_),
    .S(_05532_),
    .Z(_05569_));
 XNOR2_X1 _11073_ (.A(_05226_),
    .B(_05569_),
    .ZN(_05570_));
 MUX2_X1 _11074_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][55] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][55] ),
    .S(net708),
    .Z(_05571_));
 MUX2_X1 _11075_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][55] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][55] ),
    .S(_05455_),
    .Z(_05572_));
 MUX2_X1 _11076_ (.A(_05571_),
    .B(_05572_),
    .S(_05462_),
    .Z(_05573_));
 XNOR2_X1 _11077_ (.A(_05209_),
    .B(_05573_),
    .ZN(_05574_));
 MUX2_X1 _11078_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][63] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][63] ),
    .S(net698),
    .Z(_05575_));
 MUX2_X1 _11079_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][63] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][63] ),
    .S(net698),
    .Z(_05576_));
 MUX2_X1 _11080_ (.A(_05575_),
    .B(_05576_),
    .S(_05462_),
    .Z(_05577_));
 XNOR2_X1 _11081_ (.A(_05221_),
    .B(_05577_),
    .ZN(_05578_));
 NAND4_X2 _11082_ (.A1(_05566_),
    .A2(_05570_),
    .A3(_05574_),
    .A4(_05578_),
    .ZN(_05579_));
 MUX2_X1 _11083_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][53] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][53] ),
    .S(_05536_),
    .Z(_05580_));
 MUX2_X1 _11084_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][53] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][53] ),
    .S(_05536_),
    .Z(_05581_));
 MUX2_X1 _11085_ (.A(_05580_),
    .B(_05581_),
    .S(_05532_),
    .Z(_05582_));
 XNOR2_X1 _11086_ (.A(_05242_),
    .B(_05582_),
    .ZN(_05583_));
 MUX2_X1 _11087_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][52] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][52] ),
    .S(_05536_),
    .Z(_05584_));
 MUX2_X1 _11088_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][52] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][52] ),
    .S(net708),
    .Z(_05585_));
 MUX2_X1 _11089_ (.A(_05584_),
    .B(_05585_),
    .S(_05532_),
    .Z(_05586_));
 XNOR2_X1 _11090_ (.A(_05257_),
    .B(_05586_),
    .ZN(_05587_));
 NAND2_X1 _11091_ (.A1(_05583_),
    .A2(_05587_),
    .ZN(_05588_));
 NOR4_X4 _11092_ (.A1(_05562_),
    .A2(_05579_),
    .A3(_05544_),
    .A4(_05588_),
    .ZN(_05589_));
 MUX2_X2 _11093_ (.A(_05503_),
    .B(_05525_),
    .S(_05589_),
    .Z(_05590_));
 BUF_X4 rebuffer107 (.A(net625),
    .Z(net756));
 AOI21_X4 _11095_ (.A(_05487_),
    .B1(_05590_),
    .B2(_00052_),
    .ZN(net625));
 CLKBUF_X3 _11096_ (.A(_00054_),
    .Z(_05592_));
 INV_X2 _11097_ (.A(_05592_),
    .ZN(_05593_));
 CLKBUF_X3 _11098_ (.A(\dynamic_node_top.proc_output.control.current_route_f[2] ),
    .Z(_05594_));
 CLKBUF_X3 _11099_ (.A(\dynamic_node_top.proc_output.control.current_route_f[3] ),
    .Z(_05595_));
 BUF_X2 _11100_ (.A(\dynamic_node_top.proc_output.control.current_route_f[1] ),
    .Z(_05596_));
 NOR4_X4 _11101_ (.A1(\dynamic_node_top.proc_output.control.current_route_f[4] ),
    .A2(_05594_),
    .A3(_05595_),
    .A4(_05596_),
    .ZN(_05597_));
 INV_X1 _11102_ (.A(_05597_),
    .ZN(_05598_));
 NOR2_X2 _11103_ (.A1(_05593_),
    .A2(_05598_),
    .ZN(_05599_));
 INV_X1 _11104_ (.A(\dynamic_node_top.proc_output.space.is_one_f ),
    .ZN(_05600_));
 NOR2_X1 _11105_ (.A1(_05600_),
    .A2(\dynamic_node_top.proc_output.space.valid_f ),
    .ZN(_05601_));
 NOR3_X1 _11106_ (.A1(\dynamic_node_top.proc_output.space.is_two_or_more_f ),
    .A2(\dynamic_node_top.proc_output.space.yummy_f ),
    .A3(_05601_),
    .ZN(_05602_));
 CLKBUF_X3 _11107_ (.A(\dynamic_node_top.proc_output.control.current_route_f[0] ),
    .Z(_05603_));
 AOI22_X1 _11108_ (.A1(_05594_),
    .A2(_05168_),
    .B1(_05170_),
    .B2(_05603_),
    .ZN(_05604_));
 BUF_X4 _11109_ (.A(\dynamic_node_top.proc_output.control.current_route_f[4] ),
    .Z(_05605_));
 AOI22_X1 _11110_ (.A1(_05595_),
    .A2(_05175_),
    .B1(_05177_),
    .B2(_05605_),
    .ZN(_05606_));
 NAND2_X1 _11111_ (.A1(_05604_),
    .A2(_05606_),
    .ZN(_05607_));
 INV_X1 _11112_ (.A(_00053_),
    .ZN(_05608_));
 AOI21_X1 _11113_ (.A(_05607_),
    .B1(_05182_),
    .B2(_05608_),
    .ZN(_05609_));
 OR3_X2 _11114_ (.A1(_05599_),
    .A2(_05602_),
    .A3(_05609_),
    .ZN(_05610_));
 MUX2_X1 _11115_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][32] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][32] ),
    .S(net746),
    .Z(_05611_));
 MUX2_X1 _11116_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][32] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][32] ),
    .S(net746),
    .Z(_05612_));
 MUX2_X2 _11117_ (.A(_05611_),
    .B(_05612_),
    .S(_05124_),
    .Z(_05613_));
 MUX2_X1 _11118_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][30] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][30] ),
    .S(net765),
    .Z(_05614_));
 MUX2_X1 _11119_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][30] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][30] ),
    .S(net746),
    .Z(_05615_));
 MUX2_X2 _11120_ (.A(_05614_),
    .B(_05615_),
    .S(_05124_),
    .Z(_05616_));
 NOR2_X2 _11121_ (.A1(_05613_),
    .A2(_05616_),
    .ZN(_05617_));
 NAND2_X1 _11122_ (.A1(\dynamic_node_top.south_input.control.header_last_temp ),
    .A2(_05170_),
    .ZN(_05618_));
 MUX2_X1 _11123_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][31] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][31] ),
    .S(net765),
    .Z(_05619_));
 MUX2_X1 _11124_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][31] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][31] ),
    .S(net765),
    .Z(_05620_));
 MUX2_X2 _11125_ (.A(_05619_),
    .B(_05620_),
    .S(_05124_),
    .Z(_05621_));
 NOR2_X1 _11126_ (.A1(_05618_),
    .A2(_05621_),
    .ZN(_05622_));
 NAND3_X1 _11127_ (.A1(_05384_),
    .A2(_05617_),
    .A3(_05622_),
    .ZN(_05623_));
 NAND2_X1 _11128_ (.A1(_05617_),
    .A2(_05622_),
    .ZN(_05624_));
 NAND4_X2 _11129_ (.A1(_10220_),
    .A2(_10214_),
    .A3(_10211_),
    .A4(_10223_),
    .ZN(_05625_));
 NAND4_X2 _11130_ (.A1(_10205_),
    .A2(_10217_),
    .A3(_10208_),
    .A4(_10227_),
    .ZN(_05626_));
 NOR2_X1 _11131_ (.A1(_05625_),
    .A2(_05626_),
    .ZN(_05627_));
 AND4_X2 _11132_ (.A1(_10190_),
    .A2(_10181_),
    .A3(_10199_),
    .A4(_10184_),
    .ZN(_05628_));
 AND2_X1 _11133_ (.A1(_10187_),
    .A2(_10202_),
    .ZN(_05629_));
 AND4_X4 _11134_ (.A1(_10193_),
    .A2(_10196_),
    .A3(_05628_),
    .A4(_05629_),
    .ZN(_05630_));
 NAND2_X1 _11135_ (.A1(_05627_),
    .A2(_05630_),
    .ZN(_05631_));
 OR2_X1 _11136_ (.A1(_05624_),
    .A2(_05631_),
    .ZN(_05632_));
 MUX2_X1 _11137_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][63] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][63] ),
    .S(net687),
    .Z(_05633_));
 MUX2_X1 _11138_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][63] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][63] ),
    .S(net687),
    .Z(_05634_));
 MUX2_X1 _11139_ (.A(_05633_),
    .B(_05634_),
    .S(_05124_),
    .Z(_05635_));
 XNOR2_X2 _11140_ (.A(_05221_),
    .B(_05635_),
    .ZN(_05636_));
 MUX2_X1 _11141_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][60] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][60] ),
    .S(net687),
    .Z(_05637_));
 MUX2_X1 _11142_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][60] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][60] ),
    .S(net687),
    .Z(_05638_));
 MUX2_X2 _11143_ (.A(_05637_),
    .B(_05638_),
    .S(_05124_),
    .Z(_05639_));
 XNOR2_X2 _11144_ (.A(_05191_),
    .B(_05639_),
    .ZN(_05640_));
 MUX2_X1 _11145_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][53] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][53] ),
    .S(_05129_),
    .Z(_05641_));
 MUX2_X1 _11146_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][53] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][53] ),
    .S(net687),
    .Z(_05642_));
 CLKBUF_X3 _11147_ (.A(_05124_),
    .Z(_05643_));
 MUX2_X1 _11148_ (.A(_05641_),
    .B(_05642_),
    .S(_05643_),
    .Z(_05644_));
 XNOR2_X2 _11149_ (.A(_05242_),
    .B(_05644_),
    .ZN(_05645_));
 BUF_X4 _11150_ (.A(net679),
    .Z(_05646_));
 MUX2_X1 _11151_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][51] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][51] ),
    .S(_05646_),
    .Z(_05647_));
 MUX2_X1 _11152_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][51] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][51] ),
    .S(_05129_),
    .Z(_05648_));
 MUX2_X2 _11153_ (.A(_05647_),
    .B(_05648_),
    .S(_05124_),
    .Z(_05649_));
 XNOR2_X2 _11154_ (.A(_05186_),
    .B(_05649_),
    .ZN(_05650_));
 NAND4_X4 _11155_ (.A1(_05636_),
    .A2(_05640_),
    .A3(_05645_),
    .A4(_05650_),
    .ZN(_05651_));
 MUX2_X1 _11156_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][52] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][52] ),
    .S(_05129_),
    .Z(_05652_));
 MUX2_X1 _11157_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][52] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][52] ),
    .S(net687),
    .Z(_05653_));
 MUX2_X1 _11158_ (.A(_05652_),
    .B(_05653_),
    .S(_05643_),
    .Z(_05654_));
 XNOR2_X2 _11159_ (.A(_05257_),
    .B(_05654_),
    .ZN(_05655_));
 MUX2_X1 _11160_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][56] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][56] ),
    .S(_05646_),
    .Z(_05656_));
 MUX2_X1 _11161_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][56] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][56] ),
    .S(_05646_),
    .Z(_05657_));
 MUX2_X1 _11162_ (.A(_05656_),
    .B(_05657_),
    .S(_05643_),
    .Z(_05658_));
 XNOR2_X2 _11163_ (.A(_05204_),
    .B(_05658_),
    .ZN(_05659_));
 MUX2_X1 _11164_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][62] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][62] ),
    .S(_05646_),
    .Z(_05660_));
 MUX2_X1 _11165_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][62] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][62] ),
    .S(_05646_),
    .Z(_05661_));
 MUX2_X1 _11166_ (.A(_05660_),
    .B(_05661_),
    .S(_05643_),
    .Z(_05662_));
 XNOR2_X2 _11167_ (.A(_05197_),
    .B(_05662_),
    .ZN(_05663_));
 MUX2_X1 _11168_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][54] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][54] ),
    .S(net668),
    .Z(_05664_));
 MUX2_X1 _11169_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][54] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][54] ),
    .S(net666),
    .Z(_05665_));
 MUX2_X1 _11170_ (.A(_05664_),
    .B(_05665_),
    .S(_05643_),
    .Z(_05666_));
 XNOR2_X2 _11171_ (.A(_05252_),
    .B(_05666_),
    .ZN(_05667_));
 NAND4_X4 _11172_ (.A1(_05655_),
    .A2(_05659_),
    .A3(_05663_),
    .A4(_05667_),
    .ZN(_05668_));
 MUX2_X1 _11173_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][57] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][57] ),
    .S(_05646_),
    .Z(_05669_));
 MUX2_X1 _11174_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][57] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][57] ),
    .S(net668),
    .Z(_05670_));
 MUX2_X1 _11175_ (.A(_05669_),
    .B(_05670_),
    .S(_05643_),
    .Z(_05671_));
 XNOR2_X2 _11176_ (.A(_05231_),
    .B(_05671_),
    .ZN(_05672_));
 MUX2_X1 _11177_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][59] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][59] ),
    .S(_05128_),
    .Z(_05673_));
 MUX2_X1 _11178_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][59] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][59] ),
    .S(net668),
    .Z(_05674_));
 MUX2_X1 _11179_ (.A(_05673_),
    .B(_05674_),
    .S(_05643_),
    .Z(_05675_));
 XNOR2_X2 _11180_ (.A(_05226_),
    .B(_05675_),
    .ZN(_05676_));
 MUX2_X1 _11181_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][61] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][61] ),
    .S(_05128_),
    .Z(_05677_));
 MUX2_X1 _11182_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][61] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][61] ),
    .S(net668),
    .Z(_05678_));
 MUX2_X1 _11183_ (.A(_05677_),
    .B(_05678_),
    .S(_05643_),
    .Z(_05679_));
 XNOR2_X2 _11184_ (.A(_05236_),
    .B(_05679_),
    .ZN(_05680_));
 MUX2_X1 _11185_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][50] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][50] ),
    .S(_05128_),
    .Z(_05681_));
 MUX2_X1 _11186_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][50] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][50] ),
    .S(net666),
    .Z(_05682_));
 MUX2_X1 _11187_ (.A(_05681_),
    .B(_05682_),
    .S(_05124_),
    .Z(_05683_));
 XNOR2_X2 _11188_ (.A(_05247_),
    .B(_05683_),
    .ZN(_05684_));
 NAND4_X4 _11189_ (.A1(_05672_),
    .A2(_05676_),
    .A3(_05680_),
    .A4(_05684_),
    .ZN(_05685_));
 MUX2_X1 _11190_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][55] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][55] ),
    .S(_05646_),
    .Z(_05686_));
 MUX2_X1 _11191_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][55] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][55] ),
    .S(_05646_),
    .Z(_05687_));
 MUX2_X1 _11192_ (.A(_05686_),
    .B(_05687_),
    .S(_05643_),
    .Z(_05688_));
 XNOR2_X1 _11193_ (.A(_05209_),
    .B(_05688_),
    .ZN(_05689_));
 MUX2_X1 _11194_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][58] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][58] ),
    .S(_05646_),
    .Z(_05690_));
 MUX2_X1 _11195_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][58] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][58] ),
    .S(_05646_),
    .Z(_05691_));
 MUX2_X1 _11196_ (.A(_05690_),
    .B(_05691_),
    .S(_05643_),
    .Z(_05692_));
 XNOR2_X1 _11197_ (.A(_05215_),
    .B(_05692_),
    .ZN(_05693_));
 NAND2_X2 _11198_ (.A1(_05689_),
    .A2(_05693_),
    .ZN(_05694_));
 NOR4_X4 _11199_ (.A1(_05668_),
    .A2(_05651_),
    .A3(_05685_),
    .A4(_05694_),
    .ZN(_05695_));
 MUX2_X2 _11200_ (.A(_05623_),
    .B(_05632_),
    .S(net748),
    .Z(_05696_));
 BUF_X2 _11201_ (.A(_00055_),
    .Z(_05697_));
 AOI21_X4 _11202_ (.A(_05610_),
    .B1(_05697_),
    .B2(_05696_),
    .ZN(net623));
 BUF_X1 rebuffer130 (.A(_00010_),
    .Z(net760));
 BUF_X8 _11204_ (.A(_00010_),
    .Z(_05699_));
 BUF_X16 _11205_ (.A(_05699_),
    .Z(_05700_));
 BUF_X1 rebuffer131 (.A(net760),
    .Z(net761));
 BUF_X16 _11207_ (.A(_05700_),
    .Z(_05702_));
 BUF_X4 _11208_ (.A(_05702_),
    .Z(_05703_));
 CLKBUF_X3 _11209_ (.A(_05703_),
    .Z(_05704_));
 MUX2_X1 _11210_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][42] ),
    .S(_05704_),
    .Z(_05705_));
 MUX2_X1 _11211_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][42] ),
    .S(_05704_),
    .Z(_05706_));
 BUF_X4 _11212_ (.A(_00009_),
    .Z(_05707_));
 BUF_X4 _11213_ (.A(_05707_),
    .Z(_05708_));
 BUF_X4 _11214_ (.A(_05708_),
    .Z(_05709_));
 BUF_X4 _11215_ (.A(_05709_),
    .Z(_05710_));
 BUF_X4 _11216_ (.A(_05710_),
    .Z(_05711_));
 MUX2_X1 _11217_ (.A(_05705_),
    .B(_05706_),
    .S(_05711_),
    .Z(_05712_));
 MUX2_X1 _11218_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][42] ),
    .S(_05704_),
    .Z(_05713_));
 MUX2_X1 _11219_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][42] ),
    .S(_05704_),
    .Z(_05714_));
 MUX2_X1 _11220_ (.A(_05713_),
    .B(_05714_),
    .S(_05711_),
    .Z(_05715_));
 BUF_X4 _11221_ (.A(_00012_),
    .Z(_05716_));
 BUF_X4 _11222_ (.A(_05716_),
    .Z(_05717_));
 INV_X4 _11223_ (.A(_05717_),
    .ZN(_05718_));
 BUF_X4 _11224_ (.A(_05718_),
    .Z(_05719_));
 BUF_X4 _11225_ (.A(_05719_),
    .Z(_05720_));
 BUF_X4 _11226_ (.A(_05720_),
    .Z(_05721_));
 MUX2_X1 _11227_ (.A(_05712_),
    .B(_05715_),
    .S(_05721_),
    .Z(_05722_));
 MUX2_X1 _11228_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][42] ),
    .S(_05704_),
    .Z(_05723_));
 BUF_X4 _11229_ (.A(_05703_),
    .Z(_05724_));
 MUX2_X1 _11230_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][42] ),
    .S(_05724_),
    .Z(_05725_));
 MUX2_X1 _11231_ (.A(_05723_),
    .B(_05725_),
    .S(_05711_),
    .Z(_05726_));
 MUX2_X1 _11232_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][42] ),
    .S(_05724_),
    .Z(_05727_));
 MUX2_X1 _11233_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][42] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][42] ),
    .S(_05724_),
    .Z(_05728_));
 BUF_X4 _11234_ (.A(_05710_),
    .Z(_05729_));
 MUX2_X1 _11235_ (.A(_05727_),
    .B(_05728_),
    .S(_05729_),
    .Z(_05730_));
 MUX2_X1 _11236_ (.A(_05726_),
    .B(_05730_),
    .S(_05721_),
    .Z(_05731_));
 BUF_X4 _11237_ (.A(_00011_),
    .Z(_05732_));
 BUF_X4 _11238_ (.A(_05732_),
    .Z(_05733_));
 BUF_X4 _11239_ (.A(_05733_),
    .Z(_05734_));
 BUF_X4 _11240_ (.A(_05734_),
    .Z(_05735_));
 BUF_X4 _11241_ (.A(_05735_),
    .Z(_05736_));
 BUF_X4 _11242_ (.A(_05736_),
    .Z(_05737_));
 BUF_X8 _11243_ (.A(_05737_),
    .Z(_05738_));
 MUX2_X2 _11244_ (.A(_05722_),
    .B(_05731_),
    .S(_05738_),
    .Z(_10372_));
 MUX2_X1 _11245_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][34] ),
    .S(_05704_),
    .Z(_05739_));
 MUX2_X1 _11246_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][34] ),
    .S(_05704_),
    .Z(_05740_));
 MUX2_X1 _11247_ (.A(_05739_),
    .B(_05740_),
    .S(_05711_),
    .Z(_05741_));
 MUX2_X1 _11248_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][34] ),
    .S(_05704_),
    .Z(_05742_));
 MUX2_X1 _11249_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][34] ),
    .S(_05704_),
    .Z(_05743_));
 MUX2_X1 _11250_ (.A(_05742_),
    .B(_05743_),
    .S(_05711_),
    .Z(_05744_));
 MUX2_X1 _11251_ (.A(_05741_),
    .B(_05744_),
    .S(_05721_),
    .Z(_05745_));
 MUX2_X1 _11252_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][34] ),
    .S(_05704_),
    .Z(_05746_));
 MUX2_X1 _11253_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][34] ),
    .S(_05724_),
    .Z(_05747_));
 MUX2_X1 _11254_ (.A(_05746_),
    .B(_05747_),
    .S(_05711_),
    .Z(_05748_));
 MUX2_X1 _11255_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][34] ),
    .S(_05724_),
    .Z(_05749_));
 MUX2_X1 _11256_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][34] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][34] ),
    .S(_05724_),
    .Z(_05750_));
 MUX2_X1 _11257_ (.A(_05749_),
    .B(_05750_),
    .S(_05729_),
    .Z(_05751_));
 MUX2_X1 _11258_ (.A(_05748_),
    .B(_05751_),
    .S(_05721_),
    .Z(_05752_));
 MUX2_X2 _11259_ (.A(_05745_),
    .B(_05752_),
    .S(_05738_),
    .Z(_10417_));
 BUF_X4 _11260_ (.A(\dynamic_node_top.north_output.control.current_route_f[1] ),
    .Z(_05753_));
 BUF_X4 _11261_ (.A(_05753_),
    .Z(_05754_));
 CLKBUF_X2 _11262_ (.A(_00056_),
    .Z(_05755_));
 CLKBUF_X3 _11263_ (.A(_05755_),
    .Z(_05756_));
 BUF_X4 _11264_ (.A(\dynamic_node_top.north_output.control.current_route_f[4] ),
    .Z(_05757_));
 MUX2_X1 _11265_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][26] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][26] ),
    .S(net711),
    .Z(_05758_));
 MUX2_X1 _11266_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][26] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][26] ),
    .S(net711),
    .Z(_05759_));
 MUX2_X2 _11267_ (.A(_05758_),
    .B(_05759_),
    .S(_05463_),
    .Z(_05760_));
 NOR2_X1 _11268_ (.A1(_05489_),
    .A2(_05760_),
    .ZN(_05761_));
 BUF_X4 _11269_ (.A(_05536_),
    .Z(_05762_));
 MUX2_X1 _11270_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][23] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][23] ),
    .S(_05762_),
    .Z(_05763_));
 MUX2_X1 _11271_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][23] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][23] ),
    .S(net711),
    .Z(_05764_));
 MUX2_X2 _11272_ (.A(_05763_),
    .B(_05764_),
    .S(_05463_),
    .Z(_05765_));
 MUX2_X1 _11273_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][25] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][25] ),
    .S(_05762_),
    .Z(_05766_));
 MUX2_X1 _11274_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][25] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][25] ),
    .S(_05762_),
    .Z(_05767_));
 MUX2_X2 _11275_ (.A(_05766_),
    .B(_05767_),
    .S(_05463_),
    .Z(_05768_));
 MUX2_X1 _11276_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][24] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][24] ),
    .S(_05762_),
    .Z(_05769_));
 MUX2_X1 _11277_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][24] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][24] ),
    .S(_05762_),
    .Z(_05770_));
 MUX2_X2 _11278_ (.A(_05769_),
    .B(_05770_),
    .S(_05463_),
    .Z(_05771_));
 NOR3_X1 _11279_ (.A1(_05765_),
    .A2(_05768_),
    .A3(_05771_),
    .ZN(_05772_));
 MUX2_X1 _11280_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][22] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][22] ),
    .S(_05762_),
    .Z(_05773_));
 MUX2_X1 _11281_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][22] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][22] ),
    .S(net711),
    .Z(_05774_));
 MUX2_X2 _11282_ (.A(_05773_),
    .B(_05774_),
    .S(_05463_),
    .Z(_05775_));
 MUX2_X1 _11283_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][29] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][29] ),
    .S(net711),
    .Z(_05776_));
 MUX2_X1 _11284_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][29] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][29] ),
    .S(_05762_),
    .Z(_05777_));
 MUX2_X2 _11285_ (.A(_05776_),
    .B(_05777_),
    .S(_05463_),
    .Z(_05778_));
 MUX2_X1 _11286_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][27] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][27] ),
    .S(_05762_),
    .Z(_05779_));
 MUX2_X1 _11287_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][27] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][27] ),
    .S(_05762_),
    .Z(_05780_));
 MUX2_X2 _11288_ (.A(_05779_),
    .B(_05780_),
    .S(_05463_),
    .Z(_05781_));
 MUX2_X1 _11289_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][28] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][28] ),
    .S(net711),
    .Z(_05782_));
 MUX2_X1 _11290_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][28] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][28] ),
    .S(_05762_),
    .Z(_05783_));
 MUX2_X2 _11291_ (.A(_05782_),
    .B(_05783_),
    .S(_05463_),
    .Z(_05784_));
 NOR4_X1 _11292_ (.A1(_05775_),
    .A2(_05778_),
    .A3(_05781_),
    .A4(_05784_),
    .ZN(_05785_));
 AND3_X1 _11293_ (.A1(_05761_),
    .A2(_05772_),
    .A3(_05785_),
    .ZN(_05786_));
 BUF_X2 _11294_ (.A(net626),
    .Z(_05787_));
 MUX2_X1 _11295_ (.A(\dynamic_node_top.east_input.control.tail_last_f ),
    .B(\dynamic_node_top.east_input.control.count_one_f ),
    .S(_05787_),
    .Z(_05788_));
 OR2_X1 _11296_ (.A1(_05786_),
    .A2(_05788_),
    .ZN(_05789_));
 MUX2_X1 _11297_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][26] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][26] ),
    .S(net738),
    .Z(_05790_));
 MUX2_X1 _11298_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][26] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][26] ),
    .S(net738),
    .Z(_05791_));
 MUX2_X2 _11299_ (.A(_05790_),
    .B(_05791_),
    .S(_05151_),
    .Z(_05792_));
 NOR2_X1 _11300_ (.A1(_05185_),
    .A2(_05792_),
    .ZN(_05793_));
 MUX2_X1 _11301_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][23] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][23] ),
    .S(net738),
    .Z(_05794_));
 MUX2_X1 _11302_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][23] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][23] ),
    .S(net738),
    .Z(_05795_));
 MUX2_X2 _11303_ (.A(_05794_),
    .B(_05795_),
    .S(_05151_),
    .Z(_05796_));
 MUX2_X1 _11304_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][24] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][24] ),
    .S(_05143_),
    .Z(_05797_));
 MUX2_X1 _11305_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][24] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][24] ),
    .S(net738),
    .Z(_05798_));
 MUX2_X2 _11306_ (.A(_05797_),
    .B(_05798_),
    .S(_05151_),
    .Z(_05799_));
 MUX2_X1 _11307_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][25] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][25] ),
    .S(net740),
    .Z(_05800_));
 MUX2_X1 _11308_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][25] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][25] ),
    .S(net740),
    .Z(_05801_));
 MUX2_X2 _11309_ (.A(_05800_),
    .B(_05801_),
    .S(_05151_),
    .Z(_05802_));
 NOR3_X2 _11310_ (.A1(_05796_),
    .A2(_05799_),
    .A3(_05802_),
    .ZN(_05803_));
 MUX2_X1 _11311_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][28] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][28] ),
    .S(net738),
    .Z(_05804_));
 MUX2_X1 _11312_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][28] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][28] ),
    .S(net738),
    .Z(_05805_));
 MUX2_X2 _11313_ (.A(_05804_),
    .B(_05805_),
    .S(_05151_),
    .Z(_05806_));
 MUX2_X1 _11314_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][27] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][27] ),
    .S(_05143_),
    .Z(_05807_));
 MUX2_X1 _11315_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][27] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][27] ),
    .S(_05143_),
    .Z(_05808_));
 MUX2_X2 _11316_ (.A(_05807_),
    .B(_05808_),
    .S(_05151_),
    .Z(_05809_));
 MUX2_X1 _11317_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][29] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][29] ),
    .S(net740),
    .Z(_05810_));
 MUX2_X1 _11318_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][29] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][29] ),
    .S(net740),
    .Z(_05811_));
 MUX2_X2 _11319_ (.A(_05810_),
    .B(_05811_),
    .S(_05151_),
    .Z(_05812_));
 MUX2_X1 _11320_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][22] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][22] ),
    .S(net740),
    .Z(_05813_));
 MUX2_X1 _11321_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][22] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][22] ),
    .S(net740),
    .Z(_05814_));
 MUX2_X2 _11322_ (.A(_05813_),
    .B(_05814_),
    .S(_05151_),
    .Z(_05815_));
 NOR4_X1 _11323_ (.A1(_05806_),
    .A2(_05809_),
    .A3(_05812_),
    .A4(_05815_),
    .ZN(_05816_));
 AND3_X1 _11324_ (.A1(_05793_),
    .A2(_05803_),
    .A3(_05816_),
    .ZN(_05817_));
 BUF_X2 _11325_ (.A(net630),
    .Z(_05818_));
 MUX2_X1 _11326_ (.A(\dynamic_node_top.west_input.control.tail_last_f ),
    .B(\dynamic_node_top.west_input.control.count_one_f ),
    .S(_05818_),
    .Z(_05819_));
 OR2_X2 _11327_ (.A1(_05817_),
    .A2(_05819_),
    .ZN(_05820_));
 CLKBUF_X3 _11328_ (.A(\dynamic_node_top.north_output.control.current_route_f[3] ),
    .Z(_05821_));
 AOI22_X2 _11329_ (.A1(_05757_),
    .A2(_05789_),
    .B1(_05820_),
    .B2(_05821_),
    .ZN(_05822_));
 BUF_X4 _11330_ (.A(\dynamic_node_top.north_output.control.current_route_f[2] ),
    .Z(_05823_));
 NOR4_X4 _11331_ (.A1(_05753_),
    .A2(_05757_),
    .A3(_05823_),
    .A4(_05821_),
    .ZN(_05824_));
 BUF_X2 _11332_ (.A(net627),
    .Z(_05825_));
 MUX2_X1 _11333_ (.A(\dynamic_node_top.north_input.control.tail_last_f ),
    .B(\dynamic_node_top.north_input.control.count_one_f ),
    .S(_05825_),
    .Z(_05826_));
 MUX2_X1 _11334_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][25] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][25] ),
    .S(_05362_),
    .Z(_05827_));
 MUX2_X1 _11335_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][25] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][25] ),
    .S(_05362_),
    .Z(_05828_));
 MUX2_X2 _11336_ (.A(_05827_),
    .B(_05828_),
    .S(_05319_),
    .Z(_05829_));
 MUX2_X1 _11337_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][26] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][26] ),
    .S(net726),
    .Z(_05830_));
 MUX2_X1 _11338_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][26] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][26] ),
    .S(_05362_),
    .Z(_05831_));
 MUX2_X2 _11339_ (.A(_05830_),
    .B(_05831_),
    .S(_05319_),
    .Z(_05832_));
 NOR3_X1 _11340_ (.A1(_05346_),
    .A2(_05829_),
    .A3(_05832_),
    .ZN(_05833_));
 MUX2_X1 _11341_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][27] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][27] ),
    .S(net726),
    .Z(_05834_));
 MUX2_X1 _11342_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][27] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][27] ),
    .S(net726),
    .Z(_05835_));
 MUX2_X2 _11343_ (.A(_05834_),
    .B(_05835_),
    .S(_05320_),
    .Z(_05836_));
 MUX2_X1 _11344_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][24] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][24] ),
    .S(_05362_),
    .Z(_05837_));
 MUX2_X1 _11345_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][24] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][24] ),
    .S(net726),
    .Z(_05838_));
 MUX2_X2 _11346_ (.A(_05837_),
    .B(_05838_),
    .S(_05319_),
    .Z(_05839_));
 NOR2_X1 _11347_ (.A1(_05836_),
    .A2(_05839_),
    .ZN(_05840_));
 MUX2_X1 _11348_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][28] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][28] ),
    .S(_05362_),
    .Z(_05841_));
 MUX2_X1 _11349_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][28] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][28] ),
    .S(_05362_),
    .Z(_05842_));
 MUX2_X2 _11350_ (.A(_05841_),
    .B(_05842_),
    .S(_05319_),
    .Z(_05843_));
 MUX2_X1 _11351_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][22] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][22] ),
    .S(_05362_),
    .Z(_05844_));
 MUX2_X1 _11352_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][22] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][22] ),
    .S(_05362_),
    .Z(_05845_));
 MUX2_X1 _11353_ (.A(_05844_),
    .B(_05845_),
    .S(_05319_),
    .Z(_05846_));
 MUX2_X1 _11354_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][23] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][23] ),
    .S(net726),
    .Z(_05847_));
 MUX2_X1 _11355_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][23] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][23] ),
    .S(net726),
    .Z(_05848_));
 MUX2_X2 _11356_ (.A(_05847_),
    .B(_05848_),
    .S(_05319_),
    .Z(_05849_));
 MUX2_X1 _11357_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][29] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][29] ),
    .S(net726),
    .Z(_05850_));
 MUX2_X1 _11358_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][29] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][29] ),
    .S(_05362_),
    .Z(_05851_));
 MUX2_X1 _11359_ (.A(_05850_),
    .B(_05851_),
    .S(_05319_),
    .Z(_05852_));
 NOR4_X1 _11360_ (.A1(_05843_),
    .A2(_05846_),
    .A3(_05849_),
    .A4(_05852_),
    .ZN(_05853_));
 AND3_X1 _11361_ (.A1(_05833_),
    .A2(_05840_),
    .A3(_05853_),
    .ZN(_05854_));
 OR2_X1 _11362_ (.A1(_05826_),
    .A2(_05854_),
    .ZN(_05855_));
 AOI21_X1 _11363_ (.A(_05824_),
    .B1(_05855_),
    .B2(_05753_),
    .ZN(_05856_));
 INV_X1 _11364_ (.A(_05823_),
    .ZN(_05857_));
 CLKBUF_X3 _11365_ (.A(net628),
    .Z(_05858_));
 INV_X1 _11366_ (.A(\dynamic_node_top.proc_input.control.tail_last_f ),
    .ZN(_05859_));
 NOR2_X1 _11367_ (.A1(_05858_),
    .A2(_05859_),
    .ZN(_05860_));
 BUF_X4 _11368_ (.A(_05717_),
    .Z(_05861_));
 MUX2_X1 _11369_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][25] ),
    .S(_05861_),
    .Z(_05862_));
 NOR2_X1 _11370_ (.A1(_05735_),
    .A2(_05862_),
    .ZN(_05863_));
 INV_X2 _11371_ (.A(_05732_),
    .ZN(_05864_));
 BUF_X4 _11372_ (.A(_05864_),
    .Z(_05865_));
 BUF_X8 _11373_ (.A(_05716_),
    .Z(_05866_));
 BUF_X4 _11374_ (.A(_05866_),
    .Z(_05867_));
 MUX2_X1 _11375_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][25] ),
    .S(_05867_),
    .Z(_05868_));
 NOR2_X1 _11376_ (.A1(_05865_),
    .A2(_05868_),
    .ZN(_05869_));
 BUF_X4 _11377_ (.A(net760),
    .Z(_05870_));
 OR2_X2 _11378_ (.A1(_05707_),
    .A2(_05870_),
    .ZN(_05871_));
 BUF_X4 _11379_ (.A(_05871_),
    .Z(_05872_));
 INV_X2 _11380_ (.A(_00009_),
    .ZN(_05873_));
 BUF_X4 _11381_ (.A(_05873_),
    .Z(_05874_));
 NAND2_X2 _11382_ (.A1(_05874_),
    .A2(_05700_),
    .ZN(_05875_));
 BUF_X8 _11383_ (.A(_05716_),
    .Z(_05876_));
 BUF_X4 _11384_ (.A(_05876_),
    .Z(_05877_));
 MUX2_X1 _11385_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][25] ),
    .S(_05877_),
    .Z(_05878_));
 NOR2_X1 _11386_ (.A1(_05734_),
    .A2(_05878_),
    .ZN(_05879_));
 MUX2_X1 _11387_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][25] ),
    .S(_05877_),
    .Z(_05880_));
 NOR2_X1 _11388_ (.A1(_05865_),
    .A2(_05880_),
    .ZN(_05881_));
 OAI33_X1 _11389_ (.A1(_05863_),
    .A2(_05869_),
    .A3(_05872_),
    .B1(_05875_),
    .B2(_05879_),
    .B3(_05881_),
    .ZN(_05882_));
 MUX2_X1 _11390_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][25] ),
    .S(_05861_),
    .Z(_05883_));
 NOR2_X1 _11391_ (.A1(_05735_),
    .A2(_05883_),
    .ZN(_05884_));
 MUX2_X1 _11392_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][25] ),
    .S(_05867_),
    .Z(_05885_));
 NOR2_X1 _11393_ (.A1(_05865_),
    .A2(_05885_),
    .ZN(_05886_));
 BUF_X4 _11394_ (.A(_05707_),
    .Z(_05887_));
 BUF_X4 _11395_ (.A(_05887_),
    .Z(_05888_));
 INV_X4 _11396_ (.A(_05870_),
    .ZN(_05889_));
 BUF_X4 _11397_ (.A(_05889_),
    .Z(_05890_));
 NAND2_X1 _11398_ (.A1(_05888_),
    .A2(_05890_),
    .ZN(_05891_));
 BUF_X4 _11399_ (.A(_05699_),
    .Z(_05892_));
 NAND2_X1 _11400_ (.A1(_05707_),
    .A2(_05892_),
    .ZN(_05893_));
 BUF_X4 _11401_ (.A(_05893_),
    .Z(_05894_));
 MUX2_X1 _11402_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][25] ),
    .S(_05877_),
    .Z(_05895_));
 NOR2_X1 _11403_ (.A1(_05734_),
    .A2(_05895_),
    .ZN(_05896_));
 BUF_X4 _11404_ (.A(_05716_),
    .Z(_05897_));
 MUX2_X1 _11405_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][25] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][25] ),
    .S(_05897_),
    .Z(_05898_));
 NOR2_X1 _11406_ (.A1(_05865_),
    .A2(_05898_),
    .ZN(_05899_));
 OAI33_X1 _11407_ (.A1(_05884_),
    .A2(_05886_),
    .A3(_05891_),
    .B1(_05894_),
    .B2(_05896_),
    .B3(_05899_),
    .ZN(_05900_));
 OR2_X2 _11408_ (.A1(_05882_),
    .A2(_05900_),
    .ZN(_05901_));
 CLKBUF_X3 _11409_ (.A(_05901_),
    .Z(_05902_));
 BUF_X4 _11410_ (.A(_05870_),
    .Z(_05903_));
 BUF_X4 _11411_ (.A(_05732_),
    .Z(_05904_));
 OR2_X2 _11412_ (.A1(_05903_),
    .A2(_05904_),
    .ZN(_05905_));
 MUX2_X1 _11413_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][26] ),
    .S(_05861_),
    .Z(_05906_));
 NOR2_X1 _11414_ (.A1(_05905_),
    .A2(_05906_),
    .ZN(_05907_));
 BUF_X4 _11415_ (.A(_05892_),
    .Z(_05908_));
 BUF_X4 _11416_ (.A(_05908_),
    .Z(_05909_));
 MUX2_X1 _11417_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][26] ),
    .S(_05877_),
    .Z(_05910_));
 NOR3_X1 _11418_ (.A1(_05909_),
    .A2(_05865_),
    .A3(_05910_),
    .ZN(_05911_));
 MUX2_X1 _11419_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][26] ),
    .S(_05897_),
    .Z(_05912_));
 NOR3_X1 _11420_ (.A1(_05890_),
    .A2(_05734_),
    .A3(_05912_),
    .ZN(_05913_));
 BUF_X4 _11421_ (.A(_05732_),
    .Z(_05914_));
 NAND2_X2 _11422_ (.A1(_05903_),
    .A2(_05914_),
    .ZN(_05915_));
 MUX2_X1 _11423_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][26] ),
    .S(_05877_),
    .Z(_05916_));
 NOR2_X1 _11424_ (.A1(_05915_),
    .A2(_05916_),
    .ZN(_05917_));
 OR4_X4 _11425_ (.A1(_05907_),
    .A2(_05911_),
    .A3(_05913_),
    .A4(_05917_),
    .ZN(_05918_));
 OAI21_X4 _11426_ (.A(\dynamic_node_top.proc_input.control.header_last_temp ),
    .B1(_05181_),
    .B2(\dynamic_node_top.proc_input.NIB.elements_in_array_f[1] ),
    .ZN(_05919_));
 NOR2_X2 _11427_ (.A1(_05709_),
    .A2(_05919_),
    .ZN(_05920_));
 BUF_X4 _11428_ (.A(_05873_),
    .Z(_05921_));
 BUF_X4 _11429_ (.A(_05921_),
    .Z(_05922_));
 NOR2_X1 _11430_ (.A1(_05922_),
    .A2(_05919_),
    .ZN(_05923_));
 MUX2_X1 _11431_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][26] ),
    .S(_05867_),
    .Z(_05924_));
 NOR2_X1 _11432_ (.A1(_05924_),
    .A2(_05905_),
    .ZN(_05925_));
 MUX2_X1 _11433_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][26] ),
    .S(_05897_),
    .Z(_05926_));
 NOR3_X1 _11434_ (.A1(_05700_),
    .A2(_05864_),
    .A3(_05926_),
    .ZN(_05927_));
 MUX2_X1 _11435_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][26] ),
    .S(_05717_),
    .Z(_05928_));
 NOR3_X1 _11436_ (.A1(_05889_),
    .A2(_05734_),
    .A3(_05928_),
    .ZN(_05929_));
 MUX2_X1 _11437_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][26] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][26] ),
    .S(_05897_),
    .Z(_05930_));
 NOR2_X1 _11438_ (.A1(_05930_),
    .A2(_05915_),
    .ZN(_05931_));
 OR4_X4 _11439_ (.A1(_05925_),
    .A2(_05927_),
    .A3(_05929_),
    .A4(_05931_),
    .ZN(_05932_));
 AOI22_X4 _11440_ (.A1(_05918_),
    .A2(_05920_),
    .B1(_05923_),
    .B2(_05932_),
    .ZN(_05933_));
 NOR2_X4 _11441_ (.A1(_05702_),
    .A2(_05719_),
    .ZN(_05934_));
 BUF_X4 _11442_ (.A(_05732_),
    .Z(_05935_));
 MUX2_X1 _11443_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][24] ),
    .S(_05935_),
    .Z(_05936_));
 MUX2_X1 _11444_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][24] ),
    .S(_05935_),
    .Z(_05937_));
 BUF_X4 _11445_ (.A(_05887_),
    .Z(_05938_));
 MUX2_X1 _11446_ (.A(_05936_),
    .B(_05937_),
    .S(_05938_),
    .Z(_05939_));
 MUX2_X1 _11447_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[4][24] ),
    .S(_05904_),
    .Z(_05940_));
 MUX2_X1 _11448_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][24] ),
    .S(_05914_),
    .Z(_05941_));
 MUX2_X1 _11449_ (.A(_05940_),
    .B(_05941_),
    .S(_05888_),
    .Z(_05942_));
 BUF_X4 _11450_ (.A(_05877_),
    .Z(_05943_));
 NOR2_X4 _11451_ (.A1(_05702_),
    .A2(_05943_),
    .ZN(_05944_));
 AOI22_X2 _11452_ (.A1(_05934_),
    .A2(_05939_),
    .B1(_05942_),
    .B2(_05944_),
    .ZN(_05945_));
 BUF_X4 _11453_ (.A(_05889_),
    .Z(_05946_));
 NOR2_X4 _11454_ (.A1(_05946_),
    .A2(_05719_),
    .ZN(_05947_));
 MUX2_X1 _11455_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][24] ),
    .S(_05914_),
    .Z(_05948_));
 MUX2_X1 _11456_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][24] ),
    .S(_05914_),
    .Z(_05949_));
 MUX2_X1 _11457_ (.A(_05948_),
    .B(_05949_),
    .S(_05938_),
    .Z(_05950_));
 MUX2_X1 _11458_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][24] ),
    .S(_05904_),
    .Z(_05951_));
 MUX2_X1 _11459_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][24] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][24] ),
    .S(_05904_),
    .Z(_05952_));
 MUX2_X1 _11460_ (.A(_05951_),
    .B(_05952_),
    .S(_05888_),
    .Z(_05953_));
 NOR2_X4 _11461_ (.A1(_05946_),
    .A2(_05943_),
    .ZN(_05954_));
 AOI22_X2 _11462_ (.A1(_05947_),
    .A2(_05950_),
    .B1(_05953_),
    .B2(_05954_),
    .ZN(_05955_));
 NAND2_X4 _11463_ (.A1(_05945_),
    .A2(_05955_),
    .ZN(_05956_));
 MUX2_X1 _11464_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][27] ),
    .S(_05935_),
    .Z(_05957_));
 MUX2_X1 _11465_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][27] ),
    .S(_05935_),
    .Z(_05958_));
 MUX2_X1 _11466_ (.A(_05957_),
    .B(_05958_),
    .S(_05938_),
    .Z(_05959_));
 MUX2_X1 _11467_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[4][27] ),
    .S(_05904_),
    .Z(_05960_));
 MUX2_X1 _11468_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][27] ),
    .S(_05904_),
    .Z(_05961_));
 MUX2_X1 _11469_ (.A(_05960_),
    .B(_05961_),
    .S(_05888_),
    .Z(_05962_));
 AOI22_X2 _11470_ (.A1(_05934_),
    .A2(_05959_),
    .B1(_05962_),
    .B2(_05944_),
    .ZN(_05963_));
 MUX2_X1 _11471_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][27] ),
    .S(_05914_),
    .Z(_05964_));
 MUX2_X1 _11472_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][27] ),
    .S(_05914_),
    .Z(_05965_));
 MUX2_X1 _11473_ (.A(_05964_),
    .B(_05965_),
    .S(_05888_),
    .Z(_05966_));
 BUF_X4 _11474_ (.A(_05732_),
    .Z(_05967_));
 MUX2_X1 _11475_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][27] ),
    .S(_05967_),
    .Z(_05968_));
 MUX2_X1 _11476_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][27] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][27] ),
    .S(_05967_),
    .Z(_05969_));
 MUX2_X1 _11477_ (.A(_05968_),
    .B(_05969_),
    .S(_05888_),
    .Z(_05970_));
 AOI22_X2 _11478_ (.A1(_05947_),
    .A2(_05966_),
    .B1(_05970_),
    .B2(_05954_),
    .ZN(_05971_));
 NAND2_X4 _11479_ (.A1(_05963_),
    .A2(_05971_),
    .ZN(_05972_));
 NOR4_X2 _11480_ (.A1(_05902_),
    .A2(_05933_),
    .A3(_05956_),
    .A4(_05972_),
    .ZN(_05973_));
 MUX2_X1 _11481_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][29] ),
    .S(_05700_),
    .Z(_05974_));
 MUX2_X1 _11482_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][29] ),
    .S(_05700_),
    .Z(_05975_));
 MUX2_X2 _11483_ (.A(_05974_),
    .B(_05975_),
    .S(_05708_),
    .Z(_05976_));
 BUF_X4 _11484_ (.A(_05864_),
    .Z(_05977_));
 NAND2_X1 _11485_ (.A1(_05977_),
    .A2(_05718_),
    .ZN(_05978_));
 NAND2_X2 _11486_ (.A1(_05734_),
    .A2(_05718_),
    .ZN(_05979_));
 MUX2_X1 _11487_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][29] ),
    .S(_05892_),
    .Z(_05980_));
 MUX2_X1 _11488_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][29] ),
    .S(_05892_),
    .Z(_05981_));
 MUX2_X2 _11489_ (.A(_05980_),
    .B(_05981_),
    .S(_05708_),
    .Z(_05982_));
 OAI22_X4 _11490_ (.A1(_05976_),
    .A2(_05978_),
    .B1(_05979_),
    .B2(_05982_),
    .ZN(_05983_));
 MUX2_X1 _11491_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][29] ),
    .S(_05733_),
    .Z(_05984_));
 MUX2_X1 _11492_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][29] ),
    .S(_05733_),
    .Z(_05985_));
 MUX2_X1 _11493_ (.A(_05984_),
    .B(_05985_),
    .S(_05708_),
    .Z(_05986_));
 NAND2_X1 _11494_ (.A1(_05946_),
    .A2(_05943_),
    .ZN(_05987_));
 NAND2_X1 _11495_ (.A1(_05909_),
    .A2(_05943_),
    .ZN(_05988_));
 MUX2_X1 _11496_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][29] ),
    .S(_05732_),
    .Z(_05989_));
 MUX2_X1 _11497_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][29] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][29] ),
    .S(_05732_),
    .Z(_05990_));
 MUX2_X1 _11498_ (.A(_05989_),
    .B(_05990_),
    .S(_05887_),
    .Z(_05991_));
 OAI22_X4 _11499_ (.A1(_05986_),
    .A2(_05987_),
    .B1(_05988_),
    .B2(_05991_),
    .ZN(_05992_));
 NOR2_X4 _11500_ (.A1(_05983_),
    .A2(_05992_),
    .ZN(_05993_));
 MUX2_X1 _11501_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][28] ),
    .S(_05935_),
    .Z(_05994_));
 MUX2_X1 _11502_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][28] ),
    .S(_05935_),
    .Z(_05995_));
 MUX2_X1 _11503_ (.A(_05994_),
    .B(_05995_),
    .S(_05938_),
    .Z(_05996_));
 MUX2_X1 _11504_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[4][28] ),
    .S(_05904_),
    .Z(_05997_));
 MUX2_X1 _11505_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][28] ),
    .S(_05904_),
    .Z(_05998_));
 MUX2_X1 _11506_ (.A(_05997_),
    .B(_05998_),
    .S(_05888_),
    .Z(_05999_));
 AOI22_X4 _11507_ (.A1(_05934_),
    .A2(_05996_),
    .B1(_05999_),
    .B2(_05944_),
    .ZN(_06000_));
 MUX2_X1 _11508_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][28] ),
    .S(_05914_),
    .Z(_06001_));
 MUX2_X1 _11509_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][28] ),
    .S(_05914_),
    .Z(_06002_));
 MUX2_X1 _11510_ (.A(_06001_),
    .B(_06002_),
    .S(_05938_),
    .Z(_06003_));
 MUX2_X1 _11511_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][28] ),
    .S(_05904_),
    .Z(_06004_));
 MUX2_X1 _11512_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][28] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][28] ),
    .S(_05904_),
    .Z(_06005_));
 MUX2_X2 _11513_ (.A(_06004_),
    .B(_06005_),
    .S(_05888_),
    .Z(_06006_));
 AOI22_X4 _11514_ (.A1(_05947_),
    .A2(_06003_),
    .B1(_06006_),
    .B2(_05954_),
    .ZN(_06007_));
 NAND2_X4 _11515_ (.A1(_06000_),
    .A2(_06007_),
    .ZN(_06008_));
 CLKBUF_X3 _11516_ (.A(_05943_),
    .Z(_06009_));
 MUX2_X1 _11517_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[4][23] ),
    .S(_05935_),
    .Z(_06010_));
 NOR2_X1 _11518_ (.A1(_05872_),
    .A2(_06010_),
    .ZN(_06011_));
 MUX2_X1 _11519_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][23] ),
    .S(_05733_),
    .Z(_06012_));
 NOR3_X2 _11520_ (.A1(_05938_),
    .A2(_05890_),
    .A3(_06012_),
    .ZN(_06013_));
 MUX2_X1 _11521_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][23] ),
    .S(_05733_),
    .Z(_06014_));
 NOR3_X2 _11522_ (.A1(_05874_),
    .A2(_05700_),
    .A3(_06014_),
    .ZN(_06015_));
 MUX2_X1 _11523_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][23] ),
    .S(_05967_),
    .Z(_06016_));
 NOR2_X1 _11524_ (.A1(_05894_),
    .A2(_06016_),
    .ZN(_06017_));
 NOR4_X4 _11525_ (.A1(_06011_),
    .A2(_06013_),
    .A3(_06015_),
    .A4(_06017_),
    .ZN(_06018_));
 MUX2_X1 _11526_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[4][22] ),
    .S(_05935_),
    .Z(_06019_));
 NOR2_X1 _11527_ (.A1(_05872_),
    .A2(_06019_),
    .ZN(_06020_));
 MUX2_X1 _11528_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][22] ),
    .S(_05733_),
    .Z(_06021_));
 NOR3_X2 _11529_ (.A1(_05888_),
    .A2(_05890_),
    .A3(_06021_),
    .ZN(_06022_));
 MUX2_X1 _11530_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][22] ),
    .S(_05732_),
    .Z(_06023_));
 NOR3_X2 _11531_ (.A1(_05874_),
    .A2(_05700_),
    .A3(_06023_),
    .ZN(_06024_));
 MUX2_X1 _11532_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][22] ),
    .S(_05733_),
    .Z(_06025_));
 NOR2_X1 _11533_ (.A1(_05894_),
    .A2(_06025_),
    .ZN(_06026_));
 NOR4_X4 _11534_ (.A1(_06020_),
    .A2(_06022_),
    .A3(_06024_),
    .A4(_06026_),
    .ZN(_06027_));
 OR3_X1 _11535_ (.A1(_06009_),
    .A2(_06018_),
    .A3(_06027_),
    .ZN(_06028_));
 MUX2_X1 _11536_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][23] ),
    .S(_05734_),
    .Z(_06029_));
 NOR2_X1 _11537_ (.A1(_05872_),
    .A2(_06029_),
    .ZN(_06030_));
 BUF_X4 _11538_ (.A(_05887_),
    .Z(_06031_));
 MUX2_X1 _11539_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][23] ),
    .S(_05967_),
    .Z(_06032_));
 NOR3_X1 _11540_ (.A1(_06031_),
    .A2(_05946_),
    .A3(_06032_),
    .ZN(_06033_));
 MUX2_X1 _11541_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][23] ),
    .S(_05733_),
    .Z(_06034_));
 NOR3_X1 _11542_ (.A1(_05922_),
    .A2(_05909_),
    .A3(_06034_),
    .ZN(_06035_));
 MUX2_X1 _11543_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][23] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][23] ),
    .S(_05967_),
    .Z(_06036_));
 NOR2_X1 _11544_ (.A1(_05894_),
    .A2(_06036_),
    .ZN(_06037_));
 OR4_X4 _11545_ (.A1(_06030_),
    .A2(_06033_),
    .A3(_06035_),
    .A4(_06037_),
    .ZN(_06038_));
 MUX2_X1 _11546_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][22] ),
    .S(_05734_),
    .Z(_06039_));
 NOR2_X1 _11547_ (.A1(_05872_),
    .A2(_06039_),
    .ZN(_06040_));
 MUX2_X1 _11548_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][22] ),
    .S(_05967_),
    .Z(_06041_));
 NOR3_X1 _11549_ (.A1(_06031_),
    .A2(_05890_),
    .A3(_06041_),
    .ZN(_06042_));
 MUX2_X1 _11550_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][22] ),
    .S(_05733_),
    .Z(_06043_));
 NOR3_X1 _11551_ (.A1(_05922_),
    .A2(_05909_),
    .A3(_06043_),
    .ZN(_06044_));
 MUX2_X1 _11552_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][22] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][22] ),
    .S(_05967_),
    .Z(_06045_));
 NOR2_X1 _11553_ (.A1(_05894_),
    .A2(_06045_),
    .ZN(_06046_));
 OR4_X4 _11554_ (.A1(_06040_),
    .A2(_06042_),
    .A3(_06044_),
    .A4(_06046_),
    .ZN(_06047_));
 NAND3_X1 _11555_ (.A1(_06009_),
    .A2(_06038_),
    .A3(_06047_),
    .ZN(_06048_));
 AOI211_X2 _11556_ (.A(_05993_),
    .B(_06008_),
    .C1(_06028_),
    .C2(_06048_),
    .ZN(_06049_));
 AOI221_X2 _11557_ (.A(_05860_),
    .B1(_05973_),
    .B2(_06049_),
    .C1(_05858_),
    .C2(\dynamic_node_top.proc_input.control.count_one_f ),
    .ZN(_06050_));
 OAI211_X2 _11558_ (.A(_05822_),
    .B(_05856_),
    .C1(_05857_),
    .C2(_06050_),
    .ZN(_06051_));
 BUF_X2 _11559_ (.A(net629),
    .Z(_06052_));
 MUX2_X1 _11560_ (.A(\dynamic_node_top.south_input.control.tail_last_f ),
    .B(\dynamic_node_top.south_input.control.count_one_f ),
    .S(_06052_),
    .Z(_06053_));
 MUX2_X1 _11561_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][26] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][26] ),
    .S(net746),
    .Z(_06054_));
 MUX2_X1 _11562_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][26] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][26] ),
    .S(net746),
    .Z(_06055_));
 MUX2_X2 _11563_ (.A(_06054_),
    .B(_06055_),
    .S(_05126_),
    .Z(_06056_));
 OR2_X1 _11564_ (.A1(_05618_),
    .A2(_06056_),
    .ZN(_06057_));
 MUX2_X1 _11565_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][23] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][23] ),
    .S(net746),
    .Z(_06058_));
 MUX2_X1 _11566_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][23] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][23] ),
    .S(net746),
    .Z(_06059_));
 MUX2_X2 _11567_ (.A(_06058_),
    .B(_06059_),
    .S(_05126_),
    .Z(_06060_));
 BUF_X8 _11568_ (.A(net746),
    .Z(_06061_));
 MUX2_X1 _11569_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][24] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][24] ),
    .S(_06061_),
    .Z(_06062_));
 MUX2_X1 _11570_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][24] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][24] ),
    .S(_06061_),
    .Z(_06063_));
 MUX2_X2 _11571_ (.A(_06062_),
    .B(_06063_),
    .S(_05126_),
    .Z(_06064_));
 MUX2_X1 _11572_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][25] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][25] ),
    .S(_06061_),
    .Z(_06065_));
 MUX2_X1 _11573_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][25] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][25] ),
    .S(_06061_),
    .Z(_06066_));
 MUX2_X2 _11574_ (.A(_06065_),
    .B(_06066_),
    .S(_05124_),
    .Z(_06067_));
 OR3_X1 _11575_ (.A1(_06060_),
    .A2(_06064_),
    .A3(_06067_),
    .ZN(_06068_));
 MUX2_X1 _11576_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][29] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][29] ),
    .S(_06061_),
    .Z(_06069_));
 MUX2_X1 _11577_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][29] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][29] ),
    .S(_06061_),
    .Z(_06070_));
 MUX2_X2 _11578_ (.A(_06069_),
    .B(_06070_),
    .S(_05124_),
    .Z(_06071_));
 MUX2_X1 _11579_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][27] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][27] ),
    .S(_06061_),
    .Z(_06072_));
 MUX2_X1 _11580_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][27] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][27] ),
    .S(_06061_),
    .Z(_06073_));
 MUX2_X2 _11581_ (.A(_06072_),
    .B(_06073_),
    .S(_05124_),
    .Z(_06074_));
 MUX2_X1 _11582_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][28] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][28] ),
    .S(_06061_),
    .Z(_06075_));
 MUX2_X1 _11583_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][28] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][28] ),
    .S(_06061_),
    .Z(_06076_));
 MUX2_X2 _11584_ (.A(_06075_),
    .B(_06076_),
    .S(_05124_),
    .Z(_06077_));
 MUX2_X1 _11585_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][22] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][22] ),
    .S(net746),
    .Z(_06078_));
 MUX2_X1 _11586_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][22] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][22] ),
    .S(net746),
    .Z(_06079_));
 MUX2_X2 _11587_ (.A(_06078_),
    .B(_06079_),
    .S(_05124_),
    .Z(_06080_));
 OR4_X2 _11588_ (.A1(_06071_),
    .A2(_06074_),
    .A3(_06077_),
    .A4(_06080_),
    .ZN(_06081_));
 NOR3_X2 _11589_ (.A1(_06057_),
    .A2(_06068_),
    .A3(_06081_),
    .ZN(_06082_));
 NOR2_X2 _11590_ (.A1(_06053_),
    .A2(_06082_),
    .ZN(_06083_));
 NAND2_X1 _11591_ (.A1(_05824_),
    .A2(_06083_),
    .ZN(_06084_));
 BUF_X4 _11592_ (.A(_00042_),
    .Z(_06085_));
 AND2_X2 _11593_ (.A1(_06085_),
    .A2(_05824_),
    .ZN(_06086_));
 INV_X1 _11594_ (.A(\dynamic_node_top.north_output.space.is_one_f ),
    .ZN(_06087_));
 NOR2_X1 _11595_ (.A1(_06087_),
    .A2(\dynamic_node_top.north_output.space.valid_f ),
    .ZN(_06088_));
 NOR3_X1 _11596_ (.A1(\dynamic_node_top.north_output.space.is_two_or_more_f ),
    .A2(\dynamic_node_top.north_output.space.yummy_f ),
    .A3(_06088_),
    .ZN(_06089_));
 CLKBUF_X2 _11597_ (.A(\dynamic_node_top.north_output.control.current_route_f[0] ),
    .Z(_06090_));
 AOI22_X1 _11598_ (.A1(_05753_),
    .A2(_05168_),
    .B1(_05170_),
    .B2(_06090_),
    .ZN(_06091_));
 AOI22_X1 _11599_ (.A1(_05821_),
    .A2(_05175_),
    .B1(_05177_),
    .B2(_05757_),
    .ZN(_06092_));
 NAND2_X1 _11600_ (.A1(_06091_),
    .A2(_06092_),
    .ZN(_06093_));
 AOI21_X1 _11601_ (.A(_06093_),
    .B1(_05182_),
    .B2(_05823_),
    .ZN(_06094_));
 OR3_X2 _11602_ (.A1(_06086_),
    .A2(_06089_),
    .A3(_06094_),
    .ZN(_06095_));
 CLKBUF_X3 _11603_ (.A(_05618_),
    .Z(_06096_));
 NOR2_X1 _11604_ (.A1(_05382_),
    .A2(_06096_),
    .ZN(_06097_));
 INV_X2 _11605_ (.A(_05613_),
    .ZN(_06098_));
 INV_X2 _11606_ (.A(_05616_),
    .ZN(_06099_));
 CLKBUF_X3 _11607_ (.A(_05621_),
    .Z(_06100_));
 NOR3_X1 _11608_ (.A1(_06098_),
    .A2(_06099_),
    .A3(_06100_),
    .ZN(_06101_));
 OAI21_X1 _11609_ (.A(_06097_),
    .B1(_06101_),
    .B2(_05383_),
    .ZN(_06102_));
 AND2_X2 _11610_ (.A1(\dynamic_node_top.south_input.control.header_last_temp ),
    .A2(_05170_),
    .ZN(_06103_));
 AND2_X4 _11611_ (.A1(_06103_),
    .A2(_05630_),
    .ZN(_06104_));
 OR2_X4 _11612_ (.A1(_05625_),
    .A2(_05626_),
    .ZN(_06105_));
 AOI21_X1 _11613_ (.A(_10204_),
    .B1(_10207_),
    .B2(net657),
    .ZN(_06106_));
 NAND2_X4 _11614_ (.A1(_06105_),
    .A2(_06106_),
    .ZN(_06107_));
 NOR3_X1 _11615_ (.A1(_10213_),
    .A2(_10210_),
    .A3(_10216_),
    .ZN(_06108_));
 OAI21_X1 _11616_ (.A(_10217_),
    .B1(_10220_),
    .B2(_10219_),
    .ZN(_06109_));
 OR2_X1 _11617_ (.A1(_10219_),
    .A2(_10222_),
    .ZN(_06110_));
 INV_X1 _11618_ (.A(_10226_),
    .ZN(_06111_));
 AOI21_X1 _11619_ (.A(_06110_),
    .B1(_06111_),
    .B2(_10223_),
    .ZN(_06112_));
 OAI21_X2 _11620_ (.A(_06108_),
    .B1(_06109_),
    .B2(_06112_),
    .ZN(_06113_));
 NAND2_X1 _11621_ (.A1(_10208_),
    .A2(_10205_),
    .ZN(_06114_));
 OAI21_X1 _11622_ (.A(_10211_),
    .B1(_10214_),
    .B2(_10213_),
    .ZN(_06115_));
 INV_X1 _11623_ (.A(_10210_),
    .ZN(_06116_));
 AOI21_X2 _11624_ (.A(_06114_),
    .B1(_06115_),
    .B2(_06116_),
    .ZN(_06117_));
 AND2_X2 _11625_ (.A1(_06113_),
    .A2(_06117_),
    .ZN(_06118_));
 OAI221_X2 _11626_ (.A(_06104_),
    .B1(_06107_),
    .B2(_06118_),
    .C1(_06105_),
    .C2(_06101_),
    .ZN(_06119_));
 MUX2_X2 _11627_ (.A(_06102_),
    .B(_06119_),
    .S(net747),
    .Z(_06120_));
 BUF_X1 rebuffer37 (.A(_10302_),
    .Z(net691));
 BUF_X2 _11629_ (.A(_00043_),
    .Z(_06122_));
 AOI21_X4 _11630_ (.A(_06095_),
    .B1(_06120_),
    .B2(_06122_),
    .ZN(net622));
 NAND3_X1 _11631_ (.A1(_06051_),
    .A2(_06084_),
    .A3(net622),
    .ZN(_06123_));
 CLKBUF_X2 _11632_ (.A(\dynamic_node_top.north_output.control.planned_f ),
    .Z(_06124_));
 OR2_X1 _11633_ (.A1(_06124_),
    .A2(net622),
    .ZN(_06125_));
 AND2_X1 _11634_ (.A1(_06123_),
    .A2(_06125_),
    .ZN(_06126_));
 BUF_X2 _11635_ (.A(_06126_),
    .Z(_06127_));
 NAND3_X1 _11636_ (.A1(_05754_),
    .A2(_05756_),
    .A3(_06127_),
    .ZN(_06128_));
 BUF_X4 _11637_ (.A(_05699_),
    .Z(_06129_));
 CLKBUF_X3 _11638_ (.A(_06129_),
    .Z(_06130_));
 MUX2_X1 _11639_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][31] ),
    .S(_06130_),
    .Z(_06131_));
 MUX2_X1 _11640_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][31] ),
    .S(_06130_),
    .Z(_06132_));
 MUX2_X1 _11641_ (.A(_06131_),
    .B(_06132_),
    .S(_05709_),
    .Z(_06133_));
 MUX2_X1 _11642_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][31] ),
    .S(_06130_),
    .Z(_06134_));
 MUX2_X1 _11643_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][31] ),
    .S(_06130_),
    .Z(_06135_));
 MUX2_X1 _11644_ (.A(_06134_),
    .B(_06135_),
    .S(_05709_),
    .Z(_06136_));
 MUX2_X1 _11645_ (.A(_06133_),
    .B(_06136_),
    .S(_05719_),
    .Z(_06137_));
 MUX2_X1 _11646_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][31] ),
    .S(_06130_),
    .Z(_06138_));
 MUX2_X1 _11647_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][31] ),
    .S(_06130_),
    .Z(_06139_));
 MUX2_X1 _11648_ (.A(_06138_),
    .B(_06139_),
    .S(_05709_),
    .Z(_06140_));
 MUX2_X1 _11649_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][31] ),
    .S(_05700_),
    .Z(_06141_));
 MUX2_X1 _11650_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][31] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][31] ),
    .S(_05700_),
    .Z(_06142_));
 MUX2_X1 _11651_ (.A(_06141_),
    .B(_06142_),
    .S(_05709_),
    .Z(_06143_));
 MUX2_X1 _11652_ (.A(_06140_),
    .B(_06143_),
    .S(_05720_),
    .Z(_06144_));
 MUX2_X1 _11653_ (.A(_06137_),
    .B(_06144_),
    .S(_05736_),
    .Z(_06145_));
 CLKBUF_X3 _11654_ (.A(_06145_),
    .Z(_06146_));
 OR2_X1 _11655_ (.A1(_05919_),
    .A2(_06146_),
    .ZN(_06147_));
 MUX2_X1 _11656_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][32] ),
    .S(_05903_),
    .Z(_06148_));
 MUX2_X1 _11657_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][32] ),
    .S(_05903_),
    .Z(_06149_));
 MUX2_X1 _11658_ (.A(_06148_),
    .B(_06149_),
    .S(_05938_),
    .Z(_06150_));
 MUX2_X1 _11659_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][32] ),
    .S(_05903_),
    .Z(_06151_));
 MUX2_X1 _11660_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][32] ),
    .S(_05903_),
    .Z(_06152_));
 MUX2_X1 _11661_ (.A(_06151_),
    .B(_06152_),
    .S(_05938_),
    .Z(_06153_));
 MUX2_X1 _11662_ (.A(_06150_),
    .B(_06153_),
    .S(_05719_),
    .Z(_06154_));
 MUX2_X1 _11663_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][32] ),
    .S(_05903_),
    .Z(_06155_));
 MUX2_X1 _11664_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][32] ),
    .S(_05908_),
    .Z(_06156_));
 MUX2_X1 _11665_ (.A(_06155_),
    .B(_06156_),
    .S(_05938_),
    .Z(_06157_));
 MUX2_X1 _11666_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][32] ),
    .S(_05908_),
    .Z(_06158_));
 MUX2_X1 _11667_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][32] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][32] ),
    .S(_05908_),
    .Z(_06159_));
 MUX2_X1 _11668_ (.A(_06158_),
    .B(_06159_),
    .S(_06031_),
    .Z(_06160_));
 MUX2_X1 _11669_ (.A(_06157_),
    .B(_06160_),
    .S(_05719_),
    .Z(_06161_));
 MUX2_X2 _11670_ (.A(_06154_),
    .B(_06161_),
    .S(_05736_),
    .Z(_06162_));
 BUF_X4 _11671_ (.A(_06162_),
    .Z(_06163_));
 MUX2_X1 _11672_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][30] ),
    .S(_05908_),
    .Z(_06164_));
 MUX2_X1 _11673_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][30] ),
    .S(_05908_),
    .Z(_06165_));
 MUX2_X1 _11674_ (.A(_06164_),
    .B(_06165_),
    .S(_06031_),
    .Z(_06166_));
 MUX2_X1 _11675_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][30] ),
    .S(_05908_),
    .Z(_06167_));
 MUX2_X1 _11676_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][30] ),
    .S(_06130_),
    .Z(_06168_));
 MUX2_X1 _11677_ (.A(_06167_),
    .B(_06168_),
    .S(_06031_),
    .Z(_06169_));
 MUX2_X1 _11678_ (.A(_06166_),
    .B(_06169_),
    .S(_05719_),
    .Z(_06170_));
 MUX2_X1 _11679_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][30] ),
    .S(_05908_),
    .Z(_06171_));
 MUX2_X1 _11680_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][30] ),
    .S(_06130_),
    .Z(_06172_));
 MUX2_X1 _11681_ (.A(_06171_),
    .B(_06172_),
    .S(_06031_),
    .Z(_06173_));
 MUX2_X1 _11682_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][30] ),
    .S(_06130_),
    .Z(_06174_));
 MUX2_X1 _11683_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][30] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][30] ),
    .S(_06130_),
    .Z(_06175_));
 MUX2_X1 _11684_ (.A(_06174_),
    .B(_06175_),
    .S(_06031_),
    .Z(_06176_));
 MUX2_X1 _11685_ (.A(_06173_),
    .B(_06176_),
    .S(_05719_),
    .Z(_06177_));
 MUX2_X2 _11686_ (.A(_06170_),
    .B(_06177_),
    .S(_05736_),
    .Z(_06178_));
 BUF_X4 _11687_ (.A(_06178_),
    .Z(_06179_));
 NAND2_X1 _11688_ (.A1(_06163_),
    .A2(_06179_),
    .ZN(_06180_));
 OR3_X1 _11689_ (.A1(_05383_),
    .A2(_06147_),
    .A3(_06180_),
    .ZN(_06181_));
 AND2_X1 _11690_ (.A1(\dynamic_node_top.proc_input.control.header_last_temp ),
    .A2(_05182_),
    .ZN(_06182_));
 CLKBUF_X3 _11691_ (.A(_06182_),
    .Z(_06183_));
 NAND2_X1 _11692_ (.A1(_05383_),
    .A2(_06183_),
    .ZN(_06184_));
 AOI21_X1 _11693_ (.A(_05382_),
    .B1(_06181_),
    .B2(_06184_),
    .ZN(_06185_));
 NAND4_X2 _11694_ (.A1(_10386_),
    .A2(_10395_),
    .A3(_10392_),
    .A4(_10389_),
    .ZN(_06186_));
 NAND4_X1 _11695_ (.A1(_10380_),
    .A2(_10374_),
    .A3(_10377_),
    .A4(_10383_),
    .ZN(_06187_));
 OR2_X1 _11696_ (.A1(_06186_),
    .A2(_06187_),
    .ZN(_06188_));
 NAND4_X2 _11697_ (.A1(_10398_),
    .A2(_10401_),
    .A3(_10404_),
    .A4(_10407_),
    .ZN(_06189_));
 NAND4_X1 _11698_ (.A1(_10410_),
    .A2(_10413_),
    .A3(_10416_),
    .A4(_10419_),
    .ZN(_06190_));
 OR2_X2 _11699_ (.A1(_06189_),
    .A2(_06190_),
    .ZN(_06191_));
 OR3_X1 _11700_ (.A1(_06147_),
    .A2(_06180_),
    .A3(_06191_),
    .ZN(_06192_));
 INV_X1 _11701_ (.A(_10400_),
    .ZN(_06193_));
 AOI21_X1 _11702_ (.A(_10403_),
    .B1(_10404_),
    .B2(_10406_),
    .ZN(_06194_));
 INV_X1 _11703_ (.A(_10401_),
    .ZN(_06195_));
 OAI21_X1 _11704_ (.A(_06193_),
    .B1(_06194_),
    .B2(_06195_),
    .ZN(_06196_));
 AOI21_X1 _11705_ (.A(_10397_),
    .B1(_06196_),
    .B2(_10398_),
    .ZN(_06197_));
 INV_X1 _11706_ (.A(_10412_),
    .ZN(_06198_));
 INV_X1 _11707_ (.A(_10418_),
    .ZN(_06199_));
 AOI21_X1 _11708_ (.A(_10415_),
    .B1(_06199_),
    .B2(_10416_),
    .ZN(_06200_));
 INV_X1 _11709_ (.A(_10413_),
    .ZN(_06201_));
 OAI21_X1 _11710_ (.A(_06198_),
    .B1(_06200_),
    .B2(_06201_),
    .ZN(_06202_));
 AOI21_X1 _11711_ (.A(_10409_),
    .B1(_06202_),
    .B2(_10410_),
    .ZN(_06203_));
 OAI21_X2 _11712_ (.A(_06197_),
    .B1(_06203_),
    .B2(_06189_),
    .ZN(_06204_));
 NAND3_X1 _11713_ (.A1(_06182_),
    .A2(_06191_),
    .A3(_06204_),
    .ZN(_06205_));
 AOI21_X1 _11714_ (.A(_06188_),
    .B1(_06192_),
    .B2(_06205_),
    .ZN(_06206_));
 NAND2_X4 _11715_ (.A1(_05707_),
    .A2(_05877_),
    .ZN(_06207_));
 MUX2_X1 _11716_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][63] ),
    .S(_05935_),
    .Z(_06208_));
 NOR2_X1 _11717_ (.A1(_05909_),
    .A2(_06208_),
    .ZN(_06209_));
 MUX2_X1 _11718_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][63] ),
    .S(_05935_),
    .Z(_06210_));
 NOR2_X1 _11719_ (.A1(_05946_),
    .A2(_06210_),
    .ZN(_06211_));
 NAND2_X1 _11720_ (.A1(_06031_),
    .A2(_05718_),
    .ZN(_06212_));
 MUX2_X1 _11721_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][63] ),
    .S(_05967_),
    .Z(_06213_));
 NOR2_X1 _11722_ (.A1(_05909_),
    .A2(_06213_),
    .ZN(_06214_));
 MUX2_X1 _11723_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][63] ),
    .S(_05967_),
    .Z(_06215_));
 NOR2_X1 _11724_ (.A1(_05890_),
    .A2(_06215_),
    .ZN(_06216_));
 OAI33_X1 _11725_ (.A1(_06207_),
    .A2(_06209_),
    .A3(_06211_),
    .B1(_06212_),
    .B2(_06214_),
    .B3(_06216_),
    .ZN(_06217_));
 NAND2_X1 _11726_ (.A1(_05922_),
    .A2(_06009_),
    .ZN(_06218_));
 MUX2_X1 _11727_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][63] ),
    .S(_05914_),
    .Z(_06219_));
 NOR2_X1 _11728_ (.A1(_05909_),
    .A2(_06219_),
    .ZN(_06220_));
 MUX2_X1 _11729_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][63] ),
    .S(_05914_),
    .Z(_06221_));
 NOR2_X1 _11730_ (.A1(_05946_),
    .A2(_06221_),
    .ZN(_06222_));
 OR2_X4 _11731_ (.A1(_05707_),
    .A2(_05717_),
    .ZN(_06223_));
 MUX2_X1 _11732_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[4][63] ),
    .S(_05967_),
    .Z(_06224_));
 NOR2_X1 _11733_ (.A1(_05909_),
    .A2(_06224_),
    .ZN(_06225_));
 MUX2_X1 _11734_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][63] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][63] ),
    .S(_05733_),
    .Z(_06226_));
 NOR2_X1 _11735_ (.A1(_05890_),
    .A2(_06226_),
    .ZN(_06227_));
 OAI33_X1 _11736_ (.A1(_06218_),
    .A2(_06220_),
    .A3(_06222_),
    .B1(_06223_),
    .B2(_06225_),
    .B3(_06227_),
    .ZN(_06228_));
 NOR2_X4 _11737_ (.A1(_06217_),
    .A2(_06228_),
    .ZN(_06229_));
 XOR2_X2 _11738_ (.A(_05221_),
    .B(_06229_),
    .Z(_06230_));
 MUX2_X1 _11739_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][51] ),
    .S(_05943_),
    .Z(_06231_));
 NOR2_X1 _11740_ (.A1(_05915_),
    .A2(_06231_),
    .ZN(_06232_));
 MUX2_X1 _11741_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][51] ),
    .S(_05867_),
    .Z(_06233_));
 NOR3_X1 _11742_ (.A1(_05946_),
    .A2(_05735_),
    .A3(_06233_),
    .ZN(_06234_));
 MUX2_X1 _11743_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][51] ),
    .S(_05867_),
    .Z(_06235_));
 NOR3_X1 _11744_ (.A1(_05909_),
    .A2(_05865_),
    .A3(_06235_),
    .ZN(_06236_));
 MUX2_X1 _11745_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][51] ),
    .S(_05861_),
    .Z(_06237_));
 NOR2_X1 _11746_ (.A1(_05905_),
    .A2(_06237_),
    .ZN(_06238_));
 NOR4_X1 _11747_ (.A1(_06232_),
    .A2(_06234_),
    .A3(_06236_),
    .A4(_06238_),
    .ZN(_06239_));
 MUX2_X1 _11748_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][51] ),
    .S(_05943_),
    .Z(_06240_));
 NOR2_X1 _11749_ (.A1(_05915_),
    .A2(_06240_),
    .ZN(_06241_));
 MUX2_X1 _11750_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][51] ),
    .S(_05861_),
    .Z(_06242_));
 NOR3_X1 _11751_ (.A1(_05909_),
    .A2(_05865_),
    .A3(_06242_),
    .ZN(_06243_));
 MUX2_X1 _11752_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][51] ),
    .S(_05867_),
    .Z(_06244_));
 NOR3_X1 _11753_ (.A1(_05946_),
    .A2(_05735_),
    .A3(_06244_),
    .ZN(_06245_));
 MUX2_X1 _11754_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][51] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][51] ),
    .S(_05861_),
    .Z(_06246_));
 NOR2_X1 _11755_ (.A1(_05905_),
    .A2(_06246_),
    .ZN(_06247_));
 NOR4_X1 _11756_ (.A1(_06241_),
    .A2(_06243_),
    .A3(_06245_),
    .A4(_06247_),
    .ZN(_06248_));
 MUX2_X2 _11757_ (.A(_06239_),
    .B(_06248_),
    .S(_05922_),
    .Z(_06249_));
 XNOR2_X1 _11758_ (.A(_05186_),
    .B(_06249_),
    .ZN(_06250_));
 NAND2_X1 _11759_ (.A1(_06230_),
    .A2(_06250_),
    .ZN(_06251_));
 MUX2_X1 _11760_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][60] ),
    .S(_05735_),
    .Z(_06252_));
 MUX2_X1 _11761_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[11][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][60] ),
    .S(_05735_),
    .Z(_06253_));
 OAI22_X2 _11762_ (.A1(_05891_),
    .A2(_06252_),
    .B1(_06253_),
    .B2(_05894_),
    .ZN(_06254_));
 MUX2_X1 _11763_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][60] ),
    .S(_05735_),
    .Z(_06255_));
 MUX2_X1 _11764_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[10][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][60] ),
    .S(_05735_),
    .Z(_06256_));
 OAI22_X2 _11765_ (.A1(_05872_),
    .A2(_06255_),
    .B1(_06256_),
    .B2(_05875_),
    .ZN(_06257_));
 NOR2_X2 _11766_ (.A1(_06254_),
    .A2(_06257_),
    .ZN(_06258_));
 XNOR2_X2 _11767_ (.A(_05191_),
    .B(_06258_),
    .ZN(_06259_));
 MUX2_X1 _11768_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][54] ),
    .S(_05870_),
    .Z(_06260_));
 MUX2_X1 _11769_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][54] ),
    .S(_05870_),
    .Z(_06261_));
 OAI22_X1 _11770_ (.A1(_06207_),
    .A2(_06260_),
    .B1(_06261_),
    .B2(_06223_),
    .ZN(_06262_));
 BUF_X4 _11771_ (.A(net761),
    .Z(_06263_));
 MUX2_X1 _11772_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][54] ),
    .S(_06263_),
    .Z(_06264_));
 NOR3_X1 _11773_ (.A1(_05887_),
    .A2(_05718_),
    .A3(_06264_),
    .ZN(_06265_));
 MUX2_X1 _11774_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][54] ),
    .S(_05699_),
    .Z(_06266_));
 NOR3_X1 _11775_ (.A1(_05921_),
    .A2(_05861_),
    .A3(_06266_),
    .ZN(_06267_));
 OR3_X2 _11776_ (.A1(_06262_),
    .A2(_06265_),
    .A3(_06267_),
    .ZN(_06268_));
 OAI21_X1 _11777_ (.A(_05736_),
    .B1(_06268_),
    .B2(_05252_),
    .ZN(_06269_));
 MUX2_X1 _11778_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][50] ),
    .S(_05870_),
    .Z(_06270_));
 MUX2_X1 _11779_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][50] ),
    .S(_05870_),
    .Z(_06271_));
 MUX2_X1 _11780_ (.A(_06270_),
    .B(_06271_),
    .S(_05707_),
    .Z(_06272_));
 XOR2_X1 _11781_ (.A(_05247_),
    .B(_06272_),
    .Z(_06273_));
 AOI221_X2 _11782_ (.A(_06269_),
    .B1(_06273_),
    .B2(_06009_),
    .C1(_05252_),
    .C2(_06268_),
    .ZN(_06274_));
 MUX2_X1 _11783_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][52] ),
    .S(_05867_),
    .Z(_06275_));
 NOR3_X2 _11784_ (.A1(_06031_),
    .A2(_05890_),
    .A3(_06275_),
    .ZN(_06276_));
 MUX2_X1 _11785_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][52] ),
    .S(_05867_),
    .Z(_06277_));
 NOR2_X1 _11786_ (.A1(_05872_),
    .A2(_06277_),
    .ZN(_06278_));
 MUX2_X1 _11787_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][52] ),
    .S(_05867_),
    .Z(_06279_));
 NOR2_X1 _11788_ (.A1(_05894_),
    .A2(_06279_),
    .ZN(_06280_));
 MUX2_X1 _11789_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][52] ),
    .S(_05897_),
    .Z(_06281_));
 NOR3_X2 _11790_ (.A1(_05874_),
    .A2(_05700_),
    .A3(_06281_),
    .ZN(_06282_));
 NOR4_X4 _11791_ (.A1(_06276_),
    .A2(_06278_),
    .A3(_06280_),
    .A4(_06282_),
    .ZN(_06283_));
 XOR2_X1 _11792_ (.A(_05257_),
    .B(_06283_),
    .Z(_06284_));
 NOR2_X1 _11793_ (.A1(_05737_),
    .A2(_06284_),
    .ZN(_06285_));
 OAI22_X4 _11794_ (.A1(_05720_),
    .A2(_06259_),
    .B1(_06274_),
    .B2(_06285_),
    .ZN(_06286_));
 INV_X1 _11795_ (.A(_05231_),
    .ZN(_06287_));
 MUX2_X1 _11796_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][57] ),
    .S(_06129_),
    .Z(_06288_));
 MUX2_X1 _11797_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][57] ),
    .S(_06129_),
    .Z(_06289_));
 MUX2_X1 _11798_ (.A(_06288_),
    .B(_06289_),
    .S(_05708_),
    .Z(_06290_));
 MUX2_X1 _11799_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][57] ),
    .S(_06129_),
    .Z(_06291_));
 MUX2_X1 _11800_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][57] ),
    .S(_06129_),
    .Z(_06292_));
 MUX2_X1 _11801_ (.A(_06291_),
    .B(_06292_),
    .S(_05708_),
    .Z(_06293_));
 MUX2_X1 _11802_ (.A(_06290_),
    .B(_06293_),
    .S(_05719_),
    .Z(_06294_));
 AOI21_X1 _11803_ (.A(_06287_),
    .B1(_05736_),
    .B2(_06294_),
    .ZN(_06295_));
 MUX2_X1 _11804_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][57] ),
    .S(_05866_),
    .Z(_06296_));
 NOR3_X2 _11805_ (.A1(_05921_),
    .A2(_05908_),
    .A3(_06296_),
    .ZN(_06297_));
 MUX2_X1 _11806_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][57] ),
    .S(_05866_),
    .Z(_06298_));
 NOR2_X1 _11807_ (.A1(_05893_),
    .A2(_06298_),
    .ZN(_06299_));
 MUX2_X1 _11808_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][57] ),
    .S(_05876_),
    .Z(_06300_));
 NOR2_X1 _11809_ (.A1(_05871_),
    .A2(_06300_),
    .ZN(_06301_));
 MUX2_X1 _11810_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][57] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][57] ),
    .S(_05716_),
    .Z(_06302_));
 NOR3_X2 _11811_ (.A1(_05707_),
    .A2(_05889_),
    .A3(_06302_),
    .ZN(_06303_));
 NOR4_X4 _11812_ (.A1(_06297_),
    .A2(_06299_),
    .A3(_06301_),
    .A4(_06303_),
    .ZN(_06304_));
 MUX2_X1 _11813_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][60] ),
    .S(_05699_),
    .Z(_06305_));
 MUX2_X1 _11814_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][60] ),
    .S(_05699_),
    .Z(_06306_));
 MUX2_X1 _11815_ (.A(_06305_),
    .B(_06306_),
    .S(_05707_),
    .Z(_06307_));
 XNOR2_X1 _11816_ (.A(_05191_),
    .B(_06307_),
    .ZN(_06308_));
 OAI21_X1 _11817_ (.A(_06304_),
    .B1(_06308_),
    .B2(_06009_),
    .ZN(_06309_));
 OAI21_X1 _11818_ (.A(_06295_),
    .B1(_06309_),
    .B2(_05737_),
    .ZN(_06310_));
 XOR2_X1 _11819_ (.A(_05191_),
    .B(_06307_),
    .Z(_06311_));
 AOI211_X2 _11820_ (.A(_05735_),
    .B(_06304_),
    .C1(_06311_),
    .C2(_05719_),
    .ZN(_06312_));
 OAI21_X1 _11821_ (.A(_06287_),
    .B1(_05977_),
    .B2(_06294_),
    .ZN(_06313_));
 OR2_X1 _11822_ (.A1(_06312_),
    .A2(_06313_),
    .ZN(_06314_));
 MUX2_X1 _11823_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][53] ),
    .S(_05866_),
    .Z(_06315_));
 MUX2_X1 _11824_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][53] ),
    .S(_05866_),
    .Z(_06316_));
 MUX2_X1 _11825_ (.A(_06315_),
    .B(_06316_),
    .S(_05903_),
    .Z(_06317_));
 MUX2_X1 _11826_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][53] ),
    .S(_05866_),
    .Z(_06318_));
 BUF_X4 _11827_ (.A(_05716_),
    .Z(_06319_));
 MUX2_X1 _11828_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][53] ),
    .S(_06319_),
    .Z(_06320_));
 MUX2_X1 _11829_ (.A(_06318_),
    .B(_06320_),
    .S(_05903_),
    .Z(_06321_));
 MUX2_X1 _11830_ (.A(_06317_),
    .B(_06321_),
    .S(_05865_),
    .Z(_06322_));
 MUX2_X1 _11831_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][53] ),
    .S(_05876_),
    .Z(_06323_));
 MUX2_X1 _11832_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][53] ),
    .S(_05876_),
    .Z(_06324_));
 MUX2_X1 _11833_ (.A(_06323_),
    .B(_06324_),
    .S(_05700_),
    .Z(_06325_));
 MUX2_X1 _11834_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][53] ),
    .S(_05866_),
    .Z(_06326_));
 MUX2_X1 _11835_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][53] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][53] ),
    .S(_05866_),
    .Z(_06327_));
 MUX2_X1 _11836_ (.A(_06326_),
    .B(_06327_),
    .S(_05700_),
    .Z(_06328_));
 MUX2_X1 _11837_ (.A(_06325_),
    .B(_06328_),
    .S(_05865_),
    .Z(_06329_));
 MUX2_X2 _11838_ (.A(_06322_),
    .B(_06329_),
    .S(_05922_),
    .Z(_06330_));
 XNOR2_X1 _11839_ (.A(_05242_),
    .B(_06330_),
    .ZN(_06331_));
 MUX2_X1 _11840_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][56] ),
    .S(_05717_),
    .Z(_06332_));
 MUX2_X1 _11841_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][56] ),
    .S(_05717_),
    .Z(_06333_));
 MUX2_X1 _11842_ (.A(_06332_),
    .B(_06333_),
    .S(_05889_),
    .Z(_06334_));
 NAND2_X2 _11843_ (.A1(_05708_),
    .A2(_05865_),
    .ZN(_06335_));
 NAND2_X1 _11844_ (.A1(_05888_),
    .A2(_05734_),
    .ZN(_06336_));
 MUX2_X1 _11845_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][56] ),
    .S(_06319_),
    .Z(_06337_));
 MUX2_X1 _11846_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][56] ),
    .S(_06319_),
    .Z(_06338_));
 MUX2_X1 _11847_ (.A(_06337_),
    .B(_06338_),
    .S(_05889_),
    .Z(_06339_));
 OAI22_X4 _11848_ (.A1(_06334_),
    .A2(_06335_),
    .B1(_06336_),
    .B2(_06339_),
    .ZN(_06340_));
 MUX2_X1 _11849_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][56] ),
    .S(_05717_),
    .Z(_06341_));
 MUX2_X1 _11850_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][56] ),
    .S(_05717_),
    .Z(_06342_));
 MUX2_X1 _11851_ (.A(_06341_),
    .B(_06342_),
    .S(_05864_),
    .Z(_06343_));
 MUX2_X1 _11852_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][56] ),
    .S(_06319_),
    .Z(_06344_));
 MUX2_X1 _11853_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][56] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][56] ),
    .S(_06319_),
    .Z(_06345_));
 MUX2_X1 _11854_ (.A(_06344_),
    .B(_06345_),
    .S(_05864_),
    .Z(_06346_));
 OAI22_X4 _11855_ (.A1(_05872_),
    .A2(_06343_),
    .B1(_06346_),
    .B2(_05875_),
    .ZN(_06347_));
 OR3_X1 _11856_ (.A1(_05204_),
    .A2(_06340_),
    .A3(_06347_),
    .ZN(_06348_));
 OAI21_X1 _11857_ (.A(_05204_),
    .B1(_06340_),
    .B2(_06347_),
    .ZN(_06349_));
 MUX2_X1 _11858_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][62] ),
    .S(_06263_),
    .Z(_06350_));
 MUX2_X1 _11859_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][62] ),
    .S(_06263_),
    .Z(_06351_));
 MUX2_X1 _11860_ (.A(_06350_),
    .B(_06351_),
    .S(_05921_),
    .Z(_06352_));
 MUX2_X1 _11861_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][62] ),
    .S(_06263_),
    .Z(_06353_));
 MUX2_X1 _11862_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][62] ),
    .S(_06263_),
    .Z(_06354_));
 MUX2_X1 _11863_ (.A(_06353_),
    .B(_06354_),
    .S(_05873_),
    .Z(_06355_));
 NAND2_X1 _11864_ (.A1(_05734_),
    .A2(_05943_),
    .ZN(_06356_));
 OAI22_X4 _11865_ (.A1(_05979_),
    .A2(_06352_),
    .B1(_06355_),
    .B2(_06356_),
    .ZN(_06357_));
 MUX2_X1 _11866_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][62] ),
    .S(_06319_),
    .Z(_06358_));
 MUX2_X1 _11867_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][62] ),
    .S(_06319_),
    .Z(_06359_));
 MUX2_X1 _11868_ (.A(_06358_),
    .B(_06359_),
    .S(_05889_),
    .Z(_06360_));
 NAND2_X1 _11869_ (.A1(_05874_),
    .A2(_05864_),
    .ZN(_06361_));
 MUX2_X1 _11870_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][62] ),
    .S(_05876_),
    .Z(_06362_));
 MUX2_X1 _11871_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][62] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][62] ),
    .S(_05876_),
    .Z(_06363_));
 MUX2_X1 _11872_ (.A(_06362_),
    .B(_06363_),
    .S(_05889_),
    .Z(_06364_));
 OAI22_X4 _11873_ (.A1(_06335_),
    .A2(_06360_),
    .B1(_06361_),
    .B2(_06364_),
    .ZN(_06365_));
 OR3_X1 _11874_ (.A1(_05197_),
    .A2(_06357_),
    .A3(_06365_),
    .ZN(_06366_));
 OAI21_X1 _11875_ (.A(_05197_),
    .B1(_06357_),
    .B2(_06365_),
    .ZN(_06367_));
 AND4_X1 _11876_ (.A1(_06348_),
    .A2(_06349_),
    .A3(_06366_),
    .A4(_06367_),
    .ZN(_06368_));
 NAND4_X2 _11877_ (.A1(_06310_),
    .A2(_06314_),
    .A3(_06331_),
    .A4(_06368_),
    .ZN(_06369_));
 MUX2_X1 _11878_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][61] ),
    .S(_05877_),
    .Z(_06370_));
 NOR3_X1 _11879_ (.A1(_05938_),
    .A2(_05890_),
    .A3(_06370_),
    .ZN(_06371_));
 MUX2_X1 _11880_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][61] ),
    .S(_05897_),
    .Z(_06372_));
 NOR3_X1 _11881_ (.A1(_05874_),
    .A2(_05700_),
    .A3(_06372_),
    .ZN(_06373_));
 MUX2_X1 _11882_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][61] ),
    .S(_05897_),
    .Z(_06374_));
 MUX2_X1 _11883_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][61] ),
    .S(_05897_),
    .Z(_06375_));
 OAI22_X2 _11884_ (.A1(_05872_),
    .A2(_06374_),
    .B1(_06375_),
    .B2(_05894_),
    .ZN(_06376_));
 NOR3_X2 _11885_ (.A1(_06371_),
    .A2(_06373_),
    .A3(_06376_),
    .ZN(_06377_));
 XOR2_X2 _11886_ (.A(_05236_),
    .B(_06377_),
    .Z(_06378_));
 MUX2_X1 _11887_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][59] ),
    .S(_05717_),
    .Z(_06379_));
 NOR2_X1 _11888_ (.A1(_05871_),
    .A2(_06379_),
    .ZN(_06380_));
 MUX2_X1 _11889_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][59] ),
    .S(_05866_),
    .Z(_06381_));
 NOR3_X2 _11890_ (.A1(_05887_),
    .A2(_05889_),
    .A3(_06381_),
    .ZN(_06382_));
 MUX2_X1 _11891_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][59] ),
    .S(_05876_),
    .Z(_06383_));
 NOR3_X2 _11892_ (.A1(_05921_),
    .A2(_05903_),
    .A3(_06383_),
    .ZN(_06384_));
 MUX2_X1 _11893_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][59] ),
    .S(_06319_),
    .Z(_06385_));
 NOR2_X1 _11894_ (.A1(_05893_),
    .A2(_06385_),
    .ZN(_06386_));
 NOR4_X4 _11895_ (.A1(_06380_),
    .A2(_06382_),
    .A3(_06384_),
    .A4(_06386_),
    .ZN(_06387_));
 XOR2_X2 _11896_ (.A(_05226_),
    .B(_06387_),
    .Z(_06388_));
 MUX2_X1 _11897_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][55] ),
    .S(_05892_),
    .Z(_06389_));
 NOR2_X1 _11898_ (.A1(_06223_),
    .A2(_06389_),
    .ZN(_06390_));
 MUX2_X1 _11899_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][55] ),
    .S(_06263_),
    .Z(_06391_));
 NOR3_X1 _11900_ (.A1(_05921_),
    .A2(_05861_),
    .A3(_06391_),
    .ZN(_06392_));
 MUX2_X1 _11901_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][55] ),
    .S(_05699_),
    .Z(_06393_));
 NOR3_X1 _11902_ (.A1(_05887_),
    .A2(_05718_),
    .A3(_06393_),
    .ZN(_06394_));
 MUX2_X1 _11903_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][55] ),
    .S(_06263_),
    .Z(_06395_));
 NOR2_X1 _11904_ (.A1(_06207_),
    .A2(_06395_),
    .ZN(_06396_));
 NOR4_X2 _11905_ (.A1(_06390_),
    .A2(_06392_),
    .A3(_06394_),
    .A4(_06396_),
    .ZN(_06397_));
 XOR2_X2 _11906_ (.A(_05209_),
    .B(_06397_),
    .Z(_06398_));
 NOR4_X2 _11907_ (.A1(_05736_),
    .A2(_06378_),
    .A3(_06388_),
    .A4(_06398_),
    .ZN(_06399_));
 MUX2_X1 _11908_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][61] ),
    .S(_05867_),
    .Z(_06400_));
 NOR3_X1 _11909_ (.A1(_06031_),
    .A2(_05890_),
    .A3(_06400_),
    .ZN(_06401_));
 MUX2_X1 _11910_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][61] ),
    .S(_05877_),
    .Z(_06402_));
 NOR3_X1 _11911_ (.A1(_05874_),
    .A2(_05700_),
    .A3(_06402_),
    .ZN(_06403_));
 MUX2_X1 _11912_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][61] ),
    .S(_05877_),
    .Z(_06404_));
 MUX2_X1 _11913_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][61] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][61] ),
    .S(_05897_),
    .Z(_06405_));
 OAI22_X1 _11914_ (.A1(_05872_),
    .A2(_06404_),
    .B1(_06405_),
    .B2(_05894_),
    .ZN(_06406_));
 NOR3_X1 _11915_ (.A1(_06401_),
    .A2(_06403_),
    .A3(_06406_),
    .ZN(_06407_));
 XOR2_X1 _11916_ (.A(_05236_),
    .B(_06407_),
    .Z(_06408_));
 MUX2_X1 _11917_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][59] ),
    .S(_05700_),
    .Z(_06409_));
 NOR2_X1 _11918_ (.A1(_06207_),
    .A2(_06409_),
    .ZN(_06410_));
 MUX2_X1 _11919_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][59] ),
    .S(_05870_),
    .Z(_06411_));
 NOR3_X1 _11920_ (.A1(_05708_),
    .A2(_05718_),
    .A3(_06411_),
    .ZN(_06412_));
 MUX2_X1 _11921_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][59] ),
    .S(_05870_),
    .Z(_06413_));
 NOR3_X1 _11922_ (.A1(_05921_),
    .A2(_05943_),
    .A3(_06413_),
    .ZN(_06414_));
 MUX2_X1 _11923_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][59] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][59] ),
    .S(_05892_),
    .Z(_06415_));
 NOR2_X1 _11924_ (.A1(_06223_),
    .A2(_06415_),
    .ZN(_06416_));
 NOR4_X2 _11925_ (.A1(_06410_),
    .A2(_06412_),
    .A3(_06414_),
    .A4(_06416_),
    .ZN(_06417_));
 XOR2_X1 _11926_ (.A(_05226_),
    .B(_06417_),
    .Z(_06418_));
 NOR3_X1 _11927_ (.A1(_05977_),
    .A2(_06408_),
    .A3(_06418_),
    .ZN(_06419_));
 MUX2_X1 _11928_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][52] ),
    .S(_05892_),
    .Z(_06420_));
 NOR3_X1 _11929_ (.A1(_05874_),
    .A2(_05943_),
    .A3(_06420_),
    .ZN(_06421_));
 MUX2_X1 _11930_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][52] ),
    .S(_05892_),
    .Z(_06422_));
 NOR2_X1 _11931_ (.A1(_06223_),
    .A2(_06422_),
    .ZN(_06423_));
 MUX2_X1 _11932_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][52] ),
    .S(_05892_),
    .Z(_06424_));
 NOR2_X1 _11933_ (.A1(_06207_),
    .A2(_06424_),
    .ZN(_06425_));
 MUX2_X1 _11934_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][52] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][52] ),
    .S(_06263_),
    .Z(_06426_));
 NOR3_X1 _11935_ (.A1(_05887_),
    .A2(_05718_),
    .A3(_06426_),
    .ZN(_06427_));
 NOR4_X2 _11936_ (.A1(_06421_),
    .A2(_06423_),
    .A3(_06425_),
    .A4(_06427_),
    .ZN(_06428_));
 XOR2_X1 _11937_ (.A(_05257_),
    .B(_06428_),
    .Z(_06429_));
 MUX2_X1 _11938_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][58] ),
    .S(_05876_),
    .Z(_06430_));
 MUX2_X1 _11939_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[7][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][58] ),
    .S(_05876_),
    .Z(_06431_));
 MUX2_X1 _11940_ (.A(_06430_),
    .B(_06431_),
    .S(_05700_),
    .Z(_06432_));
 MUX2_X1 _11941_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[12][58] ),
    .S(_05876_),
    .Z(_06433_));
 MUX2_X1 _11942_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[6][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][58] ),
    .S(_05866_),
    .Z(_06434_));
 MUX2_X1 _11943_ (.A(_06433_),
    .B(_06434_),
    .S(_05700_),
    .Z(_06435_));
 MUX2_X1 _11944_ (.A(_06432_),
    .B(_06435_),
    .S(_05874_),
    .Z(_06436_));
 OR3_X1 _11945_ (.A1(_05215_),
    .A2(_05977_),
    .A3(_06436_),
    .ZN(_06437_));
 NAND3_X1 _11946_ (.A1(_05215_),
    .A2(_05736_),
    .A3(_06436_),
    .ZN(_06438_));
 AOI21_X1 _11947_ (.A(_06429_),
    .B1(_06437_),
    .B2(_06438_),
    .ZN(_06439_));
 MUX2_X1 _11948_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][50] ),
    .S(_05897_),
    .Z(_06440_));
 NOR2_X1 _11949_ (.A1(_05894_),
    .A2(_06440_),
    .ZN(_06441_));
 MUX2_X1 _11950_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][50] ),
    .S(_06319_),
    .Z(_06442_));
 NOR3_X1 _11951_ (.A1(_05921_),
    .A2(_05908_),
    .A3(_06442_),
    .ZN(_06443_));
 MUX2_X1 _11952_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][50] ),
    .S(_06319_),
    .Z(_06444_));
 NOR3_X1 _11953_ (.A1(_05887_),
    .A2(_05889_),
    .A3(_06444_),
    .ZN(_06445_));
 MUX2_X1 _11954_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][50] ),
    .S(_05717_),
    .Z(_06446_));
 NOR2_X1 _11955_ (.A1(_05871_),
    .A2(_06446_),
    .ZN(_06447_));
 NOR4_X2 _11956_ (.A1(_06441_),
    .A2(_06443_),
    .A3(_06445_),
    .A4(_06447_),
    .ZN(_06448_));
 XOR2_X1 _11957_ (.A(_05247_),
    .B(_06448_),
    .Z(_06449_));
 MUX2_X1 _11958_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][58] ),
    .S(_05716_),
    .Z(_06450_));
 MUX2_X1 _11959_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[3][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][58] ),
    .S(_05716_),
    .Z(_06451_));
 MUX2_X1 _11960_ (.A(_06450_),
    .B(_06451_),
    .S(_05700_),
    .Z(_06452_));
 MUX2_X1 _11961_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[8][58] ),
    .S(_05716_),
    .Z(_06453_));
 MUX2_X1 _11962_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[2][58] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][58] ),
    .S(_05716_),
    .Z(_06454_));
 MUX2_X1 _11963_ (.A(_06453_),
    .B(_06454_),
    .S(_05700_),
    .Z(_06455_));
 MUX2_X2 _11964_ (.A(_06452_),
    .B(_06455_),
    .S(_05874_),
    .Z(_06456_));
 OR3_X1 _11965_ (.A1(_05215_),
    .A2(_05736_),
    .A3(_06456_),
    .ZN(_06457_));
 NAND3_X1 _11966_ (.A1(_05215_),
    .A2(_05977_),
    .A3(_06456_),
    .ZN(_06458_));
 AOI21_X1 _11967_ (.A(_06449_),
    .B1(_06457_),
    .B2(_06458_),
    .ZN(_06459_));
 MUX2_X1 _11968_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][50] ),
    .S(_06129_),
    .Z(_06460_));
 MUX2_X1 _11969_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][50] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][50] ),
    .S(_06129_),
    .Z(_06461_));
 MUX2_X1 _11970_ (.A(_06460_),
    .B(_06461_),
    .S(_05708_),
    .Z(_06462_));
 XNOR2_X1 _11971_ (.A(_05247_),
    .B(_06462_),
    .ZN(_06463_));
 MUX2_X1 _11972_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][60] ),
    .S(_06129_),
    .Z(_06464_));
 MUX2_X1 _11973_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][60] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][60] ),
    .S(_06129_),
    .Z(_06465_));
 MUX2_X1 _11974_ (.A(_06464_),
    .B(_06465_),
    .S(_05708_),
    .Z(_06466_));
 XNOR2_X1 _11975_ (.A(_05191_),
    .B(_06466_),
    .ZN(_06467_));
 AOI21_X1 _11976_ (.A(_06009_),
    .B1(_06463_),
    .B2(_06467_),
    .ZN(_06468_));
 MUX2_X1 _11977_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][55] ),
    .S(_05892_),
    .Z(_06469_));
 NOR2_X1 _11978_ (.A1(_06223_),
    .A2(_06469_),
    .ZN(_06470_));
 MUX2_X1 _11979_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][55] ),
    .S(_05699_),
    .Z(_06471_));
 NOR3_X2 _11980_ (.A1(_05921_),
    .A2(_05861_),
    .A3(_06471_),
    .ZN(_06472_));
 MUX2_X1 _11981_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][55] ),
    .S(_05699_),
    .Z(_06473_));
 NOR3_X2 _11982_ (.A1(_05707_),
    .A2(_05718_),
    .A3(_06473_),
    .ZN(_06474_));
 MUX2_X1 _11983_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][55] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][55] ),
    .S(_06263_),
    .Z(_06475_));
 NOR2_X1 _11984_ (.A1(_06207_),
    .A2(_06475_),
    .ZN(_06476_));
 NOR4_X4 _11985_ (.A1(_06470_),
    .A2(_06472_),
    .A3(_06474_),
    .A4(_06476_),
    .ZN(_06477_));
 XOR2_X1 _11986_ (.A(_05209_),
    .B(_06477_),
    .Z(_06478_));
 NOR3_X1 _11987_ (.A1(_05977_),
    .A2(_06468_),
    .A3(_06478_),
    .ZN(_06479_));
 MUX2_X1 _11988_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][54] ),
    .S(_06129_),
    .Z(_06480_));
 NOR2_X1 _11989_ (.A1(_06223_),
    .A2(_06480_),
    .ZN(_06481_));
 MUX2_X1 _11990_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][54] ),
    .S(_06263_),
    .Z(_06482_));
 NOR3_X2 _11991_ (.A1(_05921_),
    .A2(_05861_),
    .A3(_06482_),
    .ZN(_06483_));
 MUX2_X1 _11992_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][54] ),
    .S(_05699_),
    .Z(_06484_));
 NOR3_X2 _11993_ (.A1(_05887_),
    .A2(_05718_),
    .A3(_06484_),
    .ZN(_06485_));
 MUX2_X1 _11994_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][54] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][54] ),
    .S(_05870_),
    .Z(_06486_));
 NOR2_X1 _11995_ (.A1(_06207_),
    .A2(_06486_),
    .ZN(_06487_));
 NOR4_X4 _11996_ (.A1(_06481_),
    .A2(_06483_),
    .A3(_06485_),
    .A4(_06487_),
    .ZN(_06488_));
 XOR2_X1 _11997_ (.A(_05252_),
    .B(_06488_),
    .Z(_06489_));
 NOR2_X1 _11998_ (.A1(_05736_),
    .A2(_06489_),
    .ZN(_06490_));
 OAI222_X2 _11999_ (.A1(_06399_),
    .A2(_06419_),
    .B1(_06439_),
    .B2(_06459_),
    .C1(_06479_),
    .C2(_06490_),
    .ZN(_06491_));
 NOR4_X4 _12000_ (.A1(_06251_),
    .A2(_06286_),
    .A3(_06369_),
    .A4(_06491_),
    .ZN(_06492_));
 MUX2_X2 _12001_ (.A(_06185_),
    .B(_06206_),
    .S(_06492_),
    .Z(_06493_));
 NOR2_X2 _12002_ (.A1(_05263_),
    .A2(_05382_),
    .ZN(_06494_));
 NAND4_X2 _12003_ (.A1(_10260_),
    .A2(_10263_),
    .A3(_05267_),
    .A4(_05268_),
    .ZN(_06495_));
 NOR3_X1 _12004_ (.A1(_10259_),
    .A2(_10271_),
    .A3(_10274_),
    .ZN(_06496_));
 INV_X1 _12005_ (.A(_10256_),
    .ZN(_06497_));
 INV_X1 _12006_ (.A(_10257_),
    .ZN(_06498_));
 OAI21_X1 _12007_ (.A(_06497_),
    .B1(_10253_),
    .B2(_06498_),
    .ZN(_06499_));
 AOI21_X1 _12008_ (.A(_10262_),
    .B1(_06499_),
    .B2(_10263_),
    .ZN(_06500_));
 INV_X1 _12009_ (.A(_10260_),
    .ZN(_06501_));
 OAI21_X1 _12010_ (.A(_06496_),
    .B1(_06500_),
    .B2(_06501_),
    .ZN(_06502_));
 NOR2_X1 _12011_ (.A1(_10272_),
    .A2(_10271_),
    .ZN(_06503_));
 NOR3_X1 _12012_ (.A1(_10275_),
    .A2(_10271_),
    .A3(_10274_),
    .ZN(_06504_));
 NOR2_X1 _12013_ (.A1(_06503_),
    .A2(_06504_),
    .ZN(_06505_));
 NAND3_X2 _12014_ (.A1(_05268_),
    .A2(_06502_),
    .A3(_06505_),
    .ZN(_06506_));
 AOI21_X2 _12015_ (.A(_10265_),
    .B1(_10268_),
    .B2(_10266_),
    .ZN(_06507_));
 NAND3_X2 _12016_ (.A1(_06495_),
    .A2(_06506_),
    .A3(_06507_),
    .ZN(_06508_));
 AND2_X1 _12017_ (.A1(_05266_),
    .A2(_05263_),
    .ZN(_06509_));
 AOI21_X4 _12018_ (.A(_06494_),
    .B1(_06508_),
    .B2(_06509_),
    .ZN(_06510_));
 AND2_X1 _12019_ (.A1(\dynamic_node_top.west_input.control.header_last_temp ),
    .A2(_05175_),
    .ZN(_06511_));
 OR2_X1 _12020_ (.A1(_05152_),
    .A2(_05275_),
    .ZN(_06512_));
 OAI21_X4 _12021_ (.A(_06512_),
    .B1(_05276_),
    .B2(_05201_),
    .ZN(_06513_));
 MUX2_X2 _12022_ (.A(_05278_),
    .B(_05280_),
    .S(_05152_),
    .Z(_06514_));
 NOR3_X2 _12023_ (.A1(_05274_),
    .A2(_06513_),
    .A3(_06514_),
    .ZN(_06515_));
 OR4_X2 _12024_ (.A1(_05196_),
    .A2(_05220_),
    .A3(_05241_),
    .A4(_05262_),
    .ZN(_06516_));
 MUX2_X1 _12025_ (.A(_06495_),
    .B(_05383_),
    .S(_06516_),
    .Z(_06517_));
 OAI21_X2 _12026_ (.A(_06511_),
    .B1(_06515_),
    .B2(_06517_),
    .ZN(_06518_));
 OAI21_X1 _12027_ (.A(_06090_),
    .B1(_06510_),
    .B2(_06518_),
    .ZN(_06519_));
 INV_X1 _12028_ (.A(_05821_),
    .ZN(_06520_));
 AOI21_X1 _12029_ (.A(_06493_),
    .B1(_06519_),
    .B2(_06520_),
    .ZN(_06521_));
 NOR2_X1 _12030_ (.A1(_05823_),
    .A2(_06521_),
    .ZN(_06522_));
 NOR4_X4 _12031_ (.A1(_05406_),
    .A2(_05424_),
    .A3(_05441_),
    .A4(_05450_),
    .ZN(_06523_));
 MUX2_X2 _12032_ (.A(_05363_),
    .B(_05365_),
    .S(_05320_),
    .Z(_06524_));
 OAI211_X2 _12033_ (.A(_06524_),
    .B(_05370_),
    .C1(_05372_),
    .C2(_05374_),
    .ZN(_06525_));
 NAND2_X1 _12034_ (.A1(_05303_),
    .A2(_06525_),
    .ZN(_06526_));
 NAND3_X1 _12035_ (.A1(_05300_),
    .A2(_05386_),
    .A3(_06526_),
    .ZN(_06527_));
 OR2_X1 _12036_ (.A1(_06523_),
    .A2(_06527_),
    .ZN(_06528_));
 NAND4_X1 _12037_ (.A1(_05351_),
    .A2(_05377_),
    .A3(_05378_),
    .A4(_06525_),
    .ZN(_06529_));
 AOI21_X1 _12038_ (.A(_10301_),
    .B1(_05360_),
    .B2(net631),
    .ZN(_06530_));
 NAND4_X1 _12039_ (.A1(net649),
    .A2(_10305_),
    .A3(net634),
    .A4(_10311_),
    .ZN(_06531_));
 INV_X1 _12040_ (.A(_10319_),
    .ZN(_06532_));
 INV_X1 _12041_ (.A(_10320_),
    .ZN(_06533_));
 OAI21_X1 _12042_ (.A(_06532_),
    .B1(_10322_),
    .B2(_06533_),
    .ZN(_06534_));
 AOI221_X2 _12043_ (.A(_10313_),
    .B1(_06534_),
    .B2(_05377_),
    .C1(_10316_),
    .C2(net681),
    .ZN(_06535_));
 OAI211_X2 _12044_ (.A(_06530_),
    .B(_05379_),
    .C1(_06531_),
    .C2(_06535_),
    .ZN(_06536_));
 NAND3_X1 _12045_ (.A1(_05350_),
    .A2(_06529_),
    .A3(_06536_),
    .ZN(_06537_));
 OAI21_X2 _12046_ (.A(_06528_),
    .B1(_06537_),
    .B2(_05451_),
    .ZN(_06538_));
 CLKBUF_X3 _12047_ (.A(\dynamic_node_top.REG_reset_fin.q ),
    .Z(_06539_));
 BUF_X8 _12048_ (.A(_06539_),
    .Z(_06540_));
 BUF_X4 _12049_ (.A(_06540_),
    .Z(_06541_));
 AOI21_X1 _12050_ (.A(_06541_),
    .B1(_06123_),
    .B2(_06125_),
    .ZN(_06542_));
 NOR2_X1 _12051_ (.A1(_05382_),
    .A2(_05489_),
    .ZN(_06543_));
 OR2_X1 _12052_ (.A1(_05463_),
    .A2(_05490_),
    .ZN(_06544_));
 OAI21_X4 _12053_ (.A(_06544_),
    .B1(_05491_),
    .B2(_05495_),
    .ZN(_06545_));
 NOR2_X2 _12054_ (.A1(_05494_),
    .A2(_05497_),
    .ZN(_06546_));
 OR2_X1 _12055_ (.A1(_05463_),
    .A2(_05498_),
    .ZN(_06547_));
 OAI21_X4 _12056_ (.A(_06547_),
    .B1(_05499_),
    .B2(_05495_),
    .ZN(_06548_));
 NOR3_X2 _12057_ (.A1(_06545_),
    .A2(_06546_),
    .A3(_06548_),
    .ZN(_06549_));
 OAI21_X1 _12058_ (.A(_06543_),
    .B1(_06549_),
    .B2(_05383_),
    .ZN(_06550_));
 OR2_X1 _12059_ (.A1(_10365_),
    .A2(_10364_),
    .ZN(_06551_));
 AOI21_X1 _12060_ (.A(_10361_),
    .B1(_06551_),
    .B2(net654),
    .ZN(_06552_));
 NOR3_X1 _12061_ (.A1(_05489_),
    .A2(_05509_),
    .A3(_06552_),
    .ZN(_06553_));
 OR3_X1 _12062_ (.A1(_10361_),
    .A2(_10364_),
    .A3(_05513_),
    .ZN(_06554_));
 OR3_X1 _12063_ (.A1(_10355_),
    .A2(_10367_),
    .A3(_10370_),
    .ZN(_06555_));
 AOI21_X1 _12064_ (.A(_06555_),
    .B1(_10358_),
    .B2(net719),
    .ZN(_06556_));
 INV_X1 _12065_ (.A(_10349_),
    .ZN(_06557_));
 AOI21_X1 _12066_ (.A(_10352_),
    .B1(_06557_),
    .B2(net718),
    .ZN(_06558_));
 NAND2_X1 _12067_ (.A1(net719),
    .A2(net725),
    .ZN(_06559_));
 OAI21_X1 _12068_ (.A(_06556_),
    .B1(_06558_),
    .B2(_06559_),
    .ZN(_06560_));
 INV_X1 _12069_ (.A(_10367_),
    .ZN(_06561_));
 OAI21_X1 _12070_ (.A(_10368_),
    .B1(_10370_),
    .B2(_10371_),
    .ZN(_06562_));
 NAND2_X1 _12071_ (.A1(_06561_),
    .A2(_06562_),
    .ZN(_06563_));
 AND2_X1 _12072_ (.A1(_06560_),
    .A2(_06563_),
    .ZN(_06564_));
 OR3_X2 _12073_ (.A1(_05510_),
    .A2(_05511_),
    .A3(_05512_),
    .ZN(_06565_));
 OAI221_X2 _12074_ (.A(_06553_),
    .B1(_06554_),
    .B2(_06564_),
    .C1(_06565_),
    .C2(_06549_),
    .ZN(_06566_));
 CLKBUF_X3 _12075_ (.A(_05589_),
    .Z(_06567_));
 MUX2_X2 _12076_ (.A(_06550_),
    .B(_06566_),
    .S(_06567_),
    .Z(_06568_));
 NAND3_X1 _12077_ (.A1(_06538_),
    .A2(_06542_),
    .A3(_06568_),
    .ZN(_06569_));
 NAND2_X1 _12078_ (.A1(_06538_),
    .A2(_06542_),
    .ZN(_06570_));
 INV_X1 _12079_ (.A(_05757_),
    .ZN(_06571_));
 OAI221_X1 _12080_ (.A(_06128_),
    .B1(_06522_),
    .B2(_06569_),
    .C1(_06570_),
    .C2(_06571_),
    .ZN(_00018_));
 CLKBUF_X3 _12081_ (.A(_06541_),
    .Z(_06572_));
 BUF_X4 _12082_ (.A(_06572_),
    .Z(_06573_));
 NOR2_X1 _12083_ (.A1(_06510_),
    .A2(_06518_),
    .ZN(_06574_));
 BUF_X4 _12084_ (.A(_05753_),
    .Z(_06575_));
 NOR2_X1 _12085_ (.A1(_06571_),
    .A2(_06540_),
    .ZN(_06576_));
 MUX2_X1 _12086_ (.A(_06537_),
    .B(_06527_),
    .S(_05451_),
    .Z(_06577_));
 AND2_X1 _12087_ (.A1(_06120_),
    .A2(_06577_),
    .ZN(_06578_));
 AOI22_X1 _12088_ (.A1(_06575_),
    .A2(_06568_),
    .B1(_06576_),
    .B2(_06578_),
    .ZN(_06579_));
 NOR2_X1 _12089_ (.A1(_05753_),
    .A2(_06577_),
    .ZN(_06580_));
 INV_X4 _12090_ (.A(_06539_),
    .ZN(_06581_));
 AOI221_X2 _12091_ (.A(_05753_),
    .B1(_05757_),
    .B2(_06581_),
    .C1(_06568_),
    .C2(_05823_),
    .ZN(_06582_));
 OAI33_X1 _12092_ (.A1(_06493_),
    .A2(_06574_),
    .A3(_06579_),
    .B1(_06580_),
    .B2(_06582_),
    .B3(_06120_),
    .ZN(_06583_));
 NOR3_X1 _12093_ (.A1(_06573_),
    .A2(_06127_),
    .A3(_06583_),
    .ZN(_06584_));
 AND2_X1 _12094_ (.A1(_06577_),
    .A2(_06568_),
    .ZN(_06585_));
 NAND2_X1 _12095_ (.A1(_05823_),
    .A2(net667),
    .ZN(_06586_));
 NOR2_X1 _12096_ (.A1(_06574_),
    .A2(_06586_),
    .ZN(_06587_));
 OAI21_X1 _12097_ (.A(_06585_),
    .B1(_06587_),
    .B2(_06521_),
    .ZN(_06588_));
 BUF_X4 _12098_ (.A(_06541_),
    .Z(_06589_));
 AOI21_X1 _12099_ (.A(_06589_),
    .B1(_05756_),
    .B2(_06090_),
    .ZN(_06590_));
 AOI22_X1 _12100_ (.A1(_06584_),
    .A2(_06588_),
    .B1(_06590_),
    .B2(_06127_),
    .ZN(_00017_));
 BUF_X4 _12101_ (.A(_05756_),
    .Z(_06591_));
 NAND2_X1 _12102_ (.A1(_05858_),
    .A2(\dynamic_node_top.proc_input.control.count_one_f ),
    .ZN(_06592_));
 OR4_X1 _12103_ (.A1(_05902_),
    .A2(_05933_),
    .A3(_05956_),
    .A4(_05972_),
    .ZN(_06593_));
 AND2_X2 _12104_ (.A1(_06000_),
    .A2(_06007_),
    .ZN(_06594_));
 NOR3_X1 _12105_ (.A1(_06009_),
    .A2(_06018_),
    .A3(_06027_),
    .ZN(_06595_));
 AND3_X1 _12106_ (.A1(_06009_),
    .A2(_06038_),
    .A3(_06047_),
    .ZN(_06596_));
 OAI221_X2 _12107_ (.A(_06594_),
    .B1(_06595_),
    .B2(_06596_),
    .C1(_05983_),
    .C2(_05992_),
    .ZN(_06597_));
 OAI221_X2 _12108_ (.A(_06592_),
    .B1(_06593_),
    .B2(_06597_),
    .C1(_05858_),
    .C2(_05859_),
    .ZN(_06598_));
 NOR2_X1 _12109_ (.A1(_05786_),
    .A2(_05788_),
    .ZN(_06599_));
 NAND2_X1 _12110_ (.A1(_05472_),
    .A2(_06599_),
    .ZN(_06600_));
 NOR2_X4 _12111_ (.A1(_05826_),
    .A2(_05854_),
    .ZN(_06601_));
 INV_X1 _12112_ (.A(_05478_),
    .ZN(_06602_));
 INV_X1 _12113_ (.A(_05470_),
    .ZN(_06603_));
 OAI221_X2 _12114_ (.A(_05473_),
    .B1(_06601_),
    .B2(_06602_),
    .C1(_06083_),
    .C2(_06603_),
    .ZN(_06604_));
 AOI222_X2 _12115_ (.A1(_05484_),
    .A2(_06598_),
    .B1(_06600_),
    .B2(_06604_),
    .C1(_05820_),
    .C2(_05471_),
    .ZN(_06605_));
 MUX2_X1 _12116_ (.A(\dynamic_node_top.west_output.control.planned_f ),
    .B(_06605_),
    .S(net625),
    .Z(_06606_));
 BUF_X2 _12117_ (.A(_06606_),
    .Z(_06607_));
 NAND3_X1 _12118_ (.A1(_05470_),
    .A2(_06591_),
    .A3(_06607_),
    .ZN(_06608_));
 BUF_X4 _12119_ (.A(_05471_),
    .Z(_06609_));
 INV_X4 _12120_ (.A(_06609_),
    .ZN(_06610_));
 BUF_X4 _12121_ (.A(_06610_),
    .Z(_06611_));
 BUF_X4 _12122_ (.A(_06611_),
    .Z(_06612_));
 BUF_X4 _12123_ (.A(_05185_),
    .Z(_06613_));
 OR2_X1 _12124_ (.A1(net770),
    .A2(_05266_),
    .ZN(_06614_));
 MUX2_X2 _12125_ (.A(_05300_),
    .B(_06614_),
    .S(_05263_),
    .Z(_06615_));
 MUX2_X1 _12126_ (.A(_05270_),
    .B(_05304_),
    .S(_06516_),
    .Z(_06616_));
 OR4_X2 _12127_ (.A1(_05273_),
    .A2(_05277_),
    .A3(_05281_),
    .A4(_06616_),
    .ZN(_06617_));
 AOI21_X4 _12128_ (.A(_06613_),
    .B1(_06615_),
    .B2(_06617_),
    .ZN(_06618_));
 OR2_X1 _12129_ (.A1(_06524_),
    .A2(_05370_),
    .ZN(_06619_));
 NOR3_X1 _12130_ (.A1(_05383_),
    .A2(_05376_),
    .A3(_06619_),
    .ZN(_06620_));
 OR3_X1 _12131_ (.A1(_05382_),
    .A2(_06523_),
    .A3(_06620_),
    .ZN(_06621_));
 NOR3_X1 _12132_ (.A1(_05376_),
    .A2(_05379_),
    .A3(_06619_),
    .ZN(_06622_));
 AOI21_X1 _12133_ (.A(_10298_),
    .B1(_10299_),
    .B2(_10295_),
    .ZN(_06623_));
 OAI21_X1 _12134_ (.A(_10293_),
    .B1(_10290_),
    .B2(_10289_),
    .ZN(_06624_));
 INV_X1 _12135_ (.A(_06624_),
    .ZN(_06625_));
 OAI21_X1 _12136_ (.A(_05348_),
    .B1(_06625_),
    .B2(_10292_),
    .ZN(_06626_));
 OR3_X1 _12137_ (.A1(_10289_),
    .A2(_10286_),
    .A3(_10292_),
    .ZN(_06627_));
 INV_X1 _12138_ (.A(_10283_),
    .ZN(_06628_));
 INV_X1 _12139_ (.A(net695),
    .ZN(_06629_));
 INV_X1 _12140_ (.A(_10277_),
    .ZN(_06630_));
 AOI21_X1 _12141_ (.A(_10280_),
    .B1(_06630_),
    .B2(_10281_),
    .ZN(_06631_));
 OAI21_X1 _12142_ (.A(_06628_),
    .B1(_06629_),
    .B2(_06631_),
    .ZN(_06632_));
 AOI21_X1 _12143_ (.A(_06627_),
    .B1(_06632_),
    .B2(_10287_),
    .ZN(_06633_));
 OAI21_X2 _12144_ (.A(_06623_),
    .B1(_06626_),
    .B2(_06633_),
    .ZN(_06634_));
 MUX2_X1 _12145_ (.A(_06622_),
    .B(_06634_),
    .S(_05349_),
    .Z(_06635_));
 OAI211_X4 _12146_ (.A(_05386_),
    .B(_06621_),
    .C1(_06635_),
    .C2(_05451_),
    .ZN(_06636_));
 AOI21_X1 _12147_ (.A(_05478_),
    .B1(_05484_),
    .B2(_06636_),
    .ZN(_06637_));
 OAI21_X1 _12148_ (.A(_06612_),
    .B1(_06618_),
    .B2(_06637_),
    .ZN(_06638_));
 AOI21_X1 _12149_ (.A(_05481_),
    .B1(net702),
    .B2(_06638_),
    .ZN(_06639_));
 NOR2_X1 _12150_ (.A1(_10192_),
    .A2(_05630_),
    .ZN(_06640_));
 INV_X1 _12151_ (.A(_10195_),
    .ZN(_06641_));
 OAI21_X1 _12152_ (.A(net676),
    .B1(_10198_),
    .B2(_10199_),
    .ZN(_06642_));
 NAND2_X1 _12153_ (.A1(_06641_),
    .A2(_06642_),
    .ZN(_06643_));
 NAND2_X1 _12154_ (.A1(_10193_),
    .A2(_06643_),
    .ZN(_06644_));
 OR3_X1 _12155_ (.A1(_10195_),
    .A2(_10198_),
    .A3(_10201_),
    .ZN(_06645_));
 INV_X1 _12156_ (.A(_10189_),
    .ZN(_06646_));
 INV_X1 _12157_ (.A(_10180_),
    .ZN(_06647_));
 AOI21_X1 _12158_ (.A(_10183_),
    .B1(_06647_),
    .B2(net653),
    .ZN(_06648_));
 INV_X1 _12159_ (.A(net641),
    .ZN(_06649_));
 OAI21_X1 _12160_ (.A(_06646_),
    .B1(_06648_),
    .B2(_06649_),
    .ZN(_06650_));
 AOI221_X2 _12161_ (.A(_06645_),
    .B1(_06650_),
    .B2(_05629_),
    .C1(net659),
    .C2(_10186_),
    .ZN(_06651_));
 OAI21_X1 _12162_ (.A(_06640_),
    .B1(_06644_),
    .B2(_06651_),
    .ZN(_06652_));
 NAND3_X1 _12163_ (.A1(_05617_),
    .A2(_06100_),
    .A3(_05627_),
    .ZN(_06653_));
 NAND2_X1 _12164_ (.A1(_05630_),
    .A2(_06653_),
    .ZN(_06654_));
 AND4_X1 _12165_ (.A1(_06103_),
    .A2(net747),
    .A3(_06652_),
    .A4(_06654_),
    .ZN(_06655_));
 NAND3_X1 _12166_ (.A1(_05303_),
    .A2(_05617_),
    .A3(_06100_),
    .ZN(_06656_));
 AOI21_X2 _12167_ (.A(_06096_),
    .B1(_06656_),
    .B2(_05300_),
    .ZN(_06657_));
 OR4_X4 _12168_ (.A1(_05651_),
    .A2(_05668_),
    .A3(_05685_),
    .A4(_05694_),
    .ZN(_06658_));
 AOI21_X4 _12169_ (.A(_06655_),
    .B1(_06657_),
    .B2(_06658_),
    .ZN(_06659_));
 INV_X1 _12170_ (.A(_06659_),
    .ZN(_06660_));
 NOR2_X2 _12171_ (.A1(_06541_),
    .A2(_06607_),
    .ZN(_06661_));
 NAND2_X1 _12172_ (.A1(_06660_),
    .A2(_06661_),
    .ZN(_06662_));
 OAI21_X1 _12173_ (.A(_06608_),
    .B1(_06639_),
    .B2(_06662_),
    .ZN(_00035_));
 INV_X1 _12174_ (.A(_05755_),
    .ZN(_06663_));
 CLKBUF_X3 _12175_ (.A(_06663_),
    .Z(_06664_));
 NAND2_X1 _12176_ (.A1(_05481_),
    .A2(_06659_),
    .ZN(_06665_));
 CLKBUF_X3 _12177_ (.A(_05919_),
    .Z(_06666_));
 NOR2_X1 _12178_ (.A1(_05737_),
    .A2(_06137_),
    .ZN(_06667_));
 NOR2_X1 _12179_ (.A1(_05977_),
    .A2(_06144_),
    .ZN(_06668_));
 NOR4_X4 _12180_ (.A1(_06667_),
    .A2(_06668_),
    .A3(_06163_),
    .A4(_06178_),
    .ZN(_06669_));
 AOI21_X1 _12181_ (.A(_05382_),
    .B1(_05303_),
    .B2(_06669_),
    .ZN(_06670_));
 OR2_X1 _12182_ (.A1(_06666_),
    .A2(_06670_),
    .ZN(_06671_));
 NOR2_X1 _12183_ (.A1(_06188_),
    .A2(_06191_),
    .ZN(_06672_));
 INV_X1 _12184_ (.A(_10388_),
    .ZN(_06673_));
 AOI21_X1 _12185_ (.A(_10391_),
    .B1(_10394_),
    .B2(_10392_),
    .ZN(_06674_));
 INV_X1 _12186_ (.A(_10389_),
    .ZN(_06675_));
 OAI21_X1 _12187_ (.A(_06673_),
    .B1(_06674_),
    .B2(_06675_),
    .ZN(_06676_));
 AOI21_X1 _12188_ (.A(_10385_),
    .B1(_06676_),
    .B2(_10386_),
    .ZN(_06677_));
 INV_X1 _12189_ (.A(_10382_),
    .ZN(_06678_));
 INV_X1 _12190_ (.A(_10373_),
    .ZN(_06679_));
 AOI21_X1 _12191_ (.A(_10376_),
    .B1(_06679_),
    .B2(_10377_),
    .ZN(_06680_));
 INV_X1 _12192_ (.A(_10383_),
    .ZN(_06681_));
 OAI21_X1 _12193_ (.A(_06678_),
    .B1(_06680_),
    .B2(_06681_),
    .ZN(_06682_));
 AOI21_X1 _12194_ (.A(_10379_),
    .B1(_06682_),
    .B2(_10380_),
    .ZN(_06683_));
 OAI21_X1 _12195_ (.A(_06677_),
    .B1(_06683_),
    .B2(_06186_),
    .ZN(_06684_));
 AOI22_X1 _12196_ (.A1(_06669_),
    .A2(_06672_),
    .B1(_06684_),
    .B2(_06188_),
    .ZN(_06685_));
 OR2_X1 _12197_ (.A1(_06666_),
    .A2(_06685_),
    .ZN(_06686_));
 MUX2_X1 _12198_ (.A(_06671_),
    .B(_06686_),
    .S(_06492_),
    .Z(_06687_));
 NOR3_X1 _12199_ (.A1(_06607_),
    .A2(_06665_),
    .A3(_06687_),
    .ZN(_06688_));
 AOI21_X1 _12200_ (.A(_06688_),
    .B1(_06607_),
    .B2(_05484_),
    .ZN(_06689_));
 AND2_X1 _12201_ (.A1(_05590_),
    .A2(_06659_),
    .ZN(_06690_));
 BUF_X4 _12202_ (.A(_06611_),
    .Z(_06691_));
 OAI21_X1 _12203_ (.A(_06691_),
    .B1(_06618_),
    .B2(_06602_),
    .ZN(_06692_));
 AOI21_X1 _12204_ (.A(_05470_),
    .B1(_06690_),
    .B2(_06692_),
    .ZN(_06693_));
 NOR2_X1 _12205_ (.A1(_06666_),
    .A2(_06670_),
    .ZN(_06694_));
 NOR2_X1 _12206_ (.A1(_06666_),
    .A2(_06685_),
    .ZN(_06695_));
 MUX2_X1 _12207_ (.A(_06694_),
    .B(_06695_),
    .S(_06492_),
    .Z(_06696_));
 BUF_X4 _12208_ (.A(_06696_),
    .Z(_06697_));
 NAND2_X1 _12209_ (.A1(_06661_),
    .A2(_06697_),
    .ZN(_06698_));
 OAI22_X1 _12210_ (.A1(_06664_),
    .A2(_06689_),
    .B1(_06693_),
    .B2(_06698_),
    .ZN(_00034_));
 BUF_X4 _12211_ (.A(_06611_),
    .Z(_06699_));
 INV_X1 _12212_ (.A(_06607_),
    .ZN(_06700_));
 BUF_X4 _12213_ (.A(_06511_),
    .Z(_06701_));
 AOI21_X2 _12214_ (.A(_06494_),
    .B1(_06614_),
    .B2(_05263_),
    .ZN(_06702_));
 NOR3_X1 _12215_ (.A1(_05277_),
    .A2(_05281_),
    .A3(_05304_),
    .ZN(_06703_));
 NOR3_X1 _12216_ (.A1(_05270_),
    .A2(_05277_),
    .A3(_05281_),
    .ZN(_06704_));
 MUX2_X2 _12217_ (.A(_06703_),
    .B(_06704_),
    .S(_05263_),
    .Z(_06705_));
 NOR2_X1 _12218_ (.A1(_06613_),
    .A2(_05273_),
    .ZN(_06706_));
 AOI22_X4 _12219_ (.A1(_06701_),
    .A2(_06702_),
    .B1(_06705_),
    .B2(_06706_),
    .ZN(_06707_));
 NOR2_X1 _12220_ (.A1(_05478_),
    .A2(_06636_),
    .ZN(_06708_));
 NOR2_X1 _12221_ (.A1(_05478_),
    .A2(_05484_),
    .ZN(_06709_));
 AOI21_X1 _12222_ (.A(_05470_),
    .B1(_05481_),
    .B2(_06659_),
    .ZN(_06710_));
 OAI21_X1 _12223_ (.A(_06709_),
    .B1(_06697_),
    .B2(_06710_),
    .ZN(_06711_));
 NAND2_X1 _12224_ (.A1(_06661_),
    .A2(_06711_),
    .ZN(_06712_));
 OAI33_X1 _12225_ (.A1(_06699_),
    .A2(_06664_),
    .A3(_06700_),
    .B1(_06707_),
    .B2(_06708_),
    .B3(_06712_),
    .ZN(_00033_));
 NOR2_X2 _12226_ (.A1(_05817_),
    .A2(_05819_),
    .ZN(_06713_));
 NAND2_X1 _12227_ (.A1(_05160_),
    .A2(_06713_),
    .ZN(_06714_));
 OR2_X2 _12228_ (.A1(_06053_),
    .A2(_06082_),
    .ZN(_06715_));
 AOI22_X2 _12229_ (.A1(_05167_),
    .A2(_05855_),
    .B1(_06715_),
    .B2(_05171_),
    .ZN(_06716_));
 AOI21_X1 _12230_ (.A(_05160_),
    .B1(_05789_),
    .B2(_05159_),
    .ZN(_06717_));
 INV_X1 _12231_ (.A(_05158_),
    .ZN(_06718_));
 OAI211_X2 _12232_ (.A(_06716_),
    .B(_06717_),
    .C1(_06718_),
    .C2(_06050_),
    .ZN(_06719_));
 NAND2_X1 _12233_ (.A1(_06714_),
    .A2(_06719_),
    .ZN(_06720_));
 BUF_X1 _12234_ (.A(\dynamic_node_top.east_output.control.planned_f ),
    .Z(_06721_));
 MUX2_X2 _12235_ (.A(_06720_),
    .B(_06721_),
    .S(_05308_),
    .Z(_06722_));
 NAND3_X1 _12236_ (.A1(_05171_),
    .A2(_06591_),
    .A3(_06722_),
    .ZN(_06723_));
 BUF_X4 _12237_ (.A(_05159_),
    .Z(_06724_));
 OR2_X1 _12238_ (.A1(_05270_),
    .A2(_05282_),
    .ZN(_06725_));
 AOI21_X1 _12239_ (.A(_10229_),
    .B1(_05295_),
    .B2(net636),
    .ZN(_06726_));
 INV_X1 _12240_ (.A(_10244_),
    .ZN(_06727_));
 INV_X1 _12241_ (.A(_10250_),
    .ZN(_06728_));
 AOI21_X1 _12242_ (.A(_10247_),
    .B1(_06728_),
    .B2(_10248_),
    .ZN(_06729_));
 INV_X1 _12243_ (.A(_10245_),
    .ZN(_06730_));
 OAI21_X1 _12244_ (.A(_06727_),
    .B1(_06729_),
    .B2(_06730_),
    .ZN(_06731_));
 AOI21_X1 _12245_ (.A(_10241_),
    .B1(_06731_),
    .B2(_10242_),
    .ZN(_06732_));
 OAI21_X2 _12246_ (.A(_06726_),
    .B1(_06732_),
    .B2(net734),
    .ZN(_06733_));
 AOI21_X2 _12247_ (.A(_06516_),
    .B1(_06725_),
    .B2(_06733_),
    .ZN(_06734_));
 NOR3_X2 _12248_ (.A1(_05282_),
    .A2(_05263_),
    .A3(_05304_),
    .ZN(_06735_));
 OAI21_X4 _12249_ (.A(_06701_),
    .B1(_06734_),
    .B2(_06735_),
    .ZN(_06736_));
 AOI21_X2 _12250_ (.A(_05173_),
    .B1(_06724_),
    .B2(_06736_),
    .ZN(_06737_));
 INV_X1 _12251_ (.A(_06162_),
    .ZN(_06738_));
 NOR3_X2 _12252_ (.A1(_05919_),
    .A2(_06146_),
    .A3(_06179_),
    .ZN(_06739_));
 INV_X1 _12253_ (.A(_06739_),
    .ZN(_06740_));
 NOR3_X1 _12254_ (.A1(_05304_),
    .A2(_06738_),
    .A3(_06740_),
    .ZN(_06741_));
 OR2_X1 _12255_ (.A1(_06666_),
    .A2(_06684_),
    .ZN(_06742_));
 NAND3_X1 _12256_ (.A1(_06163_),
    .A2(_06672_),
    .A3(_06739_),
    .ZN(_06743_));
 NAND2_X1 _12257_ (.A1(_06742_),
    .A2(_06743_),
    .ZN(_06744_));
 MUX2_X2 _12258_ (.A(_06741_),
    .B(_06744_),
    .S(_06492_),
    .Z(_06745_));
 OAI21_X1 _12259_ (.A(_06718_),
    .B1(_06737_),
    .B2(_06745_),
    .ZN(_06746_));
 NAND3_X1 _12260_ (.A1(_05366_),
    .A2(_05370_),
    .A3(_05376_),
    .ZN(_06747_));
 NOR3_X2 _12261_ (.A1(_05304_),
    .A2(_06523_),
    .A3(_06747_),
    .ZN(_06748_));
 OR2_X1 _12262_ (.A1(_05349_),
    .A2(_05379_),
    .ZN(_06749_));
 OR2_X1 _12263_ (.A1(_06747_),
    .A2(_06749_),
    .ZN(_06750_));
 AOI21_X2 _12264_ (.A(_05451_),
    .B1(_06634_),
    .B2(_06750_),
    .ZN(_06751_));
 OAI21_X4 _12265_ (.A(_05386_),
    .B1(_06748_),
    .B2(_06751_),
    .ZN(_06752_));
 AOI21_X1 _12266_ (.A(_05167_),
    .B1(_06746_),
    .B2(_06752_),
    .ZN(_06753_));
 BUF_X4 _12267_ (.A(_06581_),
    .Z(_06754_));
 BUF_X4 _12268_ (.A(_06754_),
    .Z(_06755_));
 AND2_X1 _12269_ (.A1(_06714_),
    .A2(_06719_),
    .ZN(_06756_));
 INV_X1 _12270_ (.A(_06721_),
    .ZN(_06757_));
 MUX2_X1 _12271_ (.A(_06756_),
    .B(_06757_),
    .S(_05308_),
    .Z(_06758_));
 NAND3_X1 _12272_ (.A1(_05613_),
    .A2(_06099_),
    .A3(_05622_),
    .ZN(_06759_));
 OR2_X1 _12273_ (.A1(_05631_),
    .A2(_06759_),
    .ZN(_06760_));
 NOR2_X1 _12274_ (.A1(_10192_),
    .A2(_06096_),
    .ZN(_06761_));
 OAI21_X1 _12275_ (.A(_06761_),
    .B1(_06644_),
    .B2(_06651_),
    .ZN(_06762_));
 AOI21_X2 _12276_ (.A(_06658_),
    .B1(_06760_),
    .B2(_06762_),
    .ZN(_06763_));
 NOR3_X2 _12277_ (.A1(_05304_),
    .A2(net749),
    .A3(_06759_),
    .ZN(_06764_));
 NOR2_X2 _12278_ (.A1(_06763_),
    .A2(_06764_),
    .ZN(_06765_));
 INV_X1 _12279_ (.A(_06765_),
    .ZN(_06766_));
 NAND3_X1 _12280_ (.A1(_06755_),
    .A2(_06758_),
    .A3(_06766_),
    .ZN(_06767_));
 OAI21_X1 _12281_ (.A(_06723_),
    .B1(_06753_),
    .B2(_06767_),
    .ZN(_00041_));
 NOR2_X1 _12282_ (.A1(_06607_),
    .A2(_06618_),
    .ZN(_06768_));
 NAND4_X1 _12283_ (.A1(_05478_),
    .A2(_06754_),
    .A3(_05590_),
    .A4(_06659_),
    .ZN(_06769_));
 NAND2_X1 _12284_ (.A1(_05470_),
    .A2(_06636_),
    .ZN(_06770_));
 AOI21_X1 _12285_ (.A(_06697_),
    .B1(_06769_),
    .B2(_06770_),
    .ZN(_06771_));
 NOR3_X1 _12286_ (.A1(_06602_),
    .A2(_06664_),
    .A3(net702),
    .ZN(_06772_));
 OAI21_X1 _12287_ (.A(_06768_),
    .B1(_06771_),
    .B2(_06772_),
    .ZN(_06773_));
 NAND2_X1 _12288_ (.A1(_05484_),
    .A2(_06636_),
    .ZN(_06774_));
 OAI21_X1 _12289_ (.A(_06612_),
    .B1(_06618_),
    .B2(_06774_),
    .ZN(_06775_));
 INV_X1 _12290_ (.A(_05484_),
    .ZN(_06776_));
 OAI211_X2 _12291_ (.A(net702),
    .B(_06697_),
    .C1(_06618_),
    .C2(_06776_),
    .ZN(_06777_));
 NAND2_X1 _12292_ (.A1(_06636_),
    .A2(_06659_),
    .ZN(_06778_));
 NAND2_X1 _12293_ (.A1(net702),
    .A2(_06778_),
    .ZN(_06779_));
 NAND4_X1 _12294_ (.A1(_06700_),
    .A2(_06775_),
    .A3(_06777_),
    .A4(_06779_),
    .ZN(_06780_));
 NOR3_X1 _12295_ (.A1(_06618_),
    .A2(_06697_),
    .A3(_06778_),
    .ZN(_06781_));
 NAND3_X1 _12296_ (.A1(_05481_),
    .A2(_06700_),
    .A3(_06781_),
    .ZN(_06782_));
 AND2_X1 _12297_ (.A1(_05481_),
    .A2(_05756_),
    .ZN(_06783_));
 AOI21_X1 _12298_ (.A(_06589_),
    .B1(_06607_),
    .B2(_06783_),
    .ZN(_06784_));
 NAND4_X1 _12299_ (.A1(_06773_),
    .A2(_06780_),
    .A3(_06782_),
    .A4(_06784_),
    .ZN(_00032_));
 INV_X1 _12300_ (.A(_05330_),
    .ZN(_06785_));
 CLKBUF_X3 _12301_ (.A(_05384_),
    .Z(_06786_));
 AND2_X2 _12302_ (.A1(_05488_),
    .A2(_05177_),
    .ZN(_06787_));
 OR2_X1 _12303_ (.A1(_05494_),
    .A2(_05497_),
    .ZN(_06788_));
 CLKBUF_X3 _12304_ (.A(_06788_),
    .Z(_06789_));
 NOR3_X2 _12305_ (.A1(_06545_),
    .A2(_06789_),
    .A3(_05500_),
    .ZN(_06790_));
 NAND3_X1 _12306_ (.A1(_06786_),
    .A2(_06787_),
    .A3(_06790_),
    .ZN(_06791_));
 NOR2_X1 _12307_ (.A1(_06567_),
    .A2(_06791_),
    .ZN(_06792_));
 BUF_X4 _12308_ (.A(_05489_),
    .Z(_06793_));
 NAND4_X1 _12309_ (.A1(net656),
    .A2(_10365_),
    .A3(_06560_),
    .A4(_06563_),
    .ZN(_06794_));
 AOI21_X1 _12310_ (.A(_10361_),
    .B1(_10364_),
    .B2(net655),
    .ZN(_06795_));
 AOI22_X2 _12311_ (.A1(_05513_),
    .A2(_06790_),
    .B1(_06794_),
    .B2(_06795_),
    .ZN(_06796_));
 NOR3_X4 _12312_ (.A1(_06793_),
    .A2(net684),
    .A3(_06796_),
    .ZN(_06797_));
 AOI21_X4 _12313_ (.A(_06792_),
    .B1(_06797_),
    .B2(_06567_),
    .ZN(_06798_));
 NAND2_X1 _12314_ (.A1(_05338_),
    .A2(_06798_),
    .ZN(_06799_));
 AND4_X1 _12315_ (.A1(_05266_),
    .A2(_05263_),
    .A3(_06506_),
    .A4(_06507_),
    .ZN(_06800_));
 AOI21_X4 _12316_ (.A(_06800_),
    .B1(_06705_),
    .B2(_05273_),
    .ZN(_06801_));
 NOR2_X2 _12317_ (.A1(_06613_),
    .A2(_06801_),
    .ZN(_06802_));
 OAI21_X1 _12318_ (.A(_06785_),
    .B1(_06799_),
    .B2(_06802_),
    .ZN(_06803_));
 NAND2_X1 _12319_ (.A1(_05331_),
    .A2(_05755_),
    .ZN(_06804_));
 NAND2_X2 _12320_ (.A1(_06581_),
    .A2(_06798_),
    .ZN(_06805_));
 BUF_X4 _12321_ (.A(_05332_),
    .Z(_06806_));
 BUF_X4 _12322_ (.A(_06806_),
    .Z(_06807_));
 NAND2_X1 _12323_ (.A1(_06807_),
    .A2(net680),
    .ZN(_06808_));
 OAI21_X1 _12324_ (.A(_06804_),
    .B1(_06805_),
    .B2(_06808_),
    .ZN(_06809_));
 INV_X1 _12325_ (.A(_06802_),
    .ZN(_06810_));
 AOI22_X1 _12326_ (.A1(_06755_),
    .A2(_06803_),
    .B1(_06809_),
    .B2(_06810_),
    .ZN(_06811_));
 BUF_X1 _12327_ (.A(\dynamic_node_top.south_output.control.planned_f ),
    .Z(_06812_));
 INV_X1 _12328_ (.A(_06812_),
    .ZN(_06813_));
 NAND2_X1 _12329_ (.A1(_05329_),
    .A2(_06598_),
    .ZN(_06814_));
 AOI22_X1 _12330_ (.A1(_05330_),
    .A2(_05820_),
    .B1(_06715_),
    .B2(_05332_),
    .ZN(_06815_));
 AOI21_X1 _12331_ (.A(_05333_),
    .B1(_05789_),
    .B2(_05331_),
    .ZN(_06816_));
 AND2_X1 _12332_ (.A1(_06815_),
    .A2(_06816_),
    .ZN(_06817_));
 AOI22_X4 _12333_ (.A1(_05333_),
    .A2(_06601_),
    .B1(_06814_),
    .B2(_06817_),
    .ZN(_06818_));
 MUX2_X1 _12334_ (.A(_06813_),
    .B(_06818_),
    .S(net1),
    .Z(_06819_));
 BUF_X4 _12335_ (.A(_06819_),
    .Z(_06820_));
 AND3_X1 _12336_ (.A1(_06146_),
    .A2(_06738_),
    .A3(_06179_),
    .ZN(_06821_));
 AND3_X1 _12337_ (.A1(_06786_),
    .A2(_06182_),
    .A3(_06821_),
    .ZN(_06822_));
 NOR2_X1 _12338_ (.A1(_06186_),
    .A2(_06187_),
    .ZN(_06823_));
 NAND2_X1 _12339_ (.A1(_06182_),
    .A2(_06823_),
    .ZN(_06824_));
 INV_X1 _12340_ (.A(_06191_),
    .ZN(_06825_));
 NAND4_X1 _12341_ (.A1(_06146_),
    .A2(_06738_),
    .A3(_06179_),
    .A4(_06825_),
    .ZN(_06826_));
 AOI21_X1 _12342_ (.A(_06824_),
    .B1(_06826_),
    .B2(_06204_),
    .ZN(_06827_));
 MUX2_X2 _12343_ (.A(_06822_),
    .B(_06827_),
    .S(_06492_),
    .Z(_06828_));
 NAND2_X1 _12344_ (.A1(_06820_),
    .A2(_06828_),
    .ZN(_06829_));
 NAND2_X1 _12345_ (.A1(_05329_),
    .A2(_06591_),
    .ZN(_06830_));
 OAI22_X1 _12346_ (.A1(_06811_),
    .A2(_06829_),
    .B1(_06830_),
    .B2(_06820_),
    .ZN(_00031_));
 NAND3_X1 _12347_ (.A1(_06786_),
    .A2(_06163_),
    .A3(_06739_),
    .ZN(_06831_));
 AND2_X1 _12348_ (.A1(_06742_),
    .A2(_06743_),
    .ZN(_06832_));
 MUX2_X2 _12349_ (.A(_06831_),
    .B(_06832_),
    .S(_06492_),
    .Z(_06833_));
 AOI21_X1 _12350_ (.A(_05171_),
    .B1(_05167_),
    .B2(_06765_),
    .ZN(_06834_));
 NOR3_X2 _12351_ (.A1(_05492_),
    .A2(_06546_),
    .A3(_06548_),
    .ZN(_06835_));
 NAND2_X1 _12352_ (.A1(_06786_),
    .A2(_06835_),
    .ZN(_06836_));
 NOR2_X2 _12353_ (.A1(net683),
    .A2(_06565_),
    .ZN(_06837_));
 NAND4_X2 _12354_ (.A1(net639),
    .A2(net715),
    .A3(_05523_),
    .A4(_05518_),
    .ZN(_06838_));
 AOI22_X2 _12355_ (.A1(_06835_),
    .A2(_06837_),
    .B1(_06838_),
    .B2(_05505_),
    .ZN(_06839_));
 MUX2_X1 _12356_ (.A(_06836_),
    .B(_06839_),
    .S(_06567_),
    .Z(_06840_));
 OR2_X2 _12357_ (.A1(_06793_),
    .A2(_06840_),
    .ZN(_06841_));
 NAND2_X1 _12358_ (.A1(_06736_),
    .A2(_06841_),
    .ZN(_06842_));
 OAI21_X1 _12359_ (.A(_06737_),
    .B1(_06834_),
    .B2(_06842_),
    .ZN(_06843_));
 NAND2_X1 _12360_ (.A1(_06758_),
    .A2(_06843_),
    .ZN(_06844_));
 OAI33_X1 _12361_ (.A1(_06718_),
    .A2(_06664_),
    .A3(_06758_),
    .B1(_06833_),
    .B2(_06844_),
    .B3(_06589_),
    .ZN(_00040_));
 NOR2_X1 _12362_ (.A1(_05613_),
    .A2(_06096_),
    .ZN(_06845_));
 NAND4_X1 _12363_ (.A1(_05384_),
    .A2(_05616_),
    .A3(_06100_),
    .A4(_06845_),
    .ZN(_06846_));
 NAND2_X1 _12364_ (.A1(_06103_),
    .A2(_06106_),
    .ZN(_06847_));
 AOI21_X1 _12365_ (.A(_06847_),
    .B1(_06117_),
    .B2(_06113_),
    .ZN(_06848_));
 AND4_X1 _12366_ (.A1(_05616_),
    .A2(_06100_),
    .A3(_06845_),
    .A4(_05627_),
    .ZN(_06849_));
 OAI21_X1 _12367_ (.A(_05630_),
    .B1(_06848_),
    .B2(_06849_),
    .ZN(_06850_));
 MUX2_X2 _12368_ (.A(_06846_),
    .B(_06850_),
    .S(net748),
    .Z(_06851_));
 AND2_X1 _12369_ (.A1(_05329_),
    .A2(_06851_),
    .ZN(_06852_));
 NAND2_X1 _12370_ (.A1(_05452_),
    .A2(_06852_),
    .ZN(_06853_));
 INV_X1 _12371_ (.A(_05338_),
    .ZN(_06854_));
 AOI21_X1 _12372_ (.A(_06541_),
    .B1(_06853_),
    .B2(_06854_),
    .ZN(_06855_));
 INV_X1 _12373_ (.A(net680),
    .ZN(_06856_));
 NOR2_X1 _12374_ (.A1(_06664_),
    .A2(_06856_),
    .ZN(_06857_));
 INV_X4 _12375_ (.A(_05332_),
    .ZN(_06858_));
 BUF_X4 _12376_ (.A(_06858_),
    .Z(_06859_));
 BUF_X4 _12377_ (.A(_06859_),
    .Z(_06860_));
 NAND2_X1 _12378_ (.A1(_05330_),
    .A2(_06851_),
    .ZN(_06861_));
 OAI21_X1 _12379_ (.A(_06860_),
    .B1(_06828_),
    .B2(_06861_),
    .ZN(_06862_));
 AOI21_X1 _12380_ (.A(_06855_),
    .B1(_06857_),
    .B2(_06862_),
    .ZN(_06863_));
 NAND2_X1 _12381_ (.A1(_06567_),
    .A2(_06797_),
    .ZN(_06864_));
 OAI21_X1 _12382_ (.A(_06864_),
    .B1(_06791_),
    .B2(_06567_),
    .ZN(_06865_));
 NAND2_X1 _12383_ (.A1(_06820_),
    .A2(_06865_),
    .ZN(_06866_));
 OAI22_X1 _12384_ (.A1(_06820_),
    .A2(_06804_),
    .B1(_06863_),
    .B2(_06866_),
    .ZN(_00030_));
 AOI21_X1 _12385_ (.A(_06820_),
    .B1(_05756_),
    .B2(_06807_),
    .ZN(_06867_));
 NOR2_X1 _12386_ (.A1(_06812_),
    .A2(net1),
    .ZN(_06868_));
 AOI21_X2 _12387_ (.A(_06868_),
    .B1(_06818_),
    .B2(net1),
    .ZN(_06869_));
 NOR2_X1 _12388_ (.A1(_05329_),
    .A2(_06869_),
    .ZN(_06870_));
 NAND3_X1 _12389_ (.A1(_06786_),
    .A2(_06183_),
    .A3(_06821_),
    .ZN(_06871_));
 NOR2_X1 _12390_ (.A1(_06666_),
    .A2(_06188_),
    .ZN(_06872_));
 AND4_X1 _12391_ (.A1(_06146_),
    .A2(_06738_),
    .A3(_06179_),
    .A4(_06825_),
    .ZN(_06873_));
 INV_X1 _12392_ (.A(_06204_),
    .ZN(_06874_));
 OAI21_X1 _12393_ (.A(_06872_),
    .B1(_06873_),
    .B2(_06874_),
    .ZN(_06875_));
 MUX2_X2 _12394_ (.A(_06871_),
    .B(_06875_),
    .S(_06492_),
    .Z(_06876_));
 AOI21_X2 _12395_ (.A(_05331_),
    .B1(_05338_),
    .B2(_06798_),
    .ZN(_06877_));
 NOR3_X2 _12396_ (.A1(_06541_),
    .A2(_06802_),
    .A3(_06877_),
    .ZN(_06878_));
 OAI21_X1 _12397_ (.A(_06876_),
    .B1(_06878_),
    .B2(_05330_),
    .ZN(_06879_));
 BUF_X4 _12398_ (.A(_06581_),
    .Z(_06880_));
 INV_X1 _12399_ (.A(_06851_),
    .ZN(_06881_));
 NAND2_X1 _12400_ (.A1(_06880_),
    .A2(_06881_),
    .ZN(_06882_));
 AOI221_X1 _12401_ (.A(_06867_),
    .B1(_06870_),
    .B2(_06879_),
    .C1(_06820_),
    .C2(_06882_),
    .ZN(_00028_));
 NOR2_X1 _12402_ (.A1(_06541_),
    .A2(_06877_),
    .ZN(_06883_));
 NOR2_X1 _12403_ (.A1(_06806_),
    .A2(_06852_),
    .ZN(_06884_));
 NOR3_X1 _12404_ (.A1(_06856_),
    .A2(_06805_),
    .A3(_06884_),
    .ZN(_06885_));
 OAI21_X1 _12405_ (.A(_06820_),
    .B1(_06883_),
    .B2(_06885_),
    .ZN(_06886_));
 OAI33_X1 _12406_ (.A1(_06785_),
    .A2(_06664_),
    .A3(_06820_),
    .B1(_06801_),
    .B2(_06886_),
    .B3(_06613_),
    .ZN(_00029_));
 NAND3_X1 _12407_ (.A1(_05167_),
    .A2(_06591_),
    .A3(_06722_),
    .ZN(_06887_));
 NOR2_X1 _12408_ (.A1(_06572_),
    .A2(_06752_),
    .ZN(_06888_));
 NAND3_X1 _12409_ (.A1(_05171_),
    .A2(_06736_),
    .A3(_06841_),
    .ZN(_06889_));
 AOI21_X1 _12410_ (.A(_06745_),
    .B1(_06889_),
    .B2(_06737_),
    .ZN(_06890_));
 OAI21_X1 _12411_ (.A(_06888_),
    .B1(_06890_),
    .B2(_05158_),
    .ZN(_06891_));
 OAI21_X1 _12412_ (.A(_06887_),
    .B1(_06891_),
    .B2(_06722_),
    .ZN(_00039_));
 BUF_X4 _12413_ (.A(_06755_),
    .Z(_06892_));
 NOR2_X1 _12414_ (.A1(_06828_),
    .A2(_06881_),
    .ZN(_06893_));
 AND2_X1 _12415_ (.A1(_05338_),
    .A2(_05756_),
    .ZN(_06894_));
 OAI211_X2 _12416_ (.A(_06893_),
    .B(_06878_),
    .C1(_06894_),
    .C2(_06820_),
    .ZN(_06895_));
 NAND3_X1 _12417_ (.A1(_05332_),
    .A2(_05452_),
    .A3(_06801_),
    .ZN(_06896_));
 NAND3_X1 _12418_ (.A1(_05332_),
    .A2(_05185_),
    .A3(_05452_),
    .ZN(_06897_));
 AND2_X1 _12419_ (.A1(_06861_),
    .A2(_06897_),
    .ZN(_06898_));
 AOI221_X2 _12420_ (.A(_06828_),
    .B1(_06896_),
    .B2(_06898_),
    .C1(_06805_),
    .C2(net680),
    .ZN(_06899_));
 NOR3_X1 _12421_ (.A1(_06802_),
    .A2(_06805_),
    .A3(_06853_),
    .ZN(_06900_));
 AOI21_X1 _12422_ (.A(_06806_),
    .B1(_05755_),
    .B2(_06852_),
    .ZN(_06901_));
 NOR2_X1 _12423_ (.A1(net680),
    .A2(_06901_),
    .ZN(_06902_));
 NOR4_X2 _12424_ (.A1(_06869_),
    .A2(_06899_),
    .A3(_06900_),
    .A4(_06902_),
    .ZN(_06903_));
 NOR2_X1 _12425_ (.A1(_06820_),
    .A2(_06894_),
    .ZN(_06904_));
 OAI211_X2 _12426_ (.A(_06892_),
    .B(_06895_),
    .C1(_06903_),
    .C2(_06904_),
    .ZN(_00027_));
 OR2_X1 _12427_ (.A1(_05492_),
    .A2(_05500_),
    .ZN(_06905_));
 NOR3_X2 _12428_ (.A1(_05489_),
    .A2(_06546_),
    .A3(_06905_),
    .ZN(_06906_));
 MUX2_X1 _12429_ (.A(_06786_),
    .B(_06837_),
    .S(_06567_),
    .Z(_06907_));
 NAND2_X1 _12430_ (.A1(_06906_),
    .A2(_06907_),
    .ZN(_06908_));
 CLKBUF_X3 _12431_ (.A(_05346_),
    .Z(_06909_));
 NOR2_X1 _12432_ (.A1(_05372_),
    .A2(_05374_),
    .ZN(_06910_));
 NOR3_X2 _12433_ (.A1(_06909_),
    .A2(_06910_),
    .A3(_06619_),
    .ZN(_06911_));
 INV_X1 _12434_ (.A(_06749_),
    .ZN(_06912_));
 MUX2_X1 _12435_ (.A(_06786_),
    .B(_06912_),
    .S(_06523_),
    .Z(_06913_));
 AND2_X2 _12436_ (.A1(_06911_),
    .A2(_06913_),
    .ZN(_06914_));
 INV_X1 _12437_ (.A(_05595_),
    .ZN(_06915_));
 BUF_X4 _12438_ (.A(_05596_),
    .Z(_06916_));
 NOR3_X2 _12439_ (.A1(_05185_),
    .A2(_05273_),
    .A3(_06514_),
    .ZN(_06917_));
 NAND3_X1 _12440_ (.A1(_06513_),
    .A2(_06786_),
    .A3(_06917_),
    .ZN(_06918_));
 NAND4_X1 _12441_ (.A1(_05266_),
    .A2(_05269_),
    .A3(_06513_),
    .A4(_06917_),
    .ZN(_06919_));
 MUX2_X2 _12442_ (.A(_06918_),
    .B(_06919_),
    .S(_05263_),
    .Z(_06920_));
 NAND3_X1 _12443_ (.A1(_06916_),
    .A2(_05696_),
    .A3(_06920_),
    .ZN(_06921_));
 AND2_X1 _12444_ (.A1(_06915_),
    .A2(_06921_),
    .ZN(_06922_));
 OR3_X1 _12445_ (.A1(_06663_),
    .A2(_06914_),
    .A3(_06922_),
    .ZN(_06923_));
 INV_X1 _12446_ (.A(_05603_),
    .ZN(_06924_));
 INV_X1 _12447_ (.A(_06917_),
    .ZN(_06925_));
 NOR3_X4 _12448_ (.A1(_05277_),
    .A2(_06616_),
    .A3(_06925_),
    .ZN(_06926_));
 NOR3_X1 _12449_ (.A1(_06924_),
    .A2(_06914_),
    .A3(_06926_),
    .ZN(_06927_));
 OAI21_X1 _12450_ (.A(_06880_),
    .B1(_06927_),
    .B2(_05594_),
    .ZN(_06928_));
 AOI21_X1 _12451_ (.A(_06908_),
    .B1(_06923_),
    .B2(_06928_),
    .ZN(_06929_));
 AND2_X1 _12452_ (.A1(_05605_),
    .A2(_05756_),
    .ZN(_06930_));
 BUF_X1 _12453_ (.A(\dynamic_node_top.proc_output.control.planned_f ),
    .Z(_06931_));
 NOR2_X1 _12454_ (.A1(_06931_),
    .A2(net744),
    .ZN(_06932_));
 OAI21_X1 _12455_ (.A(_05605_),
    .B1(_05786_),
    .B2(_05788_),
    .ZN(_06933_));
 INV_X1 _12456_ (.A(_05594_),
    .ZN(_06934_));
 OAI221_X2 _12457_ (.A(_06933_),
    .B1(_06713_),
    .B2(_06915_),
    .C1(_06934_),
    .C2(_06601_),
    .ZN(_06935_));
 AOI211_X2 _12458_ (.A(_05597_),
    .B(_06935_),
    .C1(_06598_),
    .C2(_05596_),
    .ZN(_06936_));
 NOR2_X2 _12459_ (.A1(_05598_),
    .A2(_06715_),
    .ZN(_06937_));
 NOR2_X2 _12460_ (.A1(_06936_),
    .A2(_06937_),
    .ZN(_06938_));
 AOI21_X4 _12461_ (.A(_06932_),
    .B1(_06938_),
    .B2(net744),
    .ZN(_06939_));
 MUX2_X1 _12462_ (.A(_06929_),
    .B(_06930_),
    .S(_06939_),
    .Z(_00026_));
 AND3_X1 _12463_ (.A1(_05595_),
    .A2(_05756_),
    .A3(_06939_),
    .ZN(_06940_));
 NAND2_X1 _12464_ (.A1(_06581_),
    .A2(_06926_),
    .ZN(_06941_));
 AOI21_X1 _12465_ (.A(_05603_),
    .B1(_06916_),
    .B2(_05696_),
    .ZN(_06942_));
 INV_X1 _12466_ (.A(_06672_),
    .ZN(_06943_));
 MUX2_X2 _12467_ (.A(_05304_),
    .B(_06943_),
    .S(_06492_),
    .Z(_06944_));
 NAND2_X2 _12468_ (.A1(_06738_),
    .A2(_06739_),
    .ZN(_06945_));
 NAND2_X1 _12469_ (.A1(_06786_),
    .A2(_06906_),
    .ZN(_06946_));
 NAND2_X1 _12470_ (.A1(_06837_),
    .A2(_06906_),
    .ZN(_06947_));
 MUX2_X1 _12471_ (.A(_06946_),
    .B(_06947_),
    .S(_06567_),
    .Z(_06948_));
 AND2_X1 _12472_ (.A1(_05594_),
    .A2(_06948_),
    .ZN(_06949_));
 OAI221_X2 _12473_ (.A(_05696_),
    .B1(_06944_),
    .B2(_06945_),
    .C1(_06949_),
    .C2(_05605_),
    .ZN(_06950_));
 AOI211_X2 _12474_ (.A(_06939_),
    .B(_06941_),
    .C1(_06942_),
    .C2(_06950_),
    .ZN(_06951_));
 OR2_X1 _12475_ (.A1(_06940_),
    .A2(_06951_),
    .ZN(_00025_));
 AND2_X1 _12476_ (.A1(_05173_),
    .A2(_05756_),
    .ZN(_06952_));
 AOI21_X1 _12477_ (.A(_06573_),
    .B1(_06722_),
    .B2(_06952_),
    .ZN(_06953_));
 NAND3_X1 _12478_ (.A1(_06752_),
    .A2(_06765_),
    .A3(_06841_),
    .ZN(_06954_));
 NOR2_X1 _12479_ (.A1(_06718_),
    .A2(_06954_),
    .ZN(_06955_));
 INV_X1 _12480_ (.A(_05167_),
    .ZN(_06956_));
 NOR4_X1 _12481_ (.A1(_06956_),
    .A2(_06540_),
    .A3(_06763_),
    .A4(_06764_),
    .ZN(_06957_));
 OAI21_X1 _12482_ (.A(_06841_),
    .B1(_06957_),
    .B2(_05171_),
    .ZN(_06958_));
 INV_X2 _12483_ (.A(_05159_),
    .ZN(_06959_));
 BUF_X4 _12484_ (.A(_06959_),
    .Z(_06960_));
 AOI21_X1 _12485_ (.A(_06736_),
    .B1(_06958_),
    .B2(_06960_),
    .ZN(_06961_));
 AOI22_X1 _12486_ (.A1(_05171_),
    .A2(_06752_),
    .B1(_06765_),
    .B2(_05167_),
    .ZN(_06962_));
 AOI22_X1 _12487_ (.A1(_05159_),
    .A2(_06736_),
    .B1(_06841_),
    .B2(_05173_),
    .ZN(_06963_));
 INV_X1 _12488_ (.A(_06752_),
    .ZN(_06964_));
 OAI33_X1 _12489_ (.A1(_06541_),
    .A2(_06842_),
    .A3(_06962_),
    .B1(_06963_),
    .B2(_06766_),
    .B3(_06964_),
    .ZN(_06965_));
 AOI211_X2 _12490_ (.A(_06955_),
    .B(_06961_),
    .C1(_06965_),
    .C2(_06833_),
    .ZN(_06966_));
 OAI21_X1 _12491_ (.A(_06953_),
    .B1(_06966_),
    .B2(_06722_),
    .ZN(_00037_));
 NAND3_X1 _12492_ (.A1(_05594_),
    .A2(_06591_),
    .A3(_06939_),
    .ZN(_06967_));
 NAND3_X1 _12493_ (.A1(_05603_),
    .A2(_05755_),
    .A3(_06920_),
    .ZN(_06968_));
 OAI21_X1 _12494_ (.A(_06968_),
    .B1(_06922_),
    .B2(_06572_),
    .ZN(_06969_));
 AND4_X1 _12495_ (.A1(_05605_),
    .A2(_05756_),
    .A3(_05696_),
    .A4(_06920_),
    .ZN(_06970_));
 OR2_X1 _12496_ (.A1(_06944_),
    .A2(_06945_),
    .ZN(_06971_));
 AOI21_X1 _12497_ (.A(_06969_),
    .B1(_06970_),
    .B2(_06971_),
    .ZN(_06972_));
 NAND2_X1 _12498_ (.A1(_06786_),
    .A2(_06911_),
    .ZN(_06973_));
 NAND2_X1 _12499_ (.A1(_06912_),
    .A2(_06911_),
    .ZN(_06974_));
 MUX2_X1 _12500_ (.A(_06973_),
    .B(_06974_),
    .S(_06523_),
    .Z(_06975_));
 OR2_X1 _12501_ (.A1(_06939_),
    .A2(_06975_),
    .ZN(_06976_));
 OAI21_X1 _12502_ (.A(_06967_),
    .B1(_06972_),
    .B2(_06976_),
    .ZN(_00024_));
 BUF_X4 _12503_ (.A(_06916_),
    .Z(_06977_));
 NAND3_X1 _12504_ (.A1(_06977_),
    .A2(_06591_),
    .A3(_06939_),
    .ZN(_06978_));
 AOI21_X1 _12505_ (.A(_05595_),
    .B1(_05603_),
    .B2(_06920_),
    .ZN(_06979_));
 OAI21_X1 _12506_ (.A(_06934_),
    .B1(_06914_),
    .B2(_06979_),
    .ZN(_06980_));
 AOI21_X1 _12507_ (.A(_05605_),
    .B1(_06908_),
    .B2(_06980_),
    .ZN(_06981_));
 OR3_X1 _12508_ (.A1(_06572_),
    .A2(_06971_),
    .A3(_06981_),
    .ZN(_06982_));
 OAI21_X1 _12509_ (.A(_06978_),
    .B1(_06982_),
    .B2(_06939_),
    .ZN(_00023_));
 NOR2_X1 _12510_ (.A1(_06924_),
    .A2(_06664_),
    .ZN(_06983_));
 AOI21_X1 _12511_ (.A(_06573_),
    .B1(_06939_),
    .B2(_06983_),
    .ZN(_06984_));
 NOR2_X1 _12512_ (.A1(_05304_),
    .A2(_05624_),
    .ZN(_06985_));
 NOR2_X1 _12513_ (.A1(_05624_),
    .A2(_05631_),
    .ZN(_06986_));
 MUX2_X2 _12514_ (.A(_06985_),
    .B(_06986_),
    .S(net748),
    .Z(_06987_));
 AND2_X1 _12515_ (.A1(_06906_),
    .A2(_06907_),
    .ZN(_06988_));
 NOR3_X1 _12516_ (.A1(_06914_),
    .A2(_06926_),
    .A3(_06988_),
    .ZN(_06989_));
 OR2_X1 _12517_ (.A1(_06987_),
    .A2(_06989_),
    .ZN(_06990_));
 AOI21_X1 _12518_ (.A(_06987_),
    .B1(_06920_),
    .B2(_06581_),
    .ZN(_06991_));
 NOR3_X1 _12519_ (.A1(_06987_),
    .A2(_06975_),
    .A3(_06949_),
    .ZN(_06992_));
 NOR2_X1 _12520_ (.A1(_05605_),
    .A2(_06949_),
    .ZN(_06993_));
 OAI33_X1 _12521_ (.A1(_06914_),
    .A2(_06988_),
    .A3(_06979_),
    .B1(_06991_),
    .B2(_06992_),
    .B3(_06993_),
    .ZN(_06994_));
 AOI22_X1 _12522_ (.A1(_06916_),
    .A2(_06990_),
    .B1(_06994_),
    .B2(_06971_),
    .ZN(_06995_));
 OAI21_X1 _12523_ (.A(_06984_),
    .B1(_06995_),
    .B2(_06939_),
    .ZN(_00022_));
 BUF_X4 _12524_ (.A(_06724_),
    .Z(_06996_));
 NAND3_X1 _12525_ (.A1(_06996_),
    .A2(_06591_),
    .A3(_06722_),
    .ZN(_06997_));
 NAND3_X1 _12526_ (.A1(_05158_),
    .A2(_06752_),
    .A3(_06765_),
    .ZN(_06998_));
 INV_X1 _12527_ (.A(_05171_),
    .ZN(_06999_));
 AOI21_X1 _12528_ (.A(_06572_),
    .B1(_06998_),
    .B2(_06999_),
    .ZN(_07000_));
 NOR2_X1 _12529_ (.A1(_06664_),
    .A2(_06766_),
    .ZN(_07001_));
 NAND2_X1 _12530_ (.A1(_05173_),
    .A2(_06752_),
    .ZN(_07002_));
 OAI21_X1 _12531_ (.A(_06956_),
    .B1(_06745_),
    .B2(_07002_),
    .ZN(_07003_));
 AOI21_X1 _12532_ (.A(_07000_),
    .B1(_07001_),
    .B2(_07003_),
    .ZN(_07004_));
 OR2_X1 _12533_ (.A1(_06722_),
    .A2(_06841_),
    .ZN(_07005_));
 OAI21_X1 _12534_ (.A(_06997_),
    .B1(_07004_),
    .B2(_07005_),
    .ZN(_00038_));
 NAND3_X1 _12535_ (.A1(_05757_),
    .A2(_06591_),
    .A3(_06127_),
    .ZN(_07006_));
 OAI21_X1 _12536_ (.A(_05857_),
    .B1(_06493_),
    .B2(_06519_),
    .ZN(_07007_));
 NAND2_X1 _12537_ (.A1(_05754_),
    .A2(net667),
    .ZN(_07008_));
 OAI21_X1 _12538_ (.A(_06520_),
    .B1(_06574_),
    .B2(_07008_),
    .ZN(_07009_));
 NOR2_X1 _12539_ (.A1(_06664_),
    .A2(_06493_),
    .ZN(_07010_));
 AOI22_X1 _12540_ (.A1(_06755_),
    .A2(_07007_),
    .B1(_07009_),
    .B2(_07010_),
    .ZN(_07011_));
 OR2_X1 _12541_ (.A1(_06127_),
    .A2(_06568_),
    .ZN(_07012_));
 OAI21_X1 _12542_ (.A(_07006_),
    .B1(_07011_),
    .B2(_07012_),
    .ZN(_00021_));
 NOR4_X1 _12543_ (.A1(_06603_),
    .A2(_06607_),
    .A3(_06636_),
    .A4(_06697_),
    .ZN(_07013_));
 AOI21_X1 _12544_ (.A(_07013_),
    .B1(_06607_),
    .B2(_05478_),
    .ZN(_07014_));
 BUF_X4 _12545_ (.A(_06609_),
    .Z(_07015_));
 AOI21_X1 _12546_ (.A(_05481_),
    .B1(_07015_),
    .B2(net702),
    .ZN(_07016_));
 NOR3_X1 _12547_ (.A1(_06660_),
    .A2(_06697_),
    .A3(_07016_),
    .ZN(_07017_));
 OAI21_X1 _12548_ (.A(_06661_),
    .B1(_07017_),
    .B2(_05484_),
    .ZN(_07018_));
 OAI22_X1 _12549_ (.A1(_06664_),
    .A2(_07014_),
    .B1(_07018_),
    .B2(_06636_),
    .ZN(_00036_));
 NAND3_X1 _12550_ (.A1(_05821_),
    .A2(_06591_),
    .A3(_06127_),
    .ZN(_07019_));
 NOR2_X1 _12551_ (.A1(_06515_),
    .A2(_06517_),
    .ZN(_07020_));
 OR3_X2 _12552_ (.A1(_06613_),
    .A2(_06510_),
    .A3(_07020_),
    .ZN(_07021_));
 INV_X2 _12553_ (.A(_05753_),
    .ZN(_07022_));
 AOI21_X1 _12554_ (.A(_05757_),
    .B1(_05823_),
    .B2(_06568_),
    .ZN(_07023_));
 OAI21_X1 _12555_ (.A(_07022_),
    .B1(_06538_),
    .B2(_07023_),
    .ZN(_07024_));
 AOI21_X1 _12556_ (.A(_06090_),
    .B1(net667),
    .B2(_07024_),
    .ZN(_07025_));
 OR4_X1 _12557_ (.A1(_06572_),
    .A2(_06127_),
    .A3(_07021_),
    .A4(_07025_),
    .ZN(_07026_));
 NAND2_X1 _12558_ (.A1(_07019_),
    .A2(_07026_),
    .ZN(_00020_));
 NAND3_X1 _12559_ (.A1(_05823_),
    .A2(_06591_),
    .A3(_06127_),
    .ZN(_07027_));
 INV_X1 _12560_ (.A(_06090_),
    .ZN(_07028_));
 NAND2_X1 _12561_ (.A1(_06576_),
    .A2(_06578_),
    .ZN(_07029_));
 NAND3_X1 _12562_ (.A1(_07028_),
    .A2(_07029_),
    .A3(_07008_),
    .ZN(_07030_));
 AOI21_X1 _12563_ (.A(_05821_),
    .B1(_07021_),
    .B2(_07030_),
    .ZN(_07031_));
 NOR3_X1 _12564_ (.A1(_05383_),
    .A2(_06147_),
    .A3(_06180_),
    .ZN(_07032_));
 NOR2_X1 _12565_ (.A1(_05303_),
    .A2(_06666_),
    .ZN(_07033_));
 OAI21_X1 _12566_ (.A(_05300_),
    .B1(_07032_),
    .B2(_07033_),
    .ZN(_07034_));
 NOR3_X1 _12567_ (.A1(_06147_),
    .A2(_06180_),
    .A3(_06191_),
    .ZN(_07035_));
 AND3_X1 _12568_ (.A1(_06182_),
    .A2(_06191_),
    .A3(_06204_),
    .ZN(_07036_));
 OAI21_X1 _12569_ (.A(_06823_),
    .B1(_07035_),
    .B2(_07036_),
    .ZN(_07037_));
 MUX2_X2 _12570_ (.A(_07034_),
    .B(_07037_),
    .S(_06492_),
    .Z(_07038_));
 OR3_X1 _12571_ (.A1(_06572_),
    .A2(_06127_),
    .A3(_07038_),
    .ZN(_07039_));
 OAI21_X1 _12572_ (.A(_07027_),
    .B1(_07031_),
    .B2(_07039_),
    .ZN(_00019_));
 NOR4_X2 _12573_ (.A1(_05605_),
    .A2(_05594_),
    .A3(_05603_),
    .A4(_06916_),
    .ZN(_07040_));
 AOI22_X2 _12574_ (.A1(_05479_),
    .A2(net756),
    .B1(net623),
    .B2(_07040_),
    .ZN(_07041_));
 OAI21_X2 _12575_ (.A(_07041_),
    .B1(_05308_),
    .B2(_05161_),
    .ZN(_07042_));
 NOR2_X1 _12576_ (.A1(_05338_),
    .A2(_05332_),
    .ZN(_07043_));
 NAND2_X2 _12577_ (.A1(net624),
    .A2(_07043_),
    .ZN(_07044_));
 NAND3_X2 _12578_ (.A1(_07028_),
    .A2(net622),
    .A3(_07022_),
    .ZN(_07045_));
 OAI33_X1 _12579_ (.A1(_05329_),
    .A2(_05331_),
    .A3(_07044_),
    .B1(_07045_),
    .B2(_05757_),
    .B3(_05823_),
    .ZN(_07046_));
 NOR2_X4 _12580_ (.A1(_07042_),
    .A2(_07046_),
    .ZN(_10498_));
 INV_X1 _12581_ (.A(_10498_),
    .ZN(\dynamic_node_top.west_input.NIB.thanks_in ));
 XOR2_X1 _12582_ (.A(_05818_),
    .B(\dynamic_node_top.west_input.control.count_f[0] ),
    .Z(_07047_));
 MUX2_X1 _12583_ (.A(_05815_),
    .B(_07047_),
    .S(_06613_),
    .Z(_07048_));
 BUF_X1 _12584_ (.A(\dynamic_node_top.west_input.control.count_f[2] ),
    .Z(_07049_));
 NAND2_X1 _12585_ (.A1(_05818_),
    .A2(_10481_),
    .ZN(_07050_));
 OR3_X1 _12586_ (.A1(_07049_),
    .A2(\dynamic_node_top.west_input.control.count_f[3] ),
    .A3(_07050_),
    .ZN(_07051_));
 XNOR2_X1 _12587_ (.A(\dynamic_node_top.west_input.control.count_f[4] ),
    .B(_07051_),
    .ZN(_07052_));
 NOR2_X1 _12588_ (.A1(_06701_),
    .A2(_07052_),
    .ZN(_07053_));
 INV_X1 _12589_ (.A(_05818_),
    .ZN(_07054_));
 OR4_X1 _12590_ (.A1(_07054_),
    .A2(\dynamic_node_top.west_input.control.count_f[0] ),
    .A3(\dynamic_node_top.west_input.control.count_f[1] ),
    .A4(_07049_),
    .ZN(_07055_));
 XNOR2_X1 _12591_ (.A(\dynamic_node_top.west_input.control.count_f[3] ),
    .B(_07055_),
    .ZN(_07056_));
 OR3_X1 _12592_ (.A1(_05818_),
    .A2(\dynamic_node_top.west_input.control.count_f[1] ),
    .A3(_07049_),
    .ZN(_07057_));
 XNOR2_X1 _12593_ (.A(_10481_),
    .B(_07049_),
    .ZN(_07058_));
 NAND3_X1 _12594_ (.A1(_05818_),
    .A2(_10482_),
    .A3(_07058_),
    .ZN(_07059_));
 AOI21_X1 _12595_ (.A(_07056_),
    .B1(_07057_),
    .B2(_07059_),
    .ZN(_07060_));
 AOI22_X2 _12596_ (.A1(_05793_),
    .A2(_05803_),
    .B1(_07053_),
    .B2(_07060_),
    .ZN(_07061_));
 OR3_X1 _12597_ (.A1(\dynamic_node_top.west_input.control.count_f[3] ),
    .A2(\dynamic_node_top.west_input.control.count_f[4] ),
    .A3(_07055_),
    .ZN(_07062_));
 NOR3_X1 _12598_ (.A1(\dynamic_node_top.west_input.control.count_f[5] ),
    .A2(\dynamic_node_top.west_input.control.count_f[6] ),
    .A3(_07062_),
    .ZN(_07063_));
 XOR2_X1 _12599_ (.A(\dynamic_node_top.west_input.control.count_f[7] ),
    .B(_07063_),
    .Z(_07064_));
 MUX2_X1 _12600_ (.A(_05812_),
    .B(_07064_),
    .S(_06613_),
    .Z(_07065_));
 NOR3_X1 _12601_ (.A1(\dynamic_node_top.west_input.control.count_f[4] ),
    .A2(\dynamic_node_top.west_input.control.count_f[5] ),
    .A3(_07051_),
    .ZN(_07066_));
 XNOR2_X1 _12602_ (.A(\dynamic_node_top.west_input.control.count_f[6] ),
    .B(_07066_),
    .ZN(_07067_));
 NOR2_X1 _12603_ (.A1(_06701_),
    .A2(_07067_),
    .ZN(_07068_));
 AOI21_X1 _12604_ (.A(_07068_),
    .B1(_05806_),
    .B2(_06701_),
    .ZN(_07069_));
 XOR2_X1 _12605_ (.A(\dynamic_node_top.west_input.control.count_f[5] ),
    .B(_07062_),
    .Z(_07070_));
 NOR2_X1 _12606_ (.A1(_06701_),
    .A2(_07070_),
    .ZN(_07071_));
 AOI21_X1 _12607_ (.A(_07071_),
    .B1(_05809_),
    .B2(_06701_),
    .ZN(_07072_));
 NAND2_X1 _12608_ (.A1(_07069_),
    .A2(_07072_),
    .ZN(_07073_));
 NOR4_X1 _12609_ (.A1(_07048_),
    .A2(_07061_),
    .A3(_07065_),
    .A4(_07073_),
    .ZN(_07074_));
 OR2_X1 _12610_ (.A1(_06572_),
    .A2(_07074_),
    .ZN(_07075_));
 OR2_X1 _12611_ (.A1(\dynamic_node_top.west_input.control.header_last_temp ),
    .A2(_06572_),
    .ZN(_07076_));
 MUX2_X1 _12612_ (.A(_07075_),
    .B(_07076_),
    .S(_10498_),
    .Z(_00004_));
 OR2_X1 _12613_ (.A1(_05173_),
    .A2(_05159_),
    .ZN(_07077_));
 OR2_X1 _12614_ (.A1(_05171_),
    .A2(_07077_),
    .ZN(_07078_));
 NOR3_X2 _12615_ (.A1(_05158_),
    .A2(_05308_),
    .A3(_07078_),
    .ZN(_07079_));
 AOI22_X1 _12616_ (.A1(_05333_),
    .A2(net624),
    .B1(net622),
    .B2(_05753_),
    .ZN(_07080_));
 INV_X1 _12617_ (.A(_07080_),
    .ZN(_07081_));
 INV_X4 _12618_ (.A(_06916_),
    .ZN(_07082_));
 NAND4_X2 _12619_ (.A1(_06915_),
    .A2(_06924_),
    .A3(_07082_),
    .A4(net623),
    .ZN(_07083_));
 NOR3_X1 _12620_ (.A1(_05484_),
    .A2(_05481_),
    .A3(_05471_),
    .ZN(_07084_));
 NAND2_X2 _12621_ (.A1(net625),
    .A2(_07084_),
    .ZN(_07085_));
 OAI22_X4 _12622_ (.A1(_05605_),
    .A2(_07083_),
    .B1(_07085_),
    .B2(_05470_),
    .ZN(_07086_));
 NOR3_X4 _12623_ (.A1(_07079_),
    .A2(_07081_),
    .A3(_07086_),
    .ZN(_10472_));
 INV_X1 _12624_ (.A(_10472_),
    .ZN(\dynamic_node_top.north_input.NIB.thanks_in ));
 XOR2_X1 _12625_ (.A(_05825_),
    .B(\dynamic_node_top.north_input.control.count_f[0] ),
    .Z(_07087_));
 MUX2_X1 _12626_ (.A(_05846_),
    .B(_07087_),
    .S(_06909_),
    .Z(_07088_));
 NOR2_X1 _12627_ (.A1(_05825_),
    .A2(\dynamic_node_top.north_input.control.count_f[1] ),
    .ZN(_07089_));
 AOI21_X1 _12628_ (.A(_07089_),
    .B1(_10423_),
    .B2(_05825_),
    .ZN(_07090_));
 MUX2_X1 _12629_ (.A(_05849_),
    .B(_07090_),
    .S(_06909_),
    .Z(_07091_));
 NAND2_X1 _12630_ (.A1(_05825_),
    .A2(_10422_),
    .ZN(_07092_));
 XNOR2_X1 _12631_ (.A(\dynamic_node_top.north_input.control.count_f[2] ),
    .B(_07092_),
    .ZN(_07093_));
 MUX2_X1 _12632_ (.A(_05839_),
    .B(_07093_),
    .S(_06909_),
    .Z(_07094_));
 INV_X1 _12633_ (.A(_05825_),
    .ZN(_07095_));
 NOR4_X1 _12634_ (.A1(_07095_),
    .A2(\dynamic_node_top.north_input.control.count_f[0] ),
    .A3(\dynamic_node_top.north_input.control.count_f[1] ),
    .A4(\dynamic_node_top.north_input.control.count_f[2] ),
    .ZN(_07096_));
 XOR2_X1 _12635_ (.A(\dynamic_node_top.north_input.control.count_f[3] ),
    .B(_07096_),
    .Z(_07097_));
 INV_X1 _12636_ (.A(_07097_),
    .ZN(_07098_));
 NOR2_X1 _12637_ (.A1(\dynamic_node_top.north_input.control.count_f[2] ),
    .A2(\dynamic_node_top.north_input.control.count_f[3] ),
    .ZN(_07099_));
 NAND3_X1 _12638_ (.A1(_05825_),
    .A2(_10422_),
    .A3(_07099_),
    .ZN(_07100_));
 XNOR2_X1 _12639_ (.A(\dynamic_node_top.north_input.control.count_f[4] ),
    .B(_07100_),
    .ZN(_07101_));
 NOR2_X1 _12640_ (.A1(_05386_),
    .A2(_07101_),
    .ZN(_07102_));
 AOI21_X1 _12641_ (.A(_05833_),
    .B1(_07098_),
    .B2(_07102_),
    .ZN(_07103_));
 NOR3_X1 _12642_ (.A1(_07091_),
    .A2(_07094_),
    .A3(_07103_),
    .ZN(_07104_));
 INV_X2 _12643_ (.A(_05852_),
    .ZN(_07105_));
 INV_X1 _12644_ (.A(\dynamic_node_top.north_input.control.count_f[4] ),
    .ZN(_07106_));
 NOR3_X1 _12645_ (.A1(_07095_),
    .A2(\dynamic_node_top.north_input.control.count_f[0] ),
    .A3(\dynamic_node_top.north_input.control.count_f[1] ),
    .ZN(_07107_));
 NAND3_X1 _12646_ (.A1(_07106_),
    .A2(_07107_),
    .A3(_07099_),
    .ZN(_07108_));
 NOR3_X1 _12647_ (.A1(\dynamic_node_top.north_input.control.count_f[5] ),
    .A2(\dynamic_node_top.north_input.control.count_f[6] ),
    .A3(_07108_),
    .ZN(_07109_));
 XNOR2_X1 _12648_ (.A(\dynamic_node_top.north_input.control.count_f[7] ),
    .B(_07109_),
    .ZN(_07110_));
 MUX2_X1 _12649_ (.A(_07105_),
    .B(_07110_),
    .S(_06909_),
    .Z(_07111_));
 NOR3_X1 _12650_ (.A1(\dynamic_node_top.north_input.control.count_f[4] ),
    .A2(\dynamic_node_top.north_input.control.count_f[5] ),
    .A3(_07100_),
    .ZN(_07112_));
 XNOR2_X1 _12651_ (.A(\dynamic_node_top.north_input.control.count_f[6] ),
    .B(_07112_),
    .ZN(_07113_));
 NOR2_X1 _12652_ (.A1(_05386_),
    .A2(_07113_),
    .ZN(_07114_));
 AOI21_X1 _12653_ (.A(_07114_),
    .B1(_05843_),
    .B2(_05386_),
    .ZN(_07115_));
 XOR2_X1 _12654_ (.A(\dynamic_node_top.north_input.control.count_f[5] ),
    .B(_07108_),
    .Z(_07116_));
 NOR2_X1 _12655_ (.A1(_05386_),
    .A2(_07116_),
    .ZN(_07117_));
 AOI21_X1 _12656_ (.A(_07117_),
    .B1(_05836_),
    .B2(_05386_),
    .ZN(_07118_));
 NAND4_X1 _12657_ (.A1(_07104_),
    .A2(_07111_),
    .A3(_07115_),
    .A4(_07118_),
    .ZN(_07119_));
 OAI21_X1 _12658_ (.A(_06880_),
    .B1(_07088_),
    .B2(_07119_),
    .ZN(_07120_));
 OR2_X1 _12659_ (.A1(\dynamic_node_top.north_input.control.header_last_temp ),
    .A2(_06541_),
    .ZN(_07121_));
 MUX2_X1 _12660_ (.A(_07120_),
    .B(_07121_),
    .S(_10472_),
    .Z(_00001_));
 NOR4_X1 _12661_ (.A1(_05478_),
    .A2(_05470_),
    .A3(_05481_),
    .A4(_06609_),
    .ZN(_07122_));
 AND2_X4 _12662_ (.A1(net625),
    .A2(_07122_),
    .ZN(_07123_));
 INV_X1 _12663_ (.A(_05697_),
    .ZN(_07124_));
 NOR2_X1 _12664_ (.A1(_07124_),
    .A2(_06987_),
    .ZN(_07125_));
 OAI33_X1 _12665_ (.A1(_00053_),
    .A2(_05610_),
    .A3(_07125_),
    .B1(_05330_),
    .B2(_07044_),
    .B3(_05331_),
    .ZN(_07126_));
 OAI33_X1 _12666_ (.A1(_07045_),
    .A2(_05821_),
    .A3(_05757_),
    .B1(_05167_),
    .B2(_05308_),
    .B3(_07078_),
    .ZN(_07127_));
 NOR3_X4 _12667_ (.A1(_07126_),
    .A2(_07123_),
    .A3(_07127_),
    .ZN(_10456_));
 INV_X2 _12668_ (.A(_10456_),
    .ZN(net620));
 XNOR2_X1 _12669_ (.A(_05858_),
    .B(\dynamic_node_top.proc_input.control.count_f[0] ),
    .ZN(_07128_));
 NOR2_X1 _12670_ (.A1(_06183_),
    .A2(_07128_),
    .ZN(_07129_));
 BUF_X4 _12671_ (.A(_06009_),
    .Z(_07130_));
 NOR2_X1 _12672_ (.A1(_07130_),
    .A2(_06027_),
    .ZN(_07131_));
 AOI21_X4 _12673_ (.A(_07131_),
    .B1(_06047_),
    .B2(_07130_),
    .ZN(_07132_));
 AOI21_X2 _12674_ (.A(_07129_),
    .B1(_07132_),
    .B2(_06183_),
    .ZN(_07133_));
 INV_X1 _12675_ (.A(_07133_),
    .ZN(_07134_));
 NAND2_X1 _12676_ (.A1(_05858_),
    .A2(_10533_),
    .ZN(_07135_));
 XOR2_X1 _12677_ (.A(\dynamic_node_top.proc_input.control.count_f[2] ),
    .B(_07135_),
    .Z(_07136_));
 NOR2_X1 _12678_ (.A1(_06183_),
    .A2(_07136_),
    .ZN(_07137_));
 AOI21_X1 _12679_ (.A(_07137_),
    .B1(_05956_),
    .B2(_06183_),
    .ZN(_07138_));
 OR3_X1 _12680_ (.A1(\dynamic_node_top.proc_input.control.count_f[2] ),
    .A2(\dynamic_node_top.proc_input.control.count_f[3] ),
    .A3(_07135_),
    .ZN(_07139_));
 NOR3_X1 _12681_ (.A1(\dynamic_node_top.proc_input.control.count_f[4] ),
    .A2(\dynamic_node_top.proc_input.control.count_f[5] ),
    .A3(_07139_),
    .ZN(_07140_));
 XNOR2_X1 _12682_ (.A(\dynamic_node_top.proc_input.control.count_f[6] ),
    .B(_07140_),
    .ZN(_07141_));
 MUX2_X1 _12683_ (.A(_06594_),
    .B(_07141_),
    .S(_06666_),
    .Z(_07142_));
 NAND2_X1 _12684_ (.A1(_07138_),
    .A2(_07142_),
    .ZN(_07143_));
 INV_X1 _12685_ (.A(_05858_),
    .ZN(_07144_));
 NOR4_X2 _12686_ (.A1(_07144_),
    .A2(\dynamic_node_top.proc_input.control.count_f[0] ),
    .A3(\dynamic_node_top.proc_input.control.count_f[1] ),
    .A4(\dynamic_node_top.proc_input.control.count_f[2] ),
    .ZN(_07145_));
 NOR2_X1 _12687_ (.A1(\dynamic_node_top.proc_input.control.count_f[3] ),
    .A2(\dynamic_node_top.proc_input.control.count_f[4] ),
    .ZN(_07146_));
 NAND2_X1 _12688_ (.A1(_07145_),
    .A2(_07146_),
    .ZN(_07147_));
 XNOR2_X1 _12689_ (.A(\dynamic_node_top.proc_input.control.count_f[5] ),
    .B(_07147_),
    .ZN(_07148_));
 MUX2_X1 _12690_ (.A(_05972_),
    .B(_07148_),
    .S(_06666_),
    .Z(_07149_));
 XOR2_X1 _12691_ (.A(\dynamic_node_top.proc_input.control.count_f[3] ),
    .B(_07145_),
    .Z(_07150_));
 MUX2_X1 _12692_ (.A(_05902_),
    .B(_07150_),
    .S(_06666_),
    .Z(_07151_));
 NOR3_X1 _12693_ (.A1(_07143_),
    .A2(_07149_),
    .A3(_07151_),
    .ZN(_07152_));
 NOR2_X1 _12694_ (.A1(_05858_),
    .A2(\dynamic_node_top.proc_input.control.count_f[1] ),
    .ZN(_07153_));
 AOI221_X2 _12695_ (.A(_07153_),
    .B1(_05182_),
    .B2(\dynamic_node_top.proc_input.control.header_last_temp ),
    .C1(_05858_),
    .C2(_10534_),
    .ZN(_07154_));
 NOR2_X1 _12696_ (.A1(_06009_),
    .A2(_06018_),
    .ZN(_07155_));
 AOI21_X4 _12697_ (.A(_07155_),
    .B1(_06038_),
    .B2(_07130_),
    .ZN(_07156_));
 AOI21_X1 _12698_ (.A(_07154_),
    .B1(_07156_),
    .B2(_06183_),
    .ZN(_07157_));
 XNOR2_X1 _12699_ (.A(\dynamic_node_top.proc_input.control.count_f[4] ),
    .B(_07139_),
    .ZN(_07158_));
 OAI21_X1 _12700_ (.A(_05933_),
    .B1(_07158_),
    .B2(_06183_),
    .ZN(_07159_));
 NOR3_X1 _12701_ (.A1(\dynamic_node_top.proc_input.control.count_f[5] ),
    .A2(\dynamic_node_top.proc_input.control.count_f[6] ),
    .A3(_07147_),
    .ZN(_07160_));
 XNOR2_X1 _12702_ (.A(\dynamic_node_top.proc_input.control.count_f[7] ),
    .B(_07160_),
    .ZN(_07161_));
 NOR2_X1 _12703_ (.A1(_06183_),
    .A2(_07161_),
    .ZN(_07162_));
 AOI21_X1 _12704_ (.A(_07162_),
    .B1(_06183_),
    .B2(_05993_),
    .ZN(_07163_));
 NAND4_X1 _12705_ (.A1(_07152_),
    .A2(_07157_),
    .A3(_07159_),
    .A4(_07163_),
    .ZN(_07164_));
 OAI21_X1 _12706_ (.A(_06880_),
    .B1(_07134_),
    .B2(_07164_),
    .ZN(_07165_));
 OR2_X1 _12707_ (.A1(\dynamic_node_top.proc_input.control.header_last_temp ),
    .A2(_06541_),
    .ZN(_07166_));
 MUX2_X1 _12708_ (.A(_07165_),
    .B(_07166_),
    .S(_10456_),
    .Z(_00002_));
 OR3_X1 _12709_ (.A1(_05167_),
    .A2(_05158_),
    .A3(_07077_),
    .ZN(_07167_));
 NOR2_X2 _12710_ (.A1(_05308_),
    .A2(_07167_),
    .ZN(_07168_));
 AOI222_X2 _12711_ (.A1(_05340_),
    .A2(net624),
    .B1(_05597_),
    .B2(net623),
    .C1(_05824_),
    .C2(net622),
    .ZN(_07169_));
 INV_X2 _12712_ (.A(_07169_),
    .ZN(_07170_));
 NOR2_X1 _12713_ (.A1(_05478_),
    .A2(_07085_),
    .ZN(_07171_));
 NOR3_X4 _12714_ (.A1(_07168_),
    .A2(_07170_),
    .A3(_07171_),
    .ZN(_10464_));
 INV_X2 _12715_ (.A(_10464_),
    .ZN(\dynamic_node_top.south_input.NIB.thanks_in ));
 XOR2_X1 _12716_ (.A(_06052_),
    .B(\dynamic_node_top.south_input.control.count_f[0] ),
    .Z(_07172_));
 MUX2_X1 _12717_ (.A(_06080_),
    .B(_07172_),
    .S(_06096_),
    .Z(_07173_));
 NOR2_X1 _12718_ (.A1(_06057_),
    .A2(_06068_),
    .ZN(_07174_));
 BUF_X1 _12719_ (.A(\dynamic_node_top.south_input.control.count_f[2] ),
    .Z(_07175_));
 NAND2_X1 _12720_ (.A1(_06052_),
    .A2(_10515_),
    .ZN(_07176_));
 OR3_X1 _12721_ (.A1(_07175_),
    .A2(\dynamic_node_top.south_input.control.count_f[3] ),
    .A3(_07176_),
    .ZN(_07177_));
 XNOR2_X1 _12722_ (.A(\dynamic_node_top.south_input.control.count_f[4] ),
    .B(_07177_),
    .ZN(_07178_));
 NOR2_X1 _12723_ (.A1(_06103_),
    .A2(_07178_),
    .ZN(_07179_));
 INV_X1 _12724_ (.A(_06052_),
    .ZN(_07180_));
 OR4_X1 _12725_ (.A1(_07180_),
    .A2(\dynamic_node_top.south_input.control.count_f[0] ),
    .A3(\dynamic_node_top.south_input.control.count_f[1] ),
    .A4(_07175_),
    .ZN(_07181_));
 XNOR2_X1 _12726_ (.A(\dynamic_node_top.south_input.control.count_f[3] ),
    .B(_07181_),
    .ZN(_07182_));
 OR3_X1 _12727_ (.A1(_06052_),
    .A2(\dynamic_node_top.south_input.control.count_f[1] ),
    .A3(_07175_),
    .ZN(_07183_));
 XNOR2_X1 _12728_ (.A(_10515_),
    .B(_07175_),
    .ZN(_07184_));
 NAND3_X1 _12729_ (.A1(_06052_),
    .A2(_10516_),
    .A3(_07184_),
    .ZN(_07185_));
 AOI21_X1 _12730_ (.A(_07182_),
    .B1(_07183_),
    .B2(_07185_),
    .ZN(_07186_));
 AOI21_X1 _12731_ (.A(_07174_),
    .B1(_07179_),
    .B2(_07186_),
    .ZN(_07187_));
 OR3_X1 _12732_ (.A1(\dynamic_node_top.south_input.control.count_f[3] ),
    .A2(\dynamic_node_top.south_input.control.count_f[4] ),
    .A3(_07181_),
    .ZN(_07188_));
 NOR3_X1 _12733_ (.A1(\dynamic_node_top.south_input.control.count_f[5] ),
    .A2(\dynamic_node_top.south_input.control.count_f[6] ),
    .A3(_07188_),
    .ZN(_07189_));
 XOR2_X1 _12734_ (.A(\dynamic_node_top.south_input.control.count_f[7] ),
    .B(_07189_),
    .Z(_07190_));
 MUX2_X1 _12735_ (.A(_06071_),
    .B(_07190_),
    .S(_06096_),
    .Z(_07191_));
 INV_X2 _12736_ (.A(_06077_),
    .ZN(_07192_));
 NOR3_X1 _12737_ (.A1(\dynamic_node_top.south_input.control.count_f[4] ),
    .A2(\dynamic_node_top.south_input.control.count_f[5] ),
    .A3(_07177_),
    .ZN(_07193_));
 XNOR2_X1 _12738_ (.A(\dynamic_node_top.south_input.control.count_f[6] ),
    .B(_07193_),
    .ZN(_07194_));
 MUX2_X1 _12739_ (.A(_07192_),
    .B(_07194_),
    .S(_06096_),
    .Z(_07195_));
 INV_X2 _12740_ (.A(_06074_),
    .ZN(_07196_));
 XOR2_X1 _12741_ (.A(\dynamic_node_top.south_input.control.count_f[5] ),
    .B(_07188_),
    .Z(_07197_));
 MUX2_X1 _12742_ (.A(_07196_),
    .B(_07197_),
    .S(_06096_),
    .Z(_07198_));
 NAND2_X1 _12743_ (.A1(_07195_),
    .A2(_07198_),
    .ZN(_07199_));
 NOR4_X1 _12744_ (.A1(_07173_),
    .A2(_07187_),
    .A3(_07191_),
    .A4(_07199_),
    .ZN(_07200_));
 MUX2_X1 _12745_ (.A(\dynamic_node_top.south_input.control.header_last_temp ),
    .B(_07200_),
    .S(\dynamic_node_top.south_input.NIB.thanks_in ),
    .Z(_07201_));
 OR2_X1 _12746_ (.A1(_06573_),
    .A2(_07201_),
    .ZN(_00003_));
 OAI211_X2 _12747_ (.A(_05178_),
    .B(_05184_),
    .C1(_05306_),
    .C2(_05307_),
    .ZN(_07202_));
 NOR2_X1 _12748_ (.A1(_05329_),
    .A2(_05330_),
    .ZN(_07203_));
 NAND3_X1 _12749_ (.A1(_07203_),
    .A2(net624),
    .A3(_07043_),
    .ZN(_07204_));
 NAND4_X1 _12750_ (.A1(_07022_),
    .A2(_05857_),
    .A3(_06520_),
    .A4(_07028_),
    .ZN(_07205_));
 AOI211_X2 _12751_ (.A(_06095_),
    .B(_07205_),
    .C1(_06120_),
    .C2(_06122_),
    .ZN(_07206_));
 NOR4_X2 _12752_ (.A1(_05594_),
    .A2(_05595_),
    .A3(_05603_),
    .A4(_05596_),
    .ZN(_07207_));
 AOI221_X2 _12753_ (.A(_07206_),
    .B1(_07207_),
    .B2(net623),
    .C1(_05472_),
    .C2(net757),
    .ZN(_07208_));
 AND3_X2 _12754_ (.A1(_07202_),
    .A2(_07204_),
    .A3(_07208_),
    .ZN(_10506_));
 INV_X1 _12755_ (.A(_10506_),
    .ZN(\dynamic_node_top.east_input.NIB.thanks_in ));
 NOR2_X1 _12756_ (.A1(_05488_),
    .A2(\dynamic_node_top.east_input.NIB.thanks_in ),
    .ZN(_07209_));
 XOR2_X1 _12757_ (.A(_05787_),
    .B(\dynamic_node_top.east_input.control.count_f[0] ),
    .Z(_07210_));
 MUX2_X1 _12758_ (.A(_05775_),
    .B(_07210_),
    .S(_06793_),
    .Z(_07211_));
 BUF_X1 _12759_ (.A(\dynamic_node_top.east_input.control.count_f[2] ),
    .Z(_07212_));
 NAND2_X1 _12760_ (.A1(_05787_),
    .A2(_10440_),
    .ZN(_07213_));
 OR3_X1 _12761_ (.A1(_07212_),
    .A2(\dynamic_node_top.east_input.control.count_f[3] ),
    .A3(_07213_),
    .ZN(_07214_));
 XNOR2_X1 _12762_ (.A(\dynamic_node_top.east_input.control.count_f[4] ),
    .B(_07214_),
    .ZN(_07215_));
 NOR2_X1 _12763_ (.A1(_06787_),
    .A2(_07215_),
    .ZN(_07216_));
 INV_X1 _12764_ (.A(_05787_),
    .ZN(_07217_));
 OR4_X1 _12765_ (.A1(_07217_),
    .A2(\dynamic_node_top.east_input.control.count_f[0] ),
    .A3(\dynamic_node_top.east_input.control.count_f[1] ),
    .A4(_07212_),
    .ZN(_07218_));
 XNOR2_X1 _12766_ (.A(\dynamic_node_top.east_input.control.count_f[3] ),
    .B(_07218_),
    .ZN(_07219_));
 OR3_X1 _12767_ (.A1(_05787_),
    .A2(\dynamic_node_top.east_input.control.count_f[1] ),
    .A3(_07212_),
    .ZN(_07220_));
 XNOR2_X1 _12768_ (.A(_10440_),
    .B(_07212_),
    .ZN(_07221_));
 NAND3_X1 _12769_ (.A1(_05787_),
    .A2(_10441_),
    .A3(_07221_),
    .ZN(_07222_));
 AOI21_X1 _12770_ (.A(_07219_),
    .B1(_07220_),
    .B2(_07222_),
    .ZN(_07223_));
 AOI22_X2 _12771_ (.A1(_05761_),
    .A2(_05772_),
    .B1(_07216_),
    .B2(_07223_),
    .ZN(_07224_));
 OR3_X1 _12772_ (.A1(\dynamic_node_top.east_input.control.count_f[3] ),
    .A2(\dynamic_node_top.east_input.control.count_f[4] ),
    .A3(_07218_),
    .ZN(_07225_));
 NOR3_X1 _12773_ (.A1(\dynamic_node_top.east_input.control.count_f[5] ),
    .A2(\dynamic_node_top.east_input.control.count_f[6] ),
    .A3(_07225_),
    .ZN(_07226_));
 XOR2_X1 _12774_ (.A(\dynamic_node_top.east_input.control.count_f[7] ),
    .B(_07226_),
    .Z(_07227_));
 MUX2_X1 _12775_ (.A(_05778_),
    .B(_07227_),
    .S(_06793_),
    .Z(_07228_));
 INV_X2 _12776_ (.A(_05784_),
    .ZN(_07229_));
 NOR3_X1 _12777_ (.A1(\dynamic_node_top.east_input.control.count_f[4] ),
    .A2(\dynamic_node_top.east_input.control.count_f[5] ),
    .A3(_07214_),
    .ZN(_07230_));
 XNOR2_X1 _12778_ (.A(\dynamic_node_top.east_input.control.count_f[6] ),
    .B(_07230_),
    .ZN(_07231_));
 MUX2_X1 _12779_ (.A(_07229_),
    .B(_07231_),
    .S(_06793_),
    .Z(_07232_));
 INV_X2 _12780_ (.A(_05781_),
    .ZN(_07233_));
 XOR2_X1 _12781_ (.A(\dynamic_node_top.east_input.control.count_f[5] ),
    .B(_07225_),
    .Z(_07234_));
 MUX2_X1 _12782_ (.A(_07233_),
    .B(_07234_),
    .S(_06793_),
    .Z(_07235_));
 NAND2_X1 _12783_ (.A1(_07232_),
    .A2(_07235_),
    .ZN(_07236_));
 NOR4_X1 _12784_ (.A1(_07211_),
    .A2(_07224_),
    .A3(_07228_),
    .A4(_07236_),
    .ZN(_07237_));
 NOR2_X1 _12785_ (.A1(_10506_),
    .A2(_07237_),
    .ZN(_07238_));
 OAI21_X1 _12786_ (.A(_06892_),
    .B1(_07209_),
    .B2(_07238_),
    .ZN(_00000_));
 MUX2_X1 _12787_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][45] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][45] ),
    .S(net765),
    .Z(_07239_));
 INV_X1 _12788_ (.A(_07239_),
    .ZN(_07240_));
 NAND2_X1 _12789_ (.A1(_05126_),
    .A2(_07240_),
    .ZN(_07241_));
 BUF_X8 _12790_ (.A(_05130_),
    .Z(_07242_));
 MUX2_X1 _12791_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][45] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][45] ),
    .S(_07242_),
    .Z(_07243_));
 OAI21_X4 _12792_ (.A(_07241_),
    .B1(_07243_),
    .B2(_05127_),
    .ZN(_10185_));
 BUF_X8 _12793_ (.A(_05126_),
    .Z(_07244_));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 BUF_X16 _12795_ (.A(_05132_),
    .Z(_07246_));
 MUX2_X1 _12796_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][49] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][49] ),
    .S(_07246_),
    .Z(_07247_));
 INV_X1 _12797_ (.A(_07247_),
    .ZN(_07248_));
 NAND2_X1 _12798_ (.A1(_07244_),
    .A2(_07248_),
    .ZN(_07249_));
 BUF_X16 _12799_ (.A(_05136_),
    .Z(_07250_));
 MUX2_X1 _12800_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][49] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][49] ),
    .S(_07250_),
    .Z(_07251_));
 OAI21_X4 _12801_ (.A(_07249_),
    .B1(_07251_),
    .B2(_07244_),
    .ZN(_10191_));
 MUX2_X1 _12802_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][47] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][47] ),
    .S(_05130_),
    .Z(_07252_));
 INV_X1 _12803_ (.A(_07252_),
    .ZN(_07253_));
 NAND2_X1 _12804_ (.A1(_05126_),
    .A2(_07253_),
    .ZN(_07254_));
 MUX2_X1 _12805_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][47] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][47] ),
    .S(_07242_),
    .Z(_07255_));
 BUF_X4 _12806_ (.A(_05126_),
    .Z(_07256_));
 OAI21_X4 _12807_ (.A(_07254_),
    .B1(_07255_),
    .B2(_07256_),
    .ZN(_10197_));
 MUX2_X1 _12808_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][46] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][46] ),
    .S(_05132_),
    .Z(_07257_));
 INV_X1 _12809_ (.A(_07257_),
    .ZN(_07258_));
 NAND2_X1 _12810_ (.A1(_07256_),
    .A2(_07258_),
    .ZN(_07259_));
 MUX2_X1 _12811_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][46] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][46] ),
    .S(_07242_),
    .Z(_07260_));
 OAI21_X4 _12812_ (.A(_07259_),
    .B1(_05127_),
    .B2(_07260_),
    .ZN(_10200_));
 MUX2_X1 _12813_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][41] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][41] ),
    .S(_07246_),
    .Z(_07261_));
 INV_X2 _12814_ (.A(_07261_),
    .ZN(_07262_));
 NAND2_X2 _12815_ (.A1(_07244_),
    .A2(_07262_),
    .ZN(_07263_));
 MUX2_X1 _12816_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][41] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][41] ),
    .S(_07250_),
    .Z(_07264_));
 OAI21_X4 _12817_ (.A(_07263_),
    .B1(_07244_),
    .B2(_07264_),
    .ZN(_10203_));
 MUX2_X1 _12818_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][37] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][37] ),
    .S(_05136_),
    .Z(_07265_));
 MUX2_X1 _12819_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][37] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][37] ),
    .S(_05136_),
    .Z(_07266_));
 MUX2_X2 _12820_ (.A(_07265_),
    .B(_07266_),
    .S(_07256_),
    .Z(_07267_));
 INV_X4 _12821_ (.A(_07267_),
    .ZN(_10215_));
 CLKBUF_X3 _12822_ (.A(_05152_),
    .Z(_07268_));
 MUX2_X1 _12823_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][45] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][45] ),
    .S(net737),
    .Z(_07269_));
 OR2_X1 _12824_ (.A1(_07268_),
    .A2(_07269_),
    .ZN(_07270_));
 MUX2_X1 _12825_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][45] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][45] ),
    .S(_05147_),
    .Z(_07271_));
 BUF_X8 _12826_ (.A(_05201_),
    .Z(_07272_));
 OAI21_X4 _12827_ (.A(_07270_),
    .B1(_07271_),
    .B2(_07272_),
    .ZN(_10240_));
 BUF_X32 _12828_ (.A(_05144_),
    .Z(_07273_));
 MUX2_X1 _12829_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][37] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][37] ),
    .S(_07273_),
    .Z(_07274_));
 OR2_X1 _12830_ (.A1(_07268_),
    .A2(_07274_),
    .ZN(_07275_));
 MUX2_X1 _12831_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][37] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][37] ),
    .S(_05147_),
    .Z(_07276_));
 OAI21_X4 _12832_ (.A(_07275_),
    .B1(_07276_),
    .B2(_07272_),
    .ZN(_10258_));
 MUX2_X1 _12833_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][39] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][39] ),
    .S(_05146_),
    .Z(_07277_));
 MUX2_X1 _12834_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][39] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][39] ),
    .S(_05146_),
    .Z(_07278_));
 MUX2_X2 _12835_ (.A(_07277_),
    .B(_07278_),
    .S(_05152_),
    .Z(_07279_));
 INV_X4 _12836_ (.A(_07279_),
    .ZN(_10270_));
 MUX2_X1 _12837_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][38] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][38] ),
    .S(_05144_),
    .Z(_07280_));
 MUX2_X1 _12838_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][38] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][38] ),
    .S(_05144_),
    .Z(_07281_));
 MUX2_X2 _12839_ (.A(_07280_),
    .B(_07281_),
    .S(_05152_),
    .Z(_07282_));
 INV_X2 _12840_ (.A(_07282_),
    .ZN(_10273_));
 MUX2_X1 _12841_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][37] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][37] ),
    .S(_05314_),
    .Z(_07283_));
 OR2_X2 _12842_ (.A1(_05321_),
    .A2(_07283_),
    .ZN(_07284_));
 MUX2_X1 _12843_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][37] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][37] ),
    .S(_05315_),
    .Z(_07285_));
 OAI21_X4 _12844_ (.A(_07284_),
    .B1(_07285_),
    .B2(_05326_),
    .ZN(_10312_));
 BUF_X16 _12845_ (.A(_05456_),
    .Z(_07286_));
 MUX2_X1 _12846_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][47] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][47] ),
    .S(_07286_),
    .Z(_07287_));
 OR2_X1 _12847_ (.A1(_05468_),
    .A2(_07287_),
    .ZN(_07288_));
 MUX2_X1 _12848_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][47] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][47] ),
    .S(net721),
    .Z(_07289_));
 BUF_X8 _12849_ (.A(_05495_),
    .Z(_07290_));
 OAI21_X4 _12850_ (.A(_07288_),
    .B1(_07289_),
    .B2(_07290_),
    .ZN(_10330_));
 MUX2_X1 _12851_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][46] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][46] ),
    .S(_05459_),
    .Z(_07291_));
 MUX2_X1 _12852_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][46] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][46] ),
    .S(_05459_),
    .Z(_07292_));
 MUX2_X2 _12853_ (.A(_07291_),
    .B(_07292_),
    .S(_05465_),
    .Z(_07293_));
 INV_X4 _12854_ (.A(_07293_),
    .ZN(_10333_));
 MUX2_X1 _12855_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][45] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][45] ),
    .S(net717),
    .Z(_07294_));
 MUX2_X1 _12856_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][45] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][45] ),
    .S(_05456_),
    .Z(_07295_));
 MUX2_X2 _12857_ (.A(_07294_),
    .B(_07295_),
    .S(_05463_),
    .Z(_07296_));
 INV_X2 _12858_ (.A(_07296_),
    .ZN(_10336_));
 MUX2_X1 _12859_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][43] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][43] ),
    .S(_05458_),
    .Z(_07297_));
 OR2_X1 _12860_ (.A1(_05468_),
    .A2(_07297_),
    .ZN(_07298_));
 MUX2_X1 _12861_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][43] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][43] ),
    .S(_07286_),
    .Z(_07299_));
 OAI21_X4 _12862_ (.A(_07298_),
    .B1(_07299_),
    .B2(_07290_),
    .ZN(_10342_));
 MUX2_X1 _12863_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][35] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][35] ),
    .S(net720),
    .Z(_07300_));
 MUX2_X1 _12864_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][35] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][35] ),
    .S(net720),
    .Z(_07301_));
 MUX2_X2 _12865_ (.A(_07300_),
    .B(_07301_),
    .S(_05463_),
    .Z(_07302_));
 INV_X4 _12866_ (.A(_07302_),
    .ZN(_10351_));
 MUX2_X1 _12867_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][37] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][37] ),
    .S(_05456_),
    .Z(_07303_));
 MUX2_X1 _12868_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][37] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][37] ),
    .S(_05456_),
    .Z(_07304_));
 MUX2_X2 _12869_ (.A(_07303_),
    .B(_07304_),
    .S(_05463_),
    .Z(_07305_));
 INV_X1 _12870_ (.A(_07305_),
    .ZN(_10354_));
 MUX2_X1 _12871_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][39] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][39] ),
    .S(net720),
    .Z(_07306_));
 OR2_X1 _12872_ (.A1(_05468_),
    .A2(_07306_),
    .ZN(_07307_));
 MUX2_X1 _12873_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][39] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][39] ),
    .S(_07286_),
    .Z(_07308_));
 OAI21_X4 _12874_ (.A(_07307_),
    .B1(_07308_),
    .B2(_07290_),
    .ZN(_10366_));
 MUX2_X1 _12875_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][38] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][38] ),
    .S(net720),
    .Z(_07309_));
 OR2_X1 _12876_ (.A1(_05468_),
    .A2(_07309_),
    .ZN(_07310_));
 MUX2_X1 _12877_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][38] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][38] ),
    .S(_07286_),
    .Z(_07311_));
 OAI21_X4 _12878_ (.A(_07310_),
    .B1(_07311_),
    .B2(_07290_),
    .ZN(_10369_));
 BUF_X4 _12879_ (.A(_05703_),
    .Z(_07312_));
 MUX2_X1 _12880_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][45] ),
    .S(_07312_),
    .Z(_07313_));
 BUF_X4 _12881_ (.A(_05703_),
    .Z(_07314_));
 MUX2_X1 _12882_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][45] ),
    .S(_07314_),
    .Z(_07315_));
 BUF_X4 _12883_ (.A(_05710_),
    .Z(_07316_));
 MUX2_X1 _12884_ (.A(_07313_),
    .B(_07315_),
    .S(_07316_),
    .Z(_07317_));
 MUX2_X1 _12885_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][45] ),
    .S(_07314_),
    .Z(_07318_));
 BUF_X4 _12886_ (.A(_05703_),
    .Z(_07319_));
 MUX2_X1 _12887_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][45] ),
    .S(_07319_),
    .Z(_07320_));
 BUF_X4 _12888_ (.A(_05710_),
    .Z(_07321_));
 MUX2_X1 _12889_ (.A(_07318_),
    .B(_07320_),
    .S(_07321_),
    .Z(_07322_));
 BUF_X4 _12890_ (.A(_05720_),
    .Z(_07323_));
 MUX2_X1 _12891_ (.A(_07317_),
    .B(_07322_),
    .S(_07323_),
    .Z(_07324_));
 BUF_X4 _12892_ (.A(_05702_),
    .Z(_07325_));
 BUF_X4 _12893_ (.A(_07325_),
    .Z(_07326_));
 MUX2_X1 _12894_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][45] ),
    .S(_07326_),
    .Z(_07327_));
 BUF_X4 _12895_ (.A(_07325_),
    .Z(_07328_));
 MUX2_X1 _12896_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][45] ),
    .S(_07328_),
    .Z(_07329_));
 BUF_X4 _12897_ (.A(_05710_),
    .Z(_07330_));
 MUX2_X1 _12898_ (.A(_07327_),
    .B(_07329_),
    .S(_07330_),
    .Z(_07331_));
 BUF_X4 _12899_ (.A(_07325_),
    .Z(_07332_));
 MUX2_X1 _12900_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][45] ),
    .S(_07332_),
    .Z(_07333_));
 BUF_X4 _12901_ (.A(_07325_),
    .Z(_07334_));
 MUX2_X1 _12902_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][45] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][45] ),
    .S(_07334_),
    .Z(_07335_));
 BUF_X4 _12903_ (.A(_05709_),
    .Z(_07336_));
 BUF_X4 _12904_ (.A(_07336_),
    .Z(_07337_));
 MUX2_X1 _12905_ (.A(_07333_),
    .B(_07335_),
    .S(_07337_),
    .Z(_07338_));
 BUF_X4 _12906_ (.A(_05720_),
    .Z(_07339_));
 MUX2_X1 _12907_ (.A(_07331_),
    .B(_07338_),
    .S(_07339_),
    .Z(_07340_));
 BUF_X4 _12908_ (.A(_05738_),
    .Z(_07341_));
 MUX2_X2 _12909_ (.A(_07324_),
    .B(_07340_),
    .S(_07341_),
    .Z(_07342_));
 INV_X1 _12910_ (.A(_07342_),
    .ZN(_10378_));
 MUX2_X1 _12911_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][47] ),
    .S(_07312_),
    .Z(_07343_));
 BUF_X4 _12912_ (.A(_05703_),
    .Z(_07344_));
 MUX2_X1 _12913_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][47] ),
    .S(_07344_),
    .Z(_07345_));
 MUX2_X1 _12914_ (.A(_07343_),
    .B(_07345_),
    .S(_05729_),
    .Z(_07346_));
 MUX2_X1 _12915_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][47] ),
    .S(_07344_),
    .Z(_07347_));
 BUF_X4 _12916_ (.A(_05703_),
    .Z(_07348_));
 MUX2_X1 _12917_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][47] ),
    .S(_07348_),
    .Z(_07349_));
 MUX2_X1 _12918_ (.A(_07347_),
    .B(_07349_),
    .S(_07316_),
    .Z(_07350_));
 MUX2_X1 _12919_ (.A(_07346_),
    .B(_07350_),
    .S(_05721_),
    .Z(_07351_));
 BUF_X4 _12920_ (.A(_07325_),
    .Z(_07352_));
 MUX2_X1 _12921_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][47] ),
    .S(_07352_),
    .Z(_07353_));
 MUX2_X1 _12922_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][47] ),
    .S(_07326_),
    .Z(_07354_));
 MUX2_X1 _12923_ (.A(_07353_),
    .B(_07354_),
    .S(_07330_),
    .Z(_07355_));
 MUX2_X1 _12924_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][47] ),
    .S(_07328_),
    .Z(_07356_));
 MUX2_X1 _12925_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][47] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][47] ),
    .S(_07334_),
    .Z(_07357_));
 BUF_X4 _12926_ (.A(_07336_),
    .Z(_07358_));
 MUX2_X1 _12927_ (.A(_07356_),
    .B(_07357_),
    .S(_07358_),
    .Z(_07359_));
 MUX2_X1 _12928_ (.A(_07355_),
    .B(_07359_),
    .S(_07339_),
    .Z(_07360_));
 MUX2_X2 _12929_ (.A(_07351_),
    .B(_07360_),
    .S(_07341_),
    .Z(_07361_));
 INV_X1 _12930_ (.A(_07361_),
    .ZN(_10390_));
 MUX2_X1 _12931_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][46] ),
    .S(_05724_),
    .Z(_07362_));
 MUX2_X1 _12932_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][46] ),
    .S(_07344_),
    .Z(_07363_));
 MUX2_X1 _12933_ (.A(_07362_),
    .B(_07363_),
    .S(_05729_),
    .Z(_07364_));
 MUX2_X1 _12934_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][46] ),
    .S(_07344_),
    .Z(_07365_));
 MUX2_X1 _12935_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][46] ),
    .S(_07348_),
    .Z(_07366_));
 MUX2_X1 _12936_ (.A(_07365_),
    .B(_07366_),
    .S(_07316_),
    .Z(_07367_));
 MUX2_X1 _12937_ (.A(_07364_),
    .B(_07367_),
    .S(_05721_),
    .Z(_07368_));
 MUX2_X1 _12938_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][46] ),
    .S(_07352_),
    .Z(_07369_));
 MUX2_X1 _12939_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][46] ),
    .S(_07326_),
    .Z(_07370_));
 MUX2_X1 _12940_ (.A(_07369_),
    .B(_07370_),
    .S(_07330_),
    .Z(_07371_));
 MUX2_X1 _12941_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][46] ),
    .S(_07328_),
    .Z(_07372_));
 MUX2_X1 _12942_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][46] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][46] ),
    .S(_07334_),
    .Z(_07373_));
 MUX2_X1 _12943_ (.A(_07372_),
    .B(_07373_),
    .S(_07358_),
    .Z(_07374_));
 MUX2_X1 _12944_ (.A(_07371_),
    .B(_07374_),
    .S(_07339_),
    .Z(_07375_));
 MUX2_X2 _12945_ (.A(_07368_),
    .B(_07375_),
    .S(_07341_),
    .Z(_07376_));
 INV_X1 _12946_ (.A(_07376_),
    .ZN(_10393_));
 MUX2_X1 _12947_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][41] ),
    .S(_07319_),
    .Z(_07377_));
 MUX2_X1 _12948_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][41] ),
    .S(_07319_),
    .Z(_07378_));
 MUX2_X1 _12949_ (.A(_07377_),
    .B(_07378_),
    .S(_07321_),
    .Z(_07379_));
 MUX2_X1 _12950_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][41] ),
    .S(_07319_),
    .Z(_07380_));
 MUX2_X1 _12951_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][41] ),
    .S(_07352_),
    .Z(_07381_));
 MUX2_X1 _12952_ (.A(_07380_),
    .B(_07381_),
    .S(_07321_),
    .Z(_07382_));
 MUX2_X1 _12953_ (.A(_07379_),
    .B(_07382_),
    .S(_07323_),
    .Z(_07383_));
 BUF_X4 _12954_ (.A(_07325_),
    .Z(_07384_));
 MUX2_X1 _12955_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][41] ),
    .S(_07384_),
    .Z(_07385_));
 MUX2_X1 _12956_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][41] ),
    .S(_07384_),
    .Z(_07386_));
 MUX2_X1 _12957_ (.A(_07385_),
    .B(_07386_),
    .S(_07337_),
    .Z(_07387_));
 MUX2_X1 _12958_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][41] ),
    .S(_07384_),
    .Z(_07388_));
 MUX2_X1 _12959_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][41] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][41] ),
    .S(_07384_),
    .Z(_07389_));
 MUX2_X1 _12960_ (.A(_07388_),
    .B(_07389_),
    .S(_07337_),
    .Z(_07390_));
 BUF_X4 _12961_ (.A(_05720_),
    .Z(_07391_));
 MUX2_X1 _12962_ (.A(_07387_),
    .B(_07390_),
    .S(_07391_),
    .Z(_07392_));
 BUF_X4 _12963_ (.A(_05737_),
    .Z(_07393_));
 MUX2_X2 _12964_ (.A(_07383_),
    .B(_07392_),
    .S(_07393_),
    .Z(_07394_));
 INV_X1 _12965_ (.A(_07394_),
    .ZN(_10396_));
 MUX2_X1 _12966_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][37] ),
    .S(_07312_),
    .Z(_07395_));
 MUX2_X1 _12967_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][37] ),
    .S(_07314_),
    .Z(_07396_));
 MUX2_X1 _12968_ (.A(_07395_),
    .B(_07396_),
    .S(_07316_),
    .Z(_07397_));
 MUX2_X1 _12969_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][37] ),
    .S(_07348_),
    .Z(_07398_));
 MUX2_X1 _12970_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][37] ),
    .S(_07319_),
    .Z(_07399_));
 MUX2_X1 _12971_ (.A(_07398_),
    .B(_07399_),
    .S(_07321_),
    .Z(_07400_));
 MUX2_X1 _12972_ (.A(_07397_),
    .B(_07400_),
    .S(_07323_),
    .Z(_07401_));
 MUX2_X1 _12973_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][37] ),
    .S(_07326_),
    .Z(_07402_));
 MUX2_X1 _12974_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][37] ),
    .S(_07332_),
    .Z(_07403_));
 MUX2_X1 _12975_ (.A(_07402_),
    .B(_07403_),
    .S(_07358_),
    .Z(_07404_));
 MUX2_X1 _12976_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][37] ),
    .S(_07332_),
    .Z(_07405_));
 MUX2_X1 _12977_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][37] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][37] ),
    .S(_07334_),
    .Z(_07406_));
 MUX2_X1 _12978_ (.A(_07405_),
    .B(_07406_),
    .S(_07337_),
    .Z(_07407_));
 MUX2_X1 _12979_ (.A(_07404_),
    .B(_07407_),
    .S(_07391_),
    .Z(_07408_));
 MUX2_X2 _12980_ (.A(_07401_),
    .B(_07408_),
    .S(_07393_),
    .Z(_07409_));
 INV_X1 _12981_ (.A(_07409_),
    .ZN(_10408_));
 INV_X2 _12982_ (.A(net293),
    .ZN(_10463_));
 INV_X2 _12983_ (.A(net291),
    .ZN(_10471_));
 INV_X2 _12984_ (.A(net294),
    .ZN(_10497_));
 INV_X2 _12985_ (.A(net290),
    .ZN(_10505_));
 MUX2_X1 _12986_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][43] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][43] ),
    .S(_05132_),
    .Z(_07410_));
 INV_X2 _12987_ (.A(_07410_),
    .ZN(_07411_));
 NAND2_X4 _12988_ (.A1(_07256_),
    .A2(_07411_),
    .ZN(_07412_));
 MUX2_X1 _12989_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][43] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][43] ),
    .S(_07242_),
    .Z(_07413_));
 OAI21_X4 _12990_ (.A(_07412_),
    .B1(_05127_),
    .B2(_07413_),
    .ZN(_10182_));
 MUX2_X1 _12991_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][44] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][44] ),
    .S(_05132_),
    .Z(_07414_));
 INV_X2 _12992_ (.A(_07414_),
    .ZN(_07415_));
 NAND2_X2 _12993_ (.A1(_07256_),
    .A2(_07415_),
    .ZN(_07416_));
 MUX2_X1 _12994_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][44] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][44] ),
    .S(_07242_),
    .Z(_07417_));
 OAI21_X4 _12995_ (.A(_07416_),
    .B1(_05127_),
    .B2(_07417_),
    .ZN(_10188_));
 MUX2_X1 _12996_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][48] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][48] ),
    .S(_07242_),
    .Z(_07418_));
 MUX2_X1 _12997_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][48] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][48] ),
    .S(_07242_),
    .Z(_07419_));
 MUX2_X2 _12998_ (.A(_07418_),
    .B(_07419_),
    .S(_05127_),
    .Z(_07420_));
 INV_X1 _12999_ (.A(_07420_),
    .ZN(_10194_));
 MUX2_X1 _13000_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][40] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][40] ),
    .S(net743),
    .Z(_07421_));
 INV_X1 _13001_ (.A(_07421_),
    .ZN(_07422_));
 NAND2_X1 _13002_ (.A1(_07256_),
    .A2(_07422_),
    .ZN(_07423_));
 MUX2_X1 _13003_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][40] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][40] ),
    .S(_07242_),
    .Z(_07424_));
 OAI21_X4 _13004_ (.A(_07423_),
    .B1(_07424_),
    .B2(_05127_),
    .ZN(_10206_));
 MUX2_X1 _13005_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][39] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][39] ),
    .S(net765),
    .Z(_07425_));
 INV_X1 _13006_ (.A(_07425_),
    .ZN(_07426_));
 NAND2_X1 _13007_ (.A1(_07256_),
    .A2(_07426_),
    .ZN(_07427_));
 MUX2_X1 _13008_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][39] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][39] ),
    .S(_07242_),
    .Z(_07428_));
 OAI21_X4 _13009_ (.A(_07427_),
    .B1(_07428_),
    .B2(_05127_),
    .ZN(_10209_));
 MUX2_X1 _13010_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][38] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][38] ),
    .S(_07242_),
    .Z(_07429_));
 MUX2_X1 _13011_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][38] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][38] ),
    .S(net745),
    .Z(_07430_));
 MUX2_X2 _13012_ (.A(_07429_),
    .B(_07430_),
    .S(_05126_),
    .Z(_07431_));
 INV_X1 _13013_ (.A(_07431_),
    .ZN(_10212_));
 MUX2_X1 _13014_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][36] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][36] ),
    .S(_05136_),
    .Z(_07432_));
 MUX2_X1 _13015_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][36] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][36] ),
    .S(_05136_),
    .Z(_07433_));
 MUX2_X2 _13016_ (.A(_07432_),
    .B(_07433_),
    .S(_07256_),
    .Z(_07434_));
 INV_X2 _13017_ (.A(_07434_),
    .ZN(_10218_));
 MUX2_X1 _13018_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][35] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][35] ),
    .S(net743),
    .Z(_07435_));
 INV_X1 _13019_ (.A(_07435_),
    .ZN(_07436_));
 NAND2_X1 _13020_ (.A1(_07256_),
    .A2(_07436_),
    .ZN(_07437_));
 MUX2_X1 _13021_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][35] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][35] ),
    .S(net743),
    .Z(_07438_));
 OAI21_X4 _13022_ (.A(_07437_),
    .B1(_07438_),
    .B2(_07256_),
    .ZN(_10221_));
 BUF_X4 _13023_ (.A(_05153_),
    .Z(_07439_));
 BUF_X16 _13024_ (.A(_07273_),
    .Z(_07440_));
 MUX2_X1 _13025_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][49] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][49] ),
    .S(_07440_),
    .Z(_07441_));
 OR2_X4 _13026_ (.A1(_07441_),
    .A2(_07439_),
    .ZN(_07442_));
 BUF_X16 _13027_ (.A(_05147_),
    .Z(_07443_));
 MUX2_X1 _13028_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][49] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][49] ),
    .S(_07443_),
    .Z(_07444_));
 BUF_X4 _13029_ (.A(_07272_),
    .Z(_07445_));
 BUF_X8 _13030_ (.A(_07445_),
    .Z(_07446_));
 OAI21_X4 _13031_ (.A(_07442_),
    .B1(_07444_),
    .B2(_07446_),
    .ZN(_10228_));
 MUX2_X1 _13032_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][48] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][48] ),
    .S(_07273_),
    .Z(_07447_));
 OR2_X1 _13033_ (.A1(_07268_),
    .A2(_07447_),
    .ZN(_07448_));
 MUX2_X1 _13034_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][48] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][48] ),
    .S(_05147_),
    .Z(_07449_));
 OAI21_X4 _13035_ (.A(_07448_),
    .B1(_07449_),
    .B2(_07272_),
    .ZN(_10231_));
 MUX2_X1 _13036_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][47] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][47] ),
    .S(_05146_),
    .Z(_07450_));
 OR2_X2 _13037_ (.A1(_07268_),
    .A2(_07450_),
    .ZN(_07451_));
 MUX2_X1 _13038_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][47] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][47] ),
    .S(_07273_),
    .Z(_07452_));
 OAI21_X4 _13039_ (.A(_07451_),
    .B1(_07452_),
    .B2(_07272_),
    .ZN(_10234_));
 MUX2_X1 _13040_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][46] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][46] ),
    .S(net737),
    .Z(_07453_));
 OR2_X1 _13041_ (.A1(_05152_),
    .A2(_07453_),
    .ZN(_07454_));
 MUX2_X1 _13042_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][46] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][46] ),
    .S(_07273_),
    .Z(_07455_));
 OAI21_X4 _13043_ (.A(_07454_),
    .B1(_07455_),
    .B2(_07272_),
    .ZN(_10237_));
 MUX2_X1 _13044_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][44] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][44] ),
    .S(net737),
    .Z(_07456_));
 OR2_X1 _13045_ (.A1(_07268_),
    .A2(_07456_),
    .ZN(_07457_));
 MUX2_X1 _13046_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][44] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][44] ),
    .S(_07273_),
    .Z(_07458_));
 OAI21_X4 _13047_ (.A(_07457_),
    .B1(_07458_),
    .B2(_07272_),
    .ZN(_10243_));
 MUX2_X1 _13048_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][43] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][43] ),
    .S(_05146_),
    .Z(_07459_));
 OR2_X2 _13049_ (.A1(_07268_),
    .A2(_07459_),
    .ZN(_07460_));
 MUX2_X1 _13050_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][43] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][43] ),
    .S(_07273_),
    .Z(_07461_));
 OAI21_X4 _13051_ (.A(_07460_),
    .B1(_07461_),
    .B2(_07272_),
    .ZN(_10246_));
 MUX2_X1 _13052_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][35] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][35] ),
    .S(net737),
    .Z(_07462_));
 OR2_X1 _13053_ (.A1(_07268_),
    .A2(_07462_),
    .ZN(_07463_));
 MUX2_X1 _13054_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][35] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][35] ),
    .S(_07273_),
    .Z(_07464_));
 OAI21_X4 _13055_ (.A(_07463_),
    .B1(_07464_),
    .B2(_07272_),
    .ZN(_10255_));
 MUX2_X1 _13056_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][36] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][36] ),
    .S(net737),
    .Z(_07465_));
 OR2_X1 _13057_ (.A1(_07268_),
    .A2(_07465_),
    .ZN(_07466_));
 MUX2_X1 _13058_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][36] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][36] ),
    .S(_05147_),
    .Z(_07467_));
 OAI21_X4 _13059_ (.A(_07466_),
    .B1(_07467_),
    .B2(_07272_),
    .ZN(_10261_));
 MUX2_X1 _13060_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][41] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][41] ),
    .S(_07440_),
    .Z(_07468_));
 OR2_X2 _13061_ (.A1(_07439_),
    .A2(_07468_),
    .ZN(_07469_));
 MUX2_X1 _13062_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][41] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][41] ),
    .S(_07443_),
    .Z(_07470_));
 OAI21_X4 _13063_ (.A(_07469_),
    .B1(_07446_),
    .B2(_07470_),
    .ZN(_10264_));
 MUX2_X1 _13064_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][40] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][40] ),
    .S(_05147_),
    .Z(_07471_));
 MUX2_X1 _13065_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][40] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][40] ),
    .S(_05147_),
    .Z(_07472_));
 MUX2_X2 _13066_ (.A(_07471_),
    .B(_07472_),
    .S(_05153_),
    .Z(_07473_));
 INV_X1 _13067_ (.A(_07473_),
    .ZN(_10267_));
 MUX2_X1 _13068_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][43] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][43] ),
    .S(_05310_),
    .Z(_07474_));
 OR2_X1 _13069_ (.A1(_05320_),
    .A2(_07474_),
    .ZN(_07475_));
 MUX2_X1 _13070_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][43] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][43] ),
    .S(_05312_),
    .Z(_07476_));
 OAI21_X4 _13071_ (.A(_07475_),
    .B1(_07476_),
    .B2(_05326_),
    .ZN(_10279_));
 MUX2_X1 _13072_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][44] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][44] ),
    .S(_05315_),
    .Z(_07477_));
 MUX2_X1 _13073_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][44] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][44] ),
    .S(_05315_),
    .Z(_07478_));
 MUX2_X2 _13074_ (.A(_07477_),
    .B(_07478_),
    .S(_05321_),
    .Z(_07479_));
 INV_X1 _13075_ (.A(_07479_),
    .ZN(_10282_));
 MUX2_X1 _13076_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][45] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][45] ),
    .S(_05314_),
    .Z(_07480_));
 OR2_X1 _13077_ (.A1(_05320_),
    .A2(_07480_),
    .ZN(_07481_));
 MUX2_X1 _13078_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][45] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][45] ),
    .S(_05312_),
    .Z(_07482_));
 OAI21_X4 _13079_ (.A(_07481_),
    .B1(_07482_),
    .B2(_05326_),
    .ZN(_10285_));
 MUX2_X1 _13080_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][46] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][46] ),
    .S(_05314_),
    .Z(_07483_));
 OR2_X1 _13081_ (.A1(_05321_),
    .A2(_07483_),
    .ZN(_07484_));
 MUX2_X1 _13082_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][46] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][46] ),
    .S(_05312_),
    .Z(_07485_));
 OAI21_X4 _13083_ (.A(_07484_),
    .B1(_07485_),
    .B2(_05326_),
    .ZN(_10288_));
 MUX2_X1 _13084_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][47] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][47] ),
    .S(_05312_),
    .Z(_07486_));
 MUX2_X1 _13085_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][47] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][47] ),
    .S(_05312_),
    .Z(_07487_));
 BUF_X4 _13086_ (.A(_05320_),
    .Z(_07488_));
 MUX2_X2 _13087_ (.A(_07486_),
    .B(_07487_),
    .S(_07488_),
    .Z(_07489_));
 INV_X1 _13088_ (.A(_07489_),
    .ZN(_10291_));
 MUX2_X1 _13089_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][48] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][48] ),
    .S(_05314_),
    .Z(_07490_));
 OR2_X1 _13090_ (.A1(_05321_),
    .A2(_07490_),
    .ZN(_07491_));
 MUX2_X1 _13091_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][48] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][48] ),
    .S(_05312_),
    .Z(_07492_));
 OAI21_X4 _13092_ (.A(_07491_),
    .B1(_07492_),
    .B2(_05326_),
    .ZN(_10294_));
 BUF_X4 _13093_ (.A(_07488_),
    .Z(_07493_));
 BUF_X16 _13094_ (.A(_05312_),
    .Z(_07494_));
 MUX2_X1 _13095_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][49] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][49] ),
    .S(_07494_),
    .Z(_07495_));
 OR2_X1 _13096_ (.A1(_07493_),
    .A2(_07495_),
    .ZN(_07496_));
 BUF_X16 _13097_ (.A(_05315_),
    .Z(_07497_));
 MUX2_X1 _13098_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][49] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][49] ),
    .S(_07497_),
    .Z(_07498_));
 BUF_X16 _13099_ (.A(_05326_),
    .Z(_07499_));
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 OAI21_X4 _13101_ (.A(_07496_),
    .B1(_07498_),
    .B2(_07499_),
    .ZN(_10297_));
 MUX2_X1 _13102_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][41] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][41] ),
    .S(_07494_),
    .Z(_07501_));
 OR2_X4 _13103_ (.A1(_07501_),
    .A2(_07493_),
    .ZN(_07502_));
 MUX2_X1 _13104_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][41] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][41] ),
    .S(_07497_),
    .Z(_07503_));
 OAI21_X4 _13105_ (.A(_07502_),
    .B1(_07499_),
    .B2(_07503_),
    .ZN(_10300_));
 MUX2_X1 _13106_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][40] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][40] ),
    .S(_05310_),
    .Z(_07504_));
 MUX2_X1 _13107_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][40] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][40] ),
    .S(_05310_),
    .Z(_07505_));
 MUX2_X2 _13108_ (.A(_07504_),
    .B(_07505_),
    .S(_05320_),
    .Z(_07506_));
 INV_X2 _13109_ (.A(_07506_),
    .ZN(_10303_));
 MUX2_X1 _13110_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][39] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][39] ),
    .S(_05315_),
    .Z(_07507_));
 MUX2_X1 _13111_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][39] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][39] ),
    .S(_05315_),
    .Z(_07508_));
 MUX2_X2 _13112_ (.A(_07507_),
    .B(_07508_),
    .S(_05321_),
    .Z(_07509_));
 INV_X2 _13113_ (.A(_07509_),
    .ZN(_10306_));
 MUX2_X1 _13114_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][38] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][38] ),
    .S(_05314_),
    .Z(_07510_));
 OR2_X1 _13115_ (.A1(_05321_),
    .A2(_07510_),
    .ZN(_07511_));
 MUX2_X1 _13116_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][38] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][38] ),
    .S(_05312_),
    .Z(_07512_));
 OAI21_X4 _13117_ (.A(_07511_),
    .B1(_07512_),
    .B2(_05326_),
    .ZN(_10309_));
 MUX2_X1 _13118_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][36] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][36] ),
    .S(net728),
    .Z(_07513_));
 OR2_X1 _13119_ (.A1(_05320_),
    .A2(_07513_),
    .ZN(_07514_));
 MUX2_X1 _13120_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][36] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][36] ),
    .S(_05314_),
    .Z(_07515_));
 OAI21_X4 _13121_ (.A(_07514_),
    .B1(_07515_),
    .B2(_05326_),
    .ZN(_10315_));
 MUX2_X1 _13122_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][35] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][35] ),
    .S(_05315_),
    .Z(_07516_));
 MUX2_X1 _13123_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][35] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][35] ),
    .S(_05315_),
    .Z(_07517_));
 MUX2_X2 _13124_ (.A(_07516_),
    .B(_07517_),
    .S(_05321_),
    .Z(_07518_));
 INV_X1 _13125_ (.A(_07518_),
    .ZN(_10318_));
 BUF_X2 _13126_ (.A(_05468_),
    .Z(_07519_));
 BUF_X16 _13127_ (.A(_07286_),
    .Z(_07520_));
 MUX2_X1 _13128_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][49] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][49] ),
    .S(_07520_),
    .Z(_07521_));
 OR2_X2 _13129_ (.A1(_07519_),
    .A2(_07521_),
    .ZN(_07522_));
 BUF_X8 _13130_ (.A(_05459_),
    .Z(_07523_));
 MUX2_X1 _13131_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][49] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][49] ),
    .S(_07523_),
    .Z(_07524_));
 BUF_X8 _13132_ (.A(_07290_),
    .Z(_07525_));
 BUF_X8 _13133_ (.A(_07525_),
    .Z(_07526_));
 OAI21_X4 _13134_ (.A(_07522_),
    .B1(_07526_),
    .B2(_07524_),
    .ZN(_10324_));
 MUX2_X1 _13135_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][48] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][48] ),
    .S(net720),
    .Z(_07527_));
 OR2_X1 _13136_ (.A1(_05463_),
    .A2(_07527_),
    .ZN(_07528_));
 MUX2_X1 _13137_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][48] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][48] ),
    .S(_07286_),
    .Z(_07529_));
 OAI21_X4 _13138_ (.A(_07528_),
    .B1(_07529_),
    .B2(_07290_),
    .ZN(_10327_));
 MUX2_X1 _13139_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][44] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][44] ),
    .S(_05458_),
    .Z(_07530_));
 OR2_X1 _13140_ (.A1(_05468_),
    .A2(_07530_),
    .ZN(_07531_));
 MUX2_X1 _13141_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][44] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][44] ),
    .S(net721),
    .Z(_07532_));
 OAI21_X4 _13142_ (.A(_07531_),
    .B1(_07532_),
    .B2(_07290_),
    .ZN(_10339_));
 MUX2_X1 _13143_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][36] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][36] ),
    .S(_05458_),
    .Z(_07533_));
 OR2_X1 _13144_ (.A1(_05463_),
    .A2(_07533_),
    .ZN(_07534_));
 MUX2_X1 _13145_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][36] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][36] ),
    .S(_07286_),
    .Z(_07535_));
 OAI21_X4 _13146_ (.A(_07534_),
    .B1(_07535_),
    .B2(_07290_),
    .ZN(_10357_));
 MUX2_X1 _13147_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][41] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][41] ),
    .S(_07520_),
    .Z(_07536_));
 OR2_X2 _13148_ (.A1(_07519_),
    .A2(_07536_),
    .ZN(_07537_));
 MUX2_X1 _13149_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][41] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][41] ),
    .S(_07523_),
    .Z(_07538_));
 OAI21_X4 _13150_ (.A(_07537_),
    .B1(_07538_),
    .B2(_07526_),
    .ZN(_10360_));
 MUX2_X1 _13151_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][40] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][40] ),
    .S(_05458_),
    .Z(_07539_));
 OR2_X2 _13152_ (.A1(_05468_),
    .A2(_07539_),
    .ZN(_07540_));
 MUX2_X1 _13153_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][40] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][40] ),
    .S(_07286_),
    .Z(_07541_));
 OAI21_X4 _13154_ (.A(_07540_),
    .B1(_07541_),
    .B2(_07290_),
    .ZN(_10363_));
 MUX2_X1 _13155_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][43] ),
    .S(_07312_),
    .Z(_07542_));
 MUX2_X1 _13156_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][43] ),
    .S(_07314_),
    .Z(_07543_));
 MUX2_X1 _13157_ (.A(_07542_),
    .B(_07543_),
    .S(_05729_),
    .Z(_07544_));
 MUX2_X1 _13158_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][43] ),
    .S(_07314_),
    .Z(_07545_));
 MUX2_X1 _13159_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][43] ),
    .S(_07348_),
    .Z(_07546_));
 MUX2_X1 _13160_ (.A(_07545_),
    .B(_07546_),
    .S(_07321_),
    .Z(_07547_));
 MUX2_X1 _13161_ (.A(_07544_),
    .B(_07547_),
    .S(_07323_),
    .Z(_07548_));
 MUX2_X1 _13162_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][43] ),
    .S(_07352_),
    .Z(_07549_));
 MUX2_X1 _13163_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][43] ),
    .S(_07328_),
    .Z(_07550_));
 MUX2_X1 _13164_ (.A(_07549_),
    .B(_07550_),
    .S(_07330_),
    .Z(_07551_));
 MUX2_X1 _13165_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][43] ),
    .S(_07332_),
    .Z(_07552_));
 MUX2_X1 _13166_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][43] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][43] ),
    .S(_07334_),
    .Z(_07553_));
 MUX2_X1 _13167_ (.A(_07552_),
    .B(_07553_),
    .S(_07358_),
    .Z(_07554_));
 MUX2_X1 _13168_ (.A(_07551_),
    .B(_07554_),
    .S(_07339_),
    .Z(_07555_));
 MUX2_X2 _13169_ (.A(_07548_),
    .B(_07555_),
    .S(_07341_),
    .Z(_07556_));
 INV_X1 _13170_ (.A(_07556_),
    .ZN(_10375_));
 MUX2_X1 _13171_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][44] ),
    .S(_05724_),
    .Z(_07557_));
 MUX2_X1 _13172_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][44] ),
    .S(_07344_),
    .Z(_07558_));
 MUX2_X1 _13173_ (.A(_07557_),
    .B(_07558_),
    .S(_05729_),
    .Z(_07559_));
 MUX2_X1 _13174_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][44] ),
    .S(_07344_),
    .Z(_07560_));
 MUX2_X1 _13175_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][44] ),
    .S(_07348_),
    .Z(_07561_));
 MUX2_X1 _13176_ (.A(_07560_),
    .B(_07561_),
    .S(_07316_),
    .Z(_07562_));
 MUX2_X1 _13177_ (.A(_07559_),
    .B(_07562_),
    .S(_05721_),
    .Z(_07563_));
 MUX2_X1 _13178_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][44] ),
    .S(_07352_),
    .Z(_07564_));
 MUX2_X1 _13179_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][44] ),
    .S(_07326_),
    .Z(_07565_));
 MUX2_X1 _13180_ (.A(_07564_),
    .B(_07565_),
    .S(_07330_),
    .Z(_07566_));
 MUX2_X1 _13181_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][44] ),
    .S(_07328_),
    .Z(_07567_));
 MUX2_X1 _13182_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][44] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][44] ),
    .S(_07334_),
    .Z(_07568_));
 MUX2_X1 _13183_ (.A(_07567_),
    .B(_07568_),
    .S(_07358_),
    .Z(_07569_));
 MUX2_X1 _13184_ (.A(_07566_),
    .B(_07569_),
    .S(_07339_),
    .Z(_07570_));
 MUX2_X2 _13185_ (.A(_07563_),
    .B(_07570_),
    .S(_07341_),
    .Z(_07571_));
 INV_X1 _13186_ (.A(_07571_),
    .ZN(_10381_));
 MUX2_X1 _13187_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][49] ),
    .S(_07319_),
    .Z(_07572_));
 MUX2_X1 _13188_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][49] ),
    .S(_07319_),
    .Z(_07573_));
 MUX2_X1 _13189_ (.A(_07572_),
    .B(_07573_),
    .S(_07321_),
    .Z(_07574_));
 MUX2_X1 _13190_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][49] ),
    .S(_07319_),
    .Z(_07575_));
 MUX2_X1 _13191_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][49] ),
    .S(_07352_),
    .Z(_07576_));
 MUX2_X1 _13192_ (.A(_07575_),
    .B(_07576_),
    .S(_07321_),
    .Z(_07577_));
 MUX2_X1 _13193_ (.A(_07574_),
    .B(_07577_),
    .S(_07323_),
    .Z(_07578_));
 MUX2_X1 _13194_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][49] ),
    .S(_07384_),
    .Z(_07579_));
 MUX2_X1 _13195_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][49] ),
    .S(_07384_),
    .Z(_07580_));
 MUX2_X1 _13196_ (.A(_07579_),
    .B(_07580_),
    .S(_07337_),
    .Z(_07581_));
 MUX2_X1 _13197_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][49] ),
    .S(_07384_),
    .Z(_07582_));
 MUX2_X1 _13198_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][49] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][49] ),
    .S(_07384_),
    .Z(_07583_));
 MUX2_X1 _13199_ (.A(_07582_),
    .B(_07583_),
    .S(_07337_),
    .Z(_07584_));
 MUX2_X1 _13200_ (.A(_07581_),
    .B(_07584_),
    .S(_07391_),
    .Z(_07585_));
 MUX2_X2 _13201_ (.A(_07578_),
    .B(_07585_),
    .S(_07393_),
    .Z(_07586_));
 INV_X1 _13202_ (.A(_07586_),
    .ZN(_10384_));
 MUX2_X1 _13203_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][48] ),
    .S(_05724_),
    .Z(_07587_));
 MUX2_X1 _13204_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][48] ),
    .S(_07312_),
    .Z(_07588_));
 MUX2_X1 _13205_ (.A(_07587_),
    .B(_07588_),
    .S(_05729_),
    .Z(_07589_));
 MUX2_X1 _13206_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][48] ),
    .S(_07344_),
    .Z(_07590_));
 MUX2_X1 _13207_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][48] ),
    .S(_07348_),
    .Z(_07591_));
 MUX2_X1 _13208_ (.A(_07590_),
    .B(_07591_),
    .S(_07316_),
    .Z(_07592_));
 MUX2_X1 _13209_ (.A(_07589_),
    .B(_07592_),
    .S(_05721_),
    .Z(_07593_));
 MUX2_X1 _13210_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][48] ),
    .S(_07352_),
    .Z(_07594_));
 MUX2_X1 _13211_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][48] ),
    .S(_07326_),
    .Z(_07595_));
 MUX2_X1 _13212_ (.A(_07594_),
    .B(_07595_),
    .S(_07330_),
    .Z(_07596_));
 MUX2_X1 _13213_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][48] ),
    .S(_07328_),
    .Z(_07597_));
 MUX2_X1 _13214_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][48] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][48] ),
    .S(_07332_),
    .Z(_07598_));
 MUX2_X1 _13215_ (.A(_07597_),
    .B(_07598_),
    .S(_07358_),
    .Z(_07599_));
 MUX2_X1 _13216_ (.A(_07596_),
    .B(_07599_),
    .S(_07339_),
    .Z(_07600_));
 MUX2_X2 _13217_ (.A(_07593_),
    .B(_07600_),
    .S(_07341_),
    .Z(_07601_));
 INV_X1 _13218_ (.A(_07601_),
    .ZN(_10387_));
 MUX2_X1 _13219_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][40] ),
    .S(_07312_),
    .Z(_07602_));
 MUX2_X1 _13220_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][40] ),
    .S(_07314_),
    .Z(_07603_));
 MUX2_X1 _13221_ (.A(_07602_),
    .B(_07603_),
    .S(_07316_),
    .Z(_07604_));
 MUX2_X1 _13222_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][40] ),
    .S(_07348_),
    .Z(_07605_));
 MUX2_X1 _13223_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][40] ),
    .S(_07319_),
    .Z(_07606_));
 MUX2_X1 _13224_ (.A(_07605_),
    .B(_07606_),
    .S(_07321_),
    .Z(_07607_));
 MUX2_X1 _13225_ (.A(_07604_),
    .B(_07607_),
    .S(_07323_),
    .Z(_07608_));
 MUX2_X1 _13226_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][40] ),
    .S(_07326_),
    .Z(_07609_));
 MUX2_X1 _13227_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][40] ),
    .S(_07332_),
    .Z(_07610_));
 MUX2_X1 _13228_ (.A(_07609_),
    .B(_07610_),
    .S(_07358_),
    .Z(_07611_));
 MUX2_X1 _13229_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][40] ),
    .S(_07332_),
    .Z(_07612_));
 MUX2_X1 _13230_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][40] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][40] ),
    .S(_07334_),
    .Z(_07613_));
 MUX2_X1 _13231_ (.A(_07612_),
    .B(_07613_),
    .S(_07337_),
    .Z(_07614_));
 MUX2_X1 _13232_ (.A(_07611_),
    .B(_07614_),
    .S(_07339_),
    .Z(_07615_));
 MUX2_X2 _13233_ (.A(_07608_),
    .B(_07615_),
    .S(_07341_),
    .Z(_07616_));
 INV_X1 _13234_ (.A(_07616_),
    .ZN(_10399_));
 MUX2_X1 _13235_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][39] ),
    .S(_07312_),
    .Z(_07617_));
 MUX2_X1 _13236_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][39] ),
    .S(_07344_),
    .Z(_07618_));
 MUX2_X1 _13237_ (.A(_07617_),
    .B(_07618_),
    .S(_05729_),
    .Z(_07619_));
 MUX2_X1 _13238_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][39] ),
    .S(_07314_),
    .Z(_07620_));
 MUX2_X1 _13239_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][39] ),
    .S(_07348_),
    .Z(_07621_));
 MUX2_X1 _13240_ (.A(_07620_),
    .B(_07621_),
    .S(_07321_),
    .Z(_07622_));
 MUX2_X1 _13241_ (.A(_07619_),
    .B(_07622_),
    .S(_07323_),
    .Z(_07623_));
 MUX2_X1 _13242_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][39] ),
    .S(_07352_),
    .Z(_07624_));
 MUX2_X1 _13243_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][39] ),
    .S(_07328_),
    .Z(_07625_));
 MUX2_X1 _13244_ (.A(_07624_),
    .B(_07625_),
    .S(_07330_),
    .Z(_07626_));
 MUX2_X1 _13245_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][39] ),
    .S(_07328_),
    .Z(_07627_));
 MUX2_X1 _13246_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][39] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][39] ),
    .S(_07334_),
    .Z(_07628_));
 MUX2_X1 _13247_ (.A(_07627_),
    .B(_07628_),
    .S(_07358_),
    .Z(_07629_));
 MUX2_X1 _13248_ (.A(_07626_),
    .B(_07629_),
    .S(_07339_),
    .Z(_07630_));
 MUX2_X2 _13249_ (.A(_07623_),
    .B(_07630_),
    .S(_07341_),
    .Z(_07631_));
 INV_X1 _13250_ (.A(_07631_),
    .ZN(_10402_));
 MUX2_X1 _13251_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][38] ),
    .S(_07312_),
    .Z(_07632_));
 MUX2_X1 _13252_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][38] ),
    .S(_07314_),
    .Z(_07633_));
 MUX2_X1 _13253_ (.A(_07632_),
    .B(_07633_),
    .S(_07316_),
    .Z(_07634_));
 MUX2_X1 _13254_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][38] ),
    .S(_07314_),
    .Z(_07635_));
 MUX2_X1 _13255_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][38] ),
    .S(_07319_),
    .Z(_07636_));
 MUX2_X1 _13256_ (.A(_07635_),
    .B(_07636_),
    .S(_07321_),
    .Z(_07637_));
 MUX2_X1 _13257_ (.A(_07634_),
    .B(_07637_),
    .S(_07323_),
    .Z(_07638_));
 MUX2_X1 _13258_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][38] ),
    .S(_07326_),
    .Z(_07639_));
 MUX2_X1 _13259_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][38] ),
    .S(_07332_),
    .Z(_07640_));
 MUX2_X1 _13260_ (.A(_07639_),
    .B(_07640_),
    .S(_07330_),
    .Z(_07641_));
 MUX2_X1 _13261_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][38] ),
    .S(_07332_),
    .Z(_07642_));
 MUX2_X1 _13262_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][38] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][38] ),
    .S(_07334_),
    .Z(_07643_));
 MUX2_X1 _13263_ (.A(_07642_),
    .B(_07643_),
    .S(_07337_),
    .Z(_07644_));
 MUX2_X1 _13264_ (.A(_07641_),
    .B(_07644_),
    .S(_07339_),
    .Z(_07645_));
 MUX2_X2 _13265_ (.A(_07638_),
    .B(_07645_),
    .S(_07341_),
    .Z(_07646_));
 INV_X1 _13266_ (.A(_07646_),
    .ZN(_10405_));
 MUX2_X1 _13267_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][36] ),
    .S(_05724_),
    .Z(_07647_));
 MUX2_X1 _13268_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][36] ),
    .S(_07312_),
    .Z(_07648_));
 MUX2_X1 _13269_ (.A(_07647_),
    .B(_07648_),
    .S(_05729_),
    .Z(_07649_));
 MUX2_X1 _13270_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][36] ),
    .S(_07344_),
    .Z(_07650_));
 MUX2_X1 _13271_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][36] ),
    .S(_07348_),
    .Z(_07651_));
 MUX2_X1 _13272_ (.A(_07650_),
    .B(_07651_),
    .S(_07316_),
    .Z(_07652_));
 MUX2_X1 _13273_ (.A(_07649_),
    .B(_07652_),
    .S(_05721_),
    .Z(_07653_));
 MUX2_X1 _13274_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][36] ),
    .S(_07352_),
    .Z(_07654_));
 MUX2_X1 _13275_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][36] ),
    .S(_07326_),
    .Z(_07655_));
 MUX2_X1 _13276_ (.A(_07654_),
    .B(_07655_),
    .S(_07330_),
    .Z(_07656_));
 MUX2_X1 _13277_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][36] ),
    .S(_07326_),
    .Z(_07657_));
 MUX2_X1 _13278_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][36] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][36] ),
    .S(_07332_),
    .Z(_07658_));
 MUX2_X1 _13279_ (.A(_07657_),
    .B(_07658_),
    .S(_07358_),
    .Z(_07659_));
 MUX2_X1 _13280_ (.A(_07656_),
    .B(_07659_),
    .S(_07323_),
    .Z(_07660_));
 MUX2_X2 _13281_ (.A(_07653_),
    .B(_07660_),
    .S(_05738_),
    .Z(_07661_));
 INV_X1 _13282_ (.A(_07661_),
    .ZN(_10411_));
 MUX2_X1 _13283_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][35] ),
    .S(_07312_),
    .Z(_07662_));
 MUX2_X1 _13284_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][35] ),
    .S(_07344_),
    .Z(_07663_));
 MUX2_X1 _13285_ (.A(_07662_),
    .B(_07663_),
    .S(_05729_),
    .Z(_07664_));
 MUX2_X1 _13286_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][35] ),
    .S(_07314_),
    .Z(_07665_));
 MUX2_X1 _13287_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][35] ),
    .S(_07348_),
    .Z(_07666_));
 MUX2_X1 _13288_ (.A(_07665_),
    .B(_07666_),
    .S(_07316_),
    .Z(_07667_));
 MUX2_X1 _13289_ (.A(_07664_),
    .B(_07667_),
    .S(_07323_),
    .Z(_07668_));
 MUX2_X1 _13290_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][35] ),
    .S(_07352_),
    .Z(_07669_));
 MUX2_X1 _13291_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][35] ),
    .S(_07328_),
    .Z(_07670_));
 MUX2_X1 _13292_ (.A(_07669_),
    .B(_07670_),
    .S(_07330_),
    .Z(_07671_));
 MUX2_X1 _13293_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][35] ),
    .S(_07328_),
    .Z(_07672_));
 MUX2_X1 _13294_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][35] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][35] ),
    .S(_07334_),
    .Z(_07673_));
 MUX2_X1 _13295_ (.A(_07672_),
    .B(_07673_),
    .S(_07358_),
    .Z(_07674_));
 MUX2_X1 _13296_ (.A(_07671_),
    .B(_07674_),
    .S(_07339_),
    .Z(_07675_));
 MUX2_X2 _13297_ (.A(_07668_),
    .B(_07675_),
    .S(_07341_),
    .Z(_07676_));
 INV_X1 _13298_ (.A(_07676_),
    .ZN(_10414_));
 BUF_X2 _13299_ (.A(net292),
    .Z(_07677_));
 INV_X1 _13300_ (.A(_07677_),
    .ZN(_10457_));
 INV_X2 _13301_ (.A(_10169_),
    .ZN(_10569_));
 INV_X1 _13302_ (.A(_10477_),
    .ZN(_10165_));
 INV_X1 _13303_ (.A(_10469_),
    .ZN(_10172_));
 INV_X1 _13304_ (.A(_10503_),
    .ZN(_10175_));
 INV_X1 _13305_ (.A(_10511_),
    .ZN(_10162_));
 NOR2_X4 _13306_ (.A1(_06540_),
    .A2(_10505_),
    .ZN(_07678_));
 NAND2_X1 _13307_ (.A1(_10577_),
    .A2(_07678_),
    .ZN(_07679_));
 BUF_X4 _13308_ (.A(_07679_),
    .Z(_07680_));
 BUF_X4 _13309_ (.A(_07680_),
    .Z(_07681_));
 MUX2_X1 _13310_ (.A(net3),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][0] ),
    .S(_07681_),
    .Z(_00093_));
 MUX2_X1 _13311_ (.A(net4),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][10] ),
    .S(_07681_),
    .Z(_00094_));
 MUX2_X1 _13312_ (.A(net5),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][11] ),
    .S(_07681_),
    .Z(_00095_));
 MUX2_X1 _13313_ (.A(net6),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][12] ),
    .S(_07681_),
    .Z(_00096_));
 MUX2_X1 _13314_ (.A(net7),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][13] ),
    .S(_07681_),
    .Z(_00097_));
 MUX2_X1 _13315_ (.A(net8),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][14] ),
    .S(_07681_),
    .Z(_00098_));
 MUX2_X1 _13316_ (.A(net9),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][15] ),
    .S(_07681_),
    .Z(_00099_));
 MUX2_X1 _13317_ (.A(net10),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][16] ),
    .S(_07681_),
    .Z(_00100_));
 MUX2_X1 _13318_ (.A(net11),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][17] ),
    .S(_07681_),
    .Z(_00101_));
 MUX2_X1 _13319_ (.A(net12),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][18] ),
    .S(_07681_),
    .Z(_00102_));
 BUF_X4 _13320_ (.A(_07680_),
    .Z(_07682_));
 MUX2_X1 _13321_ (.A(net13),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][19] ),
    .S(_07682_),
    .Z(_00103_));
 MUX2_X1 _13322_ (.A(net14),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][1] ),
    .S(_07682_),
    .Z(_00104_));
 MUX2_X1 _13323_ (.A(net15),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][20] ),
    .S(_07682_),
    .Z(_00105_));
 MUX2_X1 _13324_ (.A(net16),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][21] ),
    .S(_07682_),
    .Z(_00106_));
 MUX2_X1 _13325_ (.A(net17),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][22] ),
    .S(_07682_),
    .Z(_00107_));
 MUX2_X1 _13326_ (.A(net18),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][23] ),
    .S(_07682_),
    .Z(_00108_));
 MUX2_X1 _13327_ (.A(net19),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][24] ),
    .S(_07682_),
    .Z(_00109_));
 MUX2_X1 _13328_ (.A(net20),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][25] ),
    .S(_07682_),
    .Z(_00110_));
 MUX2_X1 _13329_ (.A(net21),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][26] ),
    .S(_07682_),
    .Z(_00111_));
 MUX2_X1 _13330_ (.A(net22),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][27] ),
    .S(_07682_),
    .Z(_00112_));
 BUF_X4 _13331_ (.A(_07680_),
    .Z(_07683_));
 MUX2_X1 _13332_ (.A(net23),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][28] ),
    .S(_07683_),
    .Z(_00113_));
 MUX2_X1 _13333_ (.A(net24),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][29] ),
    .S(_07683_),
    .Z(_00114_));
 MUX2_X1 _13334_ (.A(net25),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][2] ),
    .S(_07683_),
    .Z(_00115_));
 MUX2_X1 _13335_ (.A(net26),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][30] ),
    .S(_07683_),
    .Z(_00116_));
 MUX2_X1 _13336_ (.A(net27),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][31] ),
    .S(_07683_),
    .Z(_00117_));
 MUX2_X1 _13337_ (.A(net28),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][32] ),
    .S(_07683_),
    .Z(_00118_));
 MUX2_X1 _13338_ (.A(net29),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][33] ),
    .S(_07683_),
    .Z(_00119_));
 MUX2_X1 _13339_ (.A(net30),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][34] ),
    .S(_07683_),
    .Z(_00120_));
 MUX2_X1 _13340_ (.A(net31),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][35] ),
    .S(_07683_),
    .Z(_00121_));
 MUX2_X1 _13341_ (.A(net32),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][36] ),
    .S(_07683_),
    .Z(_00122_));
 BUF_X4 _13342_ (.A(_07680_),
    .Z(_07684_));
 MUX2_X1 _13343_ (.A(net33),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][37] ),
    .S(_07684_),
    .Z(_00123_));
 MUX2_X1 _13344_ (.A(net34),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][38] ),
    .S(_07684_),
    .Z(_00124_));
 MUX2_X1 _13345_ (.A(net35),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][39] ),
    .S(_07684_),
    .Z(_00125_));
 MUX2_X1 _13346_ (.A(net36),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][3] ),
    .S(_07684_),
    .Z(_00126_));
 MUX2_X1 _13347_ (.A(net37),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][40] ),
    .S(_07684_),
    .Z(_00127_));
 MUX2_X1 _13348_ (.A(net38),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][41] ),
    .S(_07684_),
    .Z(_00128_));
 MUX2_X1 _13349_ (.A(net39),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][42] ),
    .S(_07684_),
    .Z(_00129_));
 MUX2_X1 _13350_ (.A(net40),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][43] ),
    .S(_07684_),
    .Z(_00130_));
 MUX2_X1 _13351_ (.A(net41),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][44] ),
    .S(_07684_),
    .Z(_00131_));
 MUX2_X1 _13352_ (.A(net42),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][45] ),
    .S(_07684_),
    .Z(_00132_));
 BUF_X4 _13353_ (.A(_07680_),
    .Z(_07685_));
 MUX2_X1 _13354_ (.A(net43),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][46] ),
    .S(_07685_),
    .Z(_00133_));
 MUX2_X1 _13355_ (.A(net44),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][47] ),
    .S(_07685_),
    .Z(_00134_));
 MUX2_X1 _13356_ (.A(net45),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][48] ),
    .S(_07685_),
    .Z(_00135_));
 MUX2_X1 _13357_ (.A(net46),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][49] ),
    .S(_07685_),
    .Z(_00136_));
 MUX2_X1 _13358_ (.A(net47),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][4] ),
    .S(_07685_),
    .Z(_00137_));
 MUX2_X1 _13359_ (.A(net48),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][50] ),
    .S(_07685_),
    .Z(_00138_));
 MUX2_X1 _13360_ (.A(net49),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][51] ),
    .S(_07685_),
    .Z(_00139_));
 MUX2_X1 _13361_ (.A(net50),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][52] ),
    .S(_07685_),
    .Z(_00140_));
 MUX2_X1 _13362_ (.A(net51),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][53] ),
    .S(_07685_),
    .Z(_00141_));
 MUX2_X1 _13363_ (.A(net52),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][54] ),
    .S(_07685_),
    .Z(_00142_));
 BUF_X4 _13364_ (.A(_07680_),
    .Z(_07686_));
 MUX2_X1 _13365_ (.A(net53),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][55] ),
    .S(_07686_),
    .Z(_00143_));
 MUX2_X1 _13366_ (.A(net54),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][56] ),
    .S(_07686_),
    .Z(_00144_));
 MUX2_X1 _13367_ (.A(net55),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][57] ),
    .S(_07686_),
    .Z(_00145_));
 MUX2_X1 _13368_ (.A(net56),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][58] ),
    .S(_07686_),
    .Z(_00146_));
 MUX2_X1 _13369_ (.A(net57),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][59] ),
    .S(_07686_),
    .Z(_00147_));
 MUX2_X1 _13370_ (.A(net58),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][5] ),
    .S(_07686_),
    .Z(_00148_));
 MUX2_X1 _13371_ (.A(net59),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][60] ),
    .S(_07686_),
    .Z(_00149_));
 MUX2_X1 _13372_ (.A(net60),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][61] ),
    .S(_07686_),
    .Z(_00150_));
 MUX2_X1 _13373_ (.A(net61),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][62] ),
    .S(_07686_),
    .Z(_00151_));
 MUX2_X1 _13374_ (.A(net62),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][63] ),
    .S(_07686_),
    .Z(_00152_));
 MUX2_X1 _13375_ (.A(net63),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][6] ),
    .S(_07680_),
    .Z(_00153_));
 MUX2_X1 _13376_ (.A(net64),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][7] ),
    .S(_07680_),
    .Z(_00154_));
 MUX2_X1 _13377_ (.A(net65),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][8] ),
    .S(_07680_),
    .Z(_00155_));
 MUX2_X1 _13378_ (.A(net66),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[0][9] ),
    .S(_07680_),
    .Z(_00156_));
 NAND2_X1 _13379_ (.A1(_10580_),
    .A2(_07678_),
    .ZN(_07687_));
 BUF_X4 _13380_ (.A(_07687_),
    .Z(_07688_));
 CLKBUF_X3 _13381_ (.A(_07688_),
    .Z(_07689_));
 MUX2_X1 _13382_ (.A(net3),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][0] ),
    .S(_07689_),
    .Z(_00157_));
 MUX2_X1 _13383_ (.A(net4),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][10] ),
    .S(_07689_),
    .Z(_00158_));
 MUX2_X1 _13384_ (.A(net5),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][11] ),
    .S(_07689_),
    .Z(_00159_));
 MUX2_X1 _13385_ (.A(net6),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][12] ),
    .S(_07689_),
    .Z(_00160_));
 MUX2_X1 _13386_ (.A(net7),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][13] ),
    .S(_07689_),
    .Z(_00161_));
 MUX2_X1 _13387_ (.A(net8),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][14] ),
    .S(_07689_),
    .Z(_00162_));
 MUX2_X1 _13388_ (.A(net9),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][15] ),
    .S(_07689_),
    .Z(_00163_));
 MUX2_X1 _13389_ (.A(net10),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][16] ),
    .S(_07689_),
    .Z(_00164_));
 MUX2_X1 _13390_ (.A(net11),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][17] ),
    .S(_07689_),
    .Z(_00165_));
 MUX2_X1 _13391_ (.A(net12),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][18] ),
    .S(_07689_),
    .Z(_00166_));
 BUF_X4 _13392_ (.A(_07688_),
    .Z(_07690_));
 MUX2_X1 _13393_ (.A(net13),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][19] ),
    .S(_07690_),
    .Z(_00167_));
 MUX2_X1 _13394_ (.A(net14),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][1] ),
    .S(_07690_),
    .Z(_00168_));
 MUX2_X1 _13395_ (.A(net15),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][20] ),
    .S(_07690_),
    .Z(_00169_));
 MUX2_X1 _13396_ (.A(net16),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][21] ),
    .S(_07690_),
    .Z(_00170_));
 MUX2_X1 _13397_ (.A(net17),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][22] ),
    .S(_07690_),
    .Z(_00171_));
 MUX2_X1 _13398_ (.A(net18),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][23] ),
    .S(_07690_),
    .Z(_00172_));
 MUX2_X1 _13399_ (.A(net19),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][24] ),
    .S(_07690_),
    .Z(_00173_));
 MUX2_X1 _13400_ (.A(net20),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][25] ),
    .S(_07690_),
    .Z(_00174_));
 MUX2_X1 _13401_ (.A(net21),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][26] ),
    .S(_07690_),
    .Z(_00175_));
 MUX2_X1 _13402_ (.A(net22),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][27] ),
    .S(_07690_),
    .Z(_00176_));
 BUF_X4 _13403_ (.A(_07688_),
    .Z(_07691_));
 MUX2_X1 _13404_ (.A(net23),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][28] ),
    .S(_07691_),
    .Z(_00177_));
 MUX2_X1 _13405_ (.A(net24),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][29] ),
    .S(_07691_),
    .Z(_00178_));
 MUX2_X1 _13406_ (.A(net25),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][2] ),
    .S(_07691_),
    .Z(_00179_));
 MUX2_X1 _13407_ (.A(net26),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][30] ),
    .S(_07691_),
    .Z(_00180_));
 MUX2_X1 _13408_ (.A(net27),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][31] ),
    .S(_07691_),
    .Z(_00181_));
 MUX2_X1 _13409_ (.A(net28),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][32] ),
    .S(_07691_),
    .Z(_00182_));
 MUX2_X1 _13410_ (.A(net29),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][33] ),
    .S(_07691_),
    .Z(_00183_));
 MUX2_X1 _13411_ (.A(net30),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][34] ),
    .S(_07691_),
    .Z(_00184_));
 MUX2_X1 _13412_ (.A(net31),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][35] ),
    .S(_07691_),
    .Z(_00185_));
 MUX2_X1 _13413_ (.A(net32),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][36] ),
    .S(_07691_),
    .Z(_00186_));
 BUF_X4 _13414_ (.A(_07688_),
    .Z(_07692_));
 MUX2_X1 _13415_ (.A(net33),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][37] ),
    .S(_07692_),
    .Z(_00187_));
 MUX2_X1 _13416_ (.A(net34),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][38] ),
    .S(_07692_),
    .Z(_00188_));
 MUX2_X1 _13417_ (.A(net35),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][39] ),
    .S(_07692_),
    .Z(_00189_));
 MUX2_X1 _13418_ (.A(net36),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][3] ),
    .S(_07692_),
    .Z(_00190_));
 MUX2_X1 _13419_ (.A(net37),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][40] ),
    .S(_07692_),
    .Z(_00191_));
 MUX2_X1 _13420_ (.A(net38),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][41] ),
    .S(_07692_),
    .Z(_00192_));
 MUX2_X1 _13421_ (.A(net39),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][42] ),
    .S(_07692_),
    .Z(_00193_));
 MUX2_X1 _13422_ (.A(net40),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][43] ),
    .S(_07692_),
    .Z(_00194_));
 MUX2_X1 _13423_ (.A(net41),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][44] ),
    .S(_07692_),
    .Z(_00195_));
 MUX2_X1 _13424_ (.A(net42),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][45] ),
    .S(_07692_),
    .Z(_00196_));
 BUF_X4 _13425_ (.A(_07688_),
    .Z(_07693_));
 MUX2_X1 _13426_ (.A(net43),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][46] ),
    .S(_07693_),
    .Z(_00197_));
 MUX2_X1 _13427_ (.A(net44),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][47] ),
    .S(_07693_),
    .Z(_00198_));
 MUX2_X1 _13428_ (.A(net45),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][48] ),
    .S(_07693_),
    .Z(_00199_));
 MUX2_X1 _13429_ (.A(net46),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][49] ),
    .S(_07693_),
    .Z(_00200_));
 MUX2_X1 _13430_ (.A(net47),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][4] ),
    .S(_07693_),
    .Z(_00201_));
 MUX2_X1 _13431_ (.A(net48),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][50] ),
    .S(_07693_),
    .Z(_00202_));
 MUX2_X1 _13432_ (.A(net49),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][51] ),
    .S(_07693_),
    .Z(_00203_));
 MUX2_X1 _13433_ (.A(net50),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][52] ),
    .S(_07693_),
    .Z(_00204_));
 MUX2_X1 _13434_ (.A(net51),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][53] ),
    .S(_07693_),
    .Z(_00205_));
 MUX2_X1 _13435_ (.A(net52),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][54] ),
    .S(_07693_),
    .Z(_00206_));
 BUF_X4 _13436_ (.A(_07688_),
    .Z(_07694_));
 MUX2_X1 _13437_ (.A(net53),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][55] ),
    .S(_07694_),
    .Z(_00207_));
 MUX2_X1 _13438_ (.A(net54),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][56] ),
    .S(_07694_),
    .Z(_00208_));
 MUX2_X1 _13439_ (.A(net55),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][57] ),
    .S(_07694_),
    .Z(_00209_));
 MUX2_X1 _13440_ (.A(net56),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][58] ),
    .S(_07694_),
    .Z(_00210_));
 MUX2_X1 _13441_ (.A(net57),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][59] ),
    .S(_07694_),
    .Z(_00211_));
 MUX2_X1 _13442_ (.A(net58),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][5] ),
    .S(_07694_),
    .Z(_00212_));
 MUX2_X1 _13443_ (.A(net59),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][60] ),
    .S(_07694_),
    .Z(_00213_));
 MUX2_X1 _13444_ (.A(net60),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][61] ),
    .S(_07694_),
    .Z(_00214_));
 MUX2_X1 _13445_ (.A(net61),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][62] ),
    .S(_07694_),
    .Z(_00215_));
 MUX2_X1 _13446_ (.A(net62),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][63] ),
    .S(_07694_),
    .Z(_00216_));
 MUX2_X1 _13447_ (.A(net63),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][6] ),
    .S(_07688_),
    .Z(_00217_));
 MUX2_X1 _13448_ (.A(net64),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][7] ),
    .S(_07688_),
    .Z(_00218_));
 MUX2_X1 _13449_ (.A(net65),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][8] ),
    .S(_07688_),
    .Z(_00219_));
 MUX2_X1 _13450_ (.A(net66),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[1][9] ),
    .S(_07688_),
    .Z(_00220_));
 NAND2_X1 _13451_ (.A1(_10578_),
    .A2(_07678_),
    .ZN(_07695_));
 BUF_X4 _13452_ (.A(_07695_),
    .Z(_07696_));
 BUF_X4 _13453_ (.A(_07696_),
    .Z(_07697_));
 MUX2_X1 _13454_ (.A(net3),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][0] ),
    .S(_07697_),
    .Z(_00221_));
 MUX2_X1 _13455_ (.A(net4),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][10] ),
    .S(_07697_),
    .Z(_00222_));
 MUX2_X1 _13456_ (.A(net5),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][11] ),
    .S(_07697_),
    .Z(_00223_));
 MUX2_X1 _13457_ (.A(net6),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][12] ),
    .S(_07697_),
    .Z(_00224_));
 MUX2_X1 _13458_ (.A(net7),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][13] ),
    .S(_07697_),
    .Z(_00225_));
 MUX2_X1 _13459_ (.A(net8),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][14] ),
    .S(_07697_),
    .Z(_00226_));
 MUX2_X1 _13460_ (.A(net9),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][15] ),
    .S(_07697_),
    .Z(_00227_));
 MUX2_X1 _13461_ (.A(net10),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][16] ),
    .S(_07697_),
    .Z(_00228_));
 MUX2_X1 _13462_ (.A(net11),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][17] ),
    .S(_07697_),
    .Z(_00229_));
 MUX2_X1 _13463_ (.A(net12),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][18] ),
    .S(_07697_),
    .Z(_00230_));
 BUF_X4 _13464_ (.A(_07696_),
    .Z(_07698_));
 MUX2_X1 _13465_ (.A(net13),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][19] ),
    .S(_07698_),
    .Z(_00231_));
 MUX2_X1 _13466_ (.A(net14),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][1] ),
    .S(_07698_),
    .Z(_00232_));
 MUX2_X1 _13467_ (.A(net15),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][20] ),
    .S(_07698_),
    .Z(_00233_));
 MUX2_X1 _13468_ (.A(net16),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][21] ),
    .S(_07698_),
    .Z(_00234_));
 MUX2_X1 _13469_ (.A(net17),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][22] ),
    .S(_07698_),
    .Z(_00235_));
 MUX2_X1 _13470_ (.A(net18),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][23] ),
    .S(_07698_),
    .Z(_00236_));
 MUX2_X1 _13471_ (.A(net19),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][24] ),
    .S(_07698_),
    .Z(_00237_));
 MUX2_X1 _13472_ (.A(net20),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][25] ),
    .S(_07698_),
    .Z(_00238_));
 MUX2_X1 _13473_ (.A(net21),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][26] ),
    .S(_07698_),
    .Z(_00239_));
 MUX2_X1 _13474_ (.A(net22),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][27] ),
    .S(_07698_),
    .Z(_00240_));
 CLKBUF_X3 _13475_ (.A(_07696_),
    .Z(_07699_));
 MUX2_X1 _13476_ (.A(net23),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][28] ),
    .S(_07699_),
    .Z(_00241_));
 MUX2_X1 _13477_ (.A(net24),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][29] ),
    .S(_07699_),
    .Z(_00242_));
 MUX2_X1 _13478_ (.A(net25),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][2] ),
    .S(_07699_),
    .Z(_00243_));
 MUX2_X1 _13479_ (.A(net26),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][30] ),
    .S(_07699_),
    .Z(_00244_));
 MUX2_X1 _13480_ (.A(net27),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][31] ),
    .S(_07699_),
    .Z(_00245_));
 MUX2_X1 _13481_ (.A(net28),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][32] ),
    .S(_07699_),
    .Z(_00246_));
 MUX2_X1 _13482_ (.A(net29),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][33] ),
    .S(_07699_),
    .Z(_00247_));
 MUX2_X1 _13483_ (.A(net30),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][34] ),
    .S(_07699_),
    .Z(_00248_));
 MUX2_X1 _13484_ (.A(net31),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][35] ),
    .S(_07699_),
    .Z(_00249_));
 MUX2_X1 _13485_ (.A(net32),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][36] ),
    .S(_07699_),
    .Z(_00250_));
 BUF_X4 _13486_ (.A(_07696_),
    .Z(_07700_));
 MUX2_X1 _13487_ (.A(net33),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][37] ),
    .S(_07700_),
    .Z(_00251_));
 MUX2_X1 _13488_ (.A(net34),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][38] ),
    .S(_07700_),
    .Z(_00252_));
 MUX2_X1 _13489_ (.A(net35),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][39] ),
    .S(_07700_),
    .Z(_00253_));
 MUX2_X1 _13490_ (.A(net36),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][3] ),
    .S(_07700_),
    .Z(_00254_));
 MUX2_X1 _13491_ (.A(net37),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][40] ),
    .S(_07700_),
    .Z(_00255_));
 MUX2_X1 _13492_ (.A(net38),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][41] ),
    .S(_07700_),
    .Z(_00256_));
 MUX2_X1 _13493_ (.A(net39),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][42] ),
    .S(_07700_),
    .Z(_00257_));
 MUX2_X1 _13494_ (.A(net40),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][43] ),
    .S(_07700_),
    .Z(_00258_));
 MUX2_X1 _13495_ (.A(net41),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][44] ),
    .S(_07700_),
    .Z(_00259_));
 MUX2_X1 _13496_ (.A(net42),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][45] ),
    .S(_07700_),
    .Z(_00260_));
 BUF_X4 _13497_ (.A(_07696_),
    .Z(_07701_));
 MUX2_X1 _13498_ (.A(net43),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][46] ),
    .S(_07701_),
    .Z(_00261_));
 MUX2_X1 _13499_ (.A(net44),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][47] ),
    .S(_07701_),
    .Z(_00262_));
 MUX2_X1 _13500_ (.A(net45),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][48] ),
    .S(_07701_),
    .Z(_00263_));
 MUX2_X1 _13501_ (.A(net46),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][49] ),
    .S(_07701_),
    .Z(_00264_));
 MUX2_X1 _13502_ (.A(net47),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][4] ),
    .S(_07701_),
    .Z(_00265_));
 MUX2_X1 _13503_ (.A(net48),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][50] ),
    .S(_07701_),
    .Z(_00266_));
 MUX2_X1 _13504_ (.A(net49),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][51] ),
    .S(_07701_),
    .Z(_00267_));
 MUX2_X1 _13505_ (.A(net50),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][52] ),
    .S(_07701_),
    .Z(_00268_));
 MUX2_X1 _13506_ (.A(net51),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][53] ),
    .S(_07701_),
    .Z(_00269_));
 MUX2_X1 _13507_ (.A(net52),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][54] ),
    .S(_07701_),
    .Z(_00270_));
 BUF_X4 _13508_ (.A(_07696_),
    .Z(_07702_));
 MUX2_X1 _13509_ (.A(net53),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][55] ),
    .S(_07702_),
    .Z(_00271_));
 MUX2_X1 _13510_ (.A(net54),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][56] ),
    .S(_07702_),
    .Z(_00272_));
 MUX2_X1 _13511_ (.A(net55),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][57] ),
    .S(_07702_),
    .Z(_00273_));
 MUX2_X1 _13512_ (.A(net56),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][58] ),
    .S(_07702_),
    .Z(_00274_));
 MUX2_X1 _13513_ (.A(net57),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][59] ),
    .S(_07702_),
    .Z(_00275_));
 MUX2_X1 _13514_ (.A(net58),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][5] ),
    .S(_07702_),
    .Z(_00276_));
 MUX2_X1 _13515_ (.A(net59),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][60] ),
    .S(_07702_),
    .Z(_00277_));
 MUX2_X1 _13516_ (.A(net60),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][61] ),
    .S(_07702_),
    .Z(_00278_));
 MUX2_X1 _13517_ (.A(net61),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][62] ),
    .S(_07702_),
    .Z(_00279_));
 MUX2_X1 _13518_ (.A(net62),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][63] ),
    .S(_07702_),
    .Z(_00280_));
 MUX2_X1 _13519_ (.A(net63),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][6] ),
    .S(_07696_),
    .Z(_00281_));
 MUX2_X1 _13520_ (.A(net64),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][7] ),
    .S(_07696_),
    .Z(_00282_));
 MUX2_X1 _13521_ (.A(net65),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][8] ),
    .S(_07696_),
    .Z(_00283_));
 MUX2_X1 _13522_ (.A(net66),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][9] ),
    .S(_07696_),
    .Z(_00284_));
 NAND2_X1 _13523_ (.A1(_10582_),
    .A2(_07678_),
    .ZN(_07703_));
 BUF_X4 _13524_ (.A(_07703_),
    .Z(_07704_));
 CLKBUF_X3 _13525_ (.A(_07704_),
    .Z(_07705_));
 MUX2_X1 _13526_ (.A(net3),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][0] ),
    .S(_07705_),
    .Z(_00285_));
 MUX2_X1 _13527_ (.A(net4),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][10] ),
    .S(_07705_),
    .Z(_00286_));
 MUX2_X1 _13528_ (.A(net5),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][11] ),
    .S(_07705_),
    .Z(_00287_));
 MUX2_X1 _13529_ (.A(net6),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][12] ),
    .S(_07705_),
    .Z(_00288_));
 MUX2_X1 _13530_ (.A(net7),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][13] ),
    .S(_07705_),
    .Z(_00289_));
 MUX2_X1 _13531_ (.A(net8),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][14] ),
    .S(_07705_),
    .Z(_00290_));
 MUX2_X1 _13532_ (.A(net9),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][15] ),
    .S(_07705_),
    .Z(_00291_));
 MUX2_X1 _13533_ (.A(net10),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][16] ),
    .S(_07705_),
    .Z(_00292_));
 MUX2_X1 _13534_ (.A(net11),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][17] ),
    .S(_07705_),
    .Z(_00293_));
 MUX2_X1 _13535_ (.A(net12),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][18] ),
    .S(_07705_),
    .Z(_00294_));
 BUF_X4 _13536_ (.A(_07704_),
    .Z(_07706_));
 MUX2_X1 _13537_ (.A(net13),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][19] ),
    .S(_07706_),
    .Z(_00295_));
 MUX2_X1 _13538_ (.A(net14),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][1] ),
    .S(_07706_),
    .Z(_00296_));
 MUX2_X1 _13539_ (.A(net15),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][20] ),
    .S(_07706_),
    .Z(_00297_));
 MUX2_X1 _13540_ (.A(net16),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][21] ),
    .S(_07706_),
    .Z(_00298_));
 MUX2_X1 _13541_ (.A(net17),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][22] ),
    .S(_07706_),
    .Z(_00299_));
 MUX2_X1 _13542_ (.A(net18),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][23] ),
    .S(_07706_),
    .Z(_00300_));
 MUX2_X1 _13543_ (.A(net19),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][24] ),
    .S(_07706_),
    .Z(_00301_));
 MUX2_X1 _13544_ (.A(net20),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][25] ),
    .S(_07706_),
    .Z(_00302_));
 MUX2_X1 _13545_ (.A(net21),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][26] ),
    .S(_07706_),
    .Z(_00303_));
 MUX2_X1 _13546_ (.A(net22),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][27] ),
    .S(_07706_),
    .Z(_00304_));
 BUF_X4 _13547_ (.A(_07704_),
    .Z(_07707_));
 MUX2_X1 _13548_ (.A(net23),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][28] ),
    .S(_07707_),
    .Z(_00305_));
 MUX2_X1 _13549_ (.A(net24),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][29] ),
    .S(_07707_),
    .Z(_00306_));
 MUX2_X1 _13550_ (.A(net25),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][2] ),
    .S(_07707_),
    .Z(_00307_));
 MUX2_X1 _13551_ (.A(net26),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][30] ),
    .S(_07707_),
    .Z(_00308_));
 MUX2_X1 _13552_ (.A(net27),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][31] ),
    .S(_07707_),
    .Z(_00309_));
 MUX2_X1 _13553_ (.A(net28),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][32] ),
    .S(_07707_),
    .Z(_00310_));
 MUX2_X1 _13554_ (.A(net29),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][33] ),
    .S(_07707_),
    .Z(_00311_));
 MUX2_X1 _13555_ (.A(net30),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][34] ),
    .S(_07707_),
    .Z(_00312_));
 MUX2_X1 _13556_ (.A(net31),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][35] ),
    .S(_07707_),
    .Z(_00313_));
 MUX2_X1 _13557_ (.A(net32),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][36] ),
    .S(_07707_),
    .Z(_00314_));
 BUF_X4 _13558_ (.A(_07704_),
    .Z(_07708_));
 MUX2_X1 _13559_ (.A(net33),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][37] ),
    .S(_07708_),
    .Z(_00315_));
 MUX2_X1 _13560_ (.A(net34),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][38] ),
    .S(_07708_),
    .Z(_00316_));
 MUX2_X1 _13561_ (.A(net35),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][39] ),
    .S(_07708_),
    .Z(_00317_));
 MUX2_X1 _13562_ (.A(net36),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][3] ),
    .S(_07708_),
    .Z(_00318_));
 MUX2_X1 _13563_ (.A(net37),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][40] ),
    .S(_07708_),
    .Z(_00319_));
 MUX2_X1 _13564_ (.A(net38),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][41] ),
    .S(_07708_),
    .Z(_00320_));
 MUX2_X1 _13565_ (.A(net39),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][42] ),
    .S(_07708_),
    .Z(_00321_));
 MUX2_X1 _13566_ (.A(net40),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][43] ),
    .S(_07708_),
    .Z(_00322_));
 MUX2_X1 _13567_ (.A(net41),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][44] ),
    .S(_07708_),
    .Z(_00323_));
 MUX2_X1 _13568_ (.A(net42),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][45] ),
    .S(_07708_),
    .Z(_00324_));
 BUF_X4 _13569_ (.A(_07704_),
    .Z(_07709_));
 MUX2_X1 _13570_ (.A(net43),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][46] ),
    .S(_07709_),
    .Z(_00325_));
 MUX2_X1 _13571_ (.A(net44),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][47] ),
    .S(_07709_),
    .Z(_00326_));
 MUX2_X1 _13572_ (.A(net45),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][48] ),
    .S(_07709_),
    .Z(_00327_));
 MUX2_X1 _13573_ (.A(net46),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][49] ),
    .S(_07709_),
    .Z(_00328_));
 MUX2_X1 _13574_ (.A(net47),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][4] ),
    .S(_07709_),
    .Z(_00329_));
 MUX2_X1 _13575_ (.A(net48),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][50] ),
    .S(_07709_),
    .Z(_00330_));
 MUX2_X1 _13576_ (.A(net49),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][51] ),
    .S(_07709_),
    .Z(_00331_));
 MUX2_X1 _13577_ (.A(net50),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][52] ),
    .S(_07709_),
    .Z(_00332_));
 MUX2_X1 _13578_ (.A(net51),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][53] ),
    .S(_07709_),
    .Z(_00333_));
 MUX2_X1 _13579_ (.A(net52),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][54] ),
    .S(_07709_),
    .Z(_00334_));
 BUF_X4 _13580_ (.A(_07704_),
    .Z(_07710_));
 MUX2_X1 _13581_ (.A(net53),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][55] ),
    .S(_07710_),
    .Z(_00335_));
 MUX2_X1 _13582_ (.A(net54),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][56] ),
    .S(_07710_),
    .Z(_00336_));
 MUX2_X1 _13583_ (.A(net55),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][57] ),
    .S(_07710_),
    .Z(_00337_));
 MUX2_X1 _13584_ (.A(net56),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][58] ),
    .S(_07710_),
    .Z(_00338_));
 MUX2_X1 _13585_ (.A(net57),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][59] ),
    .S(_07710_),
    .Z(_00339_));
 MUX2_X1 _13586_ (.A(net58),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][5] ),
    .S(_07710_),
    .Z(_00340_));
 MUX2_X1 _13587_ (.A(net59),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][60] ),
    .S(_07710_),
    .Z(_00341_));
 MUX2_X1 _13588_ (.A(net60),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][61] ),
    .S(_07710_),
    .Z(_00342_));
 MUX2_X1 _13589_ (.A(net61),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][62] ),
    .S(_07710_),
    .Z(_00343_));
 MUX2_X1 _13590_ (.A(net62),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][63] ),
    .S(_07710_),
    .Z(_00344_));
 MUX2_X1 _13591_ (.A(net63),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][6] ),
    .S(_07704_),
    .Z(_00345_));
 MUX2_X1 _13592_ (.A(net64),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][7] ),
    .S(_07704_),
    .Z(_00346_));
 MUX2_X1 _13593_ (.A(net65),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][8] ),
    .S(_07704_),
    .Z(_00347_));
 MUX2_X1 _13594_ (.A(net66),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][9] ),
    .S(_07704_),
    .Z(_00348_));
 NOR2_X2 _13595_ (.A1(_06540_),
    .A2(_10471_),
    .ZN(_07711_));
 NAND2_X1 _13596_ (.A1(_10585_),
    .A2(_07711_),
    .ZN(_07712_));
 BUF_X4 _13597_ (.A(_07712_),
    .Z(_07713_));
 CLKBUF_X3 _13598_ (.A(_07713_),
    .Z(_07714_));
 MUX2_X1 _13599_ (.A(net67),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][0] ),
    .S(_07714_),
    .Z(_00404_));
 MUX2_X1 _13600_ (.A(net68),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][10] ),
    .S(_07714_),
    .Z(_00405_));
 MUX2_X1 _13601_ (.A(net69),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][11] ),
    .S(_07714_),
    .Z(_00406_));
 MUX2_X1 _13602_ (.A(net70),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][12] ),
    .S(_07714_),
    .Z(_00407_));
 MUX2_X1 _13603_ (.A(net71),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][13] ),
    .S(_07714_),
    .Z(_00408_));
 MUX2_X1 _13604_ (.A(net72),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][14] ),
    .S(_07714_),
    .Z(_00409_));
 MUX2_X1 _13605_ (.A(net73),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][15] ),
    .S(_07714_),
    .Z(_00410_));
 MUX2_X1 _13606_ (.A(net74),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][16] ),
    .S(_07714_),
    .Z(_00411_));
 MUX2_X1 _13607_ (.A(net75),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][17] ),
    .S(_07714_),
    .Z(_00412_));
 MUX2_X1 _13608_ (.A(net76),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][18] ),
    .S(_07714_),
    .Z(_00413_));
 BUF_X4 _13609_ (.A(_07713_),
    .Z(_07715_));
 MUX2_X1 _13610_ (.A(net77),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][19] ),
    .S(_07715_),
    .Z(_00414_));
 MUX2_X1 _13611_ (.A(net78),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][1] ),
    .S(_07715_),
    .Z(_00415_));
 MUX2_X1 _13612_ (.A(net79),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][20] ),
    .S(_07715_),
    .Z(_00416_));
 MUX2_X1 _13613_ (.A(net80),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][21] ),
    .S(_07715_),
    .Z(_00417_));
 MUX2_X1 _13614_ (.A(net81),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][22] ),
    .S(_07715_),
    .Z(_00418_));
 MUX2_X1 _13615_ (.A(net82),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][23] ),
    .S(_07715_),
    .Z(_00419_));
 MUX2_X1 _13616_ (.A(net83),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][24] ),
    .S(_07715_),
    .Z(_00420_));
 MUX2_X1 _13617_ (.A(net84),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][25] ),
    .S(_07715_),
    .Z(_00421_));
 MUX2_X1 _13618_ (.A(net85),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][26] ),
    .S(_07715_),
    .Z(_00422_));
 MUX2_X1 _13619_ (.A(net86),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][27] ),
    .S(_07715_),
    .Z(_00423_));
 BUF_X4 _13620_ (.A(_07713_),
    .Z(_07716_));
 MUX2_X1 _13621_ (.A(net87),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][28] ),
    .S(_07716_),
    .Z(_00424_));
 MUX2_X1 _13622_ (.A(net88),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][29] ),
    .S(_07716_),
    .Z(_00425_));
 MUX2_X1 _13623_ (.A(net89),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][2] ),
    .S(_07716_),
    .Z(_00426_));
 MUX2_X1 _13624_ (.A(net90),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][30] ),
    .S(_07716_),
    .Z(_00427_));
 MUX2_X1 _13625_ (.A(net91),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][31] ),
    .S(_07716_),
    .Z(_00428_));
 MUX2_X1 _13626_ (.A(net92),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][32] ),
    .S(_07716_),
    .Z(_00429_));
 MUX2_X1 _13627_ (.A(net93),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][33] ),
    .S(_07716_),
    .Z(_00430_));
 MUX2_X1 _13628_ (.A(net94),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][34] ),
    .S(_07716_),
    .Z(_00431_));
 MUX2_X1 _13629_ (.A(net95),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][35] ),
    .S(_07716_),
    .Z(_00432_));
 MUX2_X1 _13630_ (.A(net96),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][36] ),
    .S(_07716_),
    .Z(_00433_));
 BUF_X4 _13631_ (.A(_07713_),
    .Z(_07717_));
 MUX2_X1 _13632_ (.A(net97),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][37] ),
    .S(_07717_),
    .Z(_00434_));
 MUX2_X1 _13633_ (.A(net98),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][38] ),
    .S(_07717_),
    .Z(_00435_));
 MUX2_X1 _13634_ (.A(net99),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][39] ),
    .S(_07717_),
    .Z(_00436_));
 MUX2_X1 _13635_ (.A(net100),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][3] ),
    .S(_07717_),
    .Z(_00437_));
 MUX2_X1 _13636_ (.A(net101),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][40] ),
    .S(_07717_),
    .Z(_00438_));
 MUX2_X1 _13637_ (.A(net102),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][41] ),
    .S(_07717_),
    .Z(_00439_));
 MUX2_X1 _13638_ (.A(net103),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][42] ),
    .S(_07717_),
    .Z(_00440_));
 MUX2_X1 _13639_ (.A(net104),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][43] ),
    .S(_07717_),
    .Z(_00441_));
 MUX2_X1 _13640_ (.A(net105),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][44] ),
    .S(_07717_),
    .Z(_00442_));
 MUX2_X1 _13641_ (.A(net106),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][45] ),
    .S(_07717_),
    .Z(_00443_));
 BUF_X4 _13642_ (.A(_07713_),
    .Z(_07718_));
 MUX2_X1 _13643_ (.A(net107),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][46] ),
    .S(_07718_),
    .Z(_00444_));
 MUX2_X1 _13644_ (.A(net108),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][47] ),
    .S(_07718_),
    .Z(_00445_));
 MUX2_X1 _13645_ (.A(net109),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][48] ),
    .S(_07718_),
    .Z(_00446_));
 MUX2_X1 _13646_ (.A(net110),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][49] ),
    .S(_07718_),
    .Z(_00447_));
 MUX2_X1 _13647_ (.A(net111),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][4] ),
    .S(_07718_),
    .Z(_00448_));
 MUX2_X1 _13648_ (.A(net112),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][50] ),
    .S(_07718_),
    .Z(_00449_));
 MUX2_X1 _13649_ (.A(net113),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][51] ),
    .S(_07718_),
    .Z(_00450_));
 MUX2_X1 _13650_ (.A(net114),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][52] ),
    .S(_07718_),
    .Z(_00451_));
 MUX2_X1 _13651_ (.A(net115),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][53] ),
    .S(_07718_),
    .Z(_00452_));
 MUX2_X1 _13652_ (.A(net116),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][54] ),
    .S(_07718_),
    .Z(_00453_));
 BUF_X4 _13653_ (.A(_07713_),
    .Z(_07719_));
 MUX2_X1 _13654_ (.A(net117),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][55] ),
    .S(_07719_),
    .Z(_00454_));
 MUX2_X1 _13655_ (.A(net118),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][56] ),
    .S(_07719_),
    .Z(_00455_));
 MUX2_X1 _13656_ (.A(net119),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][57] ),
    .S(_07719_),
    .Z(_00456_));
 MUX2_X1 _13657_ (.A(net120),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][58] ),
    .S(_07719_),
    .Z(_00457_));
 MUX2_X1 _13658_ (.A(net121),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][59] ),
    .S(_07719_),
    .Z(_00458_));
 MUX2_X1 _13659_ (.A(net122),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][5] ),
    .S(_07719_),
    .Z(_00459_));
 MUX2_X1 _13660_ (.A(net123),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][60] ),
    .S(_07719_),
    .Z(_00460_));
 MUX2_X1 _13661_ (.A(net124),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][61] ),
    .S(_07719_),
    .Z(_00461_));
 MUX2_X1 _13662_ (.A(net125),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][62] ),
    .S(_07719_),
    .Z(_00462_));
 MUX2_X1 _13663_ (.A(net126),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][63] ),
    .S(_07719_),
    .Z(_00463_));
 MUX2_X1 _13664_ (.A(net127),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][6] ),
    .S(_07713_),
    .Z(_00464_));
 MUX2_X1 _13665_ (.A(net128),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][7] ),
    .S(_07713_),
    .Z(_00465_));
 MUX2_X1 _13666_ (.A(net129),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][8] ),
    .S(_07713_),
    .Z(_00466_));
 MUX2_X1 _13667_ (.A(net130),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[0][9] ),
    .S(_07713_),
    .Z(_00467_));
 NAND2_X1 _13668_ (.A1(_10588_),
    .A2(_07711_),
    .ZN(_07720_));
 BUF_X4 _13669_ (.A(_07720_),
    .Z(_07721_));
 BUF_X4 _13670_ (.A(_07721_),
    .Z(_07722_));
 MUX2_X1 _13671_ (.A(net67),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][0] ),
    .S(_07722_),
    .Z(_00468_));
 MUX2_X1 _13672_ (.A(net68),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][10] ),
    .S(_07722_),
    .Z(_00469_));
 MUX2_X1 _13673_ (.A(net69),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][11] ),
    .S(_07722_),
    .Z(_00470_));
 MUX2_X1 _13674_ (.A(net70),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][12] ),
    .S(_07722_),
    .Z(_00471_));
 MUX2_X1 _13675_ (.A(net71),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][13] ),
    .S(_07722_),
    .Z(_00472_));
 MUX2_X1 _13676_ (.A(net72),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][14] ),
    .S(_07722_),
    .Z(_00473_));
 MUX2_X1 _13677_ (.A(net73),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][15] ),
    .S(_07722_),
    .Z(_00474_));
 MUX2_X1 _13678_ (.A(net74),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][16] ),
    .S(_07722_),
    .Z(_00475_));
 MUX2_X1 _13679_ (.A(net75),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][17] ),
    .S(_07722_),
    .Z(_00476_));
 MUX2_X1 _13680_ (.A(net76),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][18] ),
    .S(_07722_),
    .Z(_00477_));
 BUF_X4 _13681_ (.A(_07721_),
    .Z(_07723_));
 MUX2_X1 _13682_ (.A(net77),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][19] ),
    .S(_07723_),
    .Z(_00478_));
 MUX2_X1 _13683_ (.A(net78),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][1] ),
    .S(_07723_),
    .Z(_00479_));
 MUX2_X1 _13684_ (.A(net79),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][20] ),
    .S(_07723_),
    .Z(_00480_));
 MUX2_X1 _13685_ (.A(net80),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][21] ),
    .S(_07723_),
    .Z(_00481_));
 MUX2_X1 _13686_ (.A(net81),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][22] ),
    .S(_07723_),
    .Z(_00482_));
 MUX2_X1 _13687_ (.A(net82),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][23] ),
    .S(_07723_),
    .Z(_00483_));
 MUX2_X1 _13688_ (.A(net83),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][24] ),
    .S(_07723_),
    .Z(_00484_));
 MUX2_X1 _13689_ (.A(net84),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][25] ),
    .S(_07723_),
    .Z(_00485_));
 MUX2_X1 _13690_ (.A(net85),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][26] ),
    .S(_07723_),
    .Z(_00486_));
 MUX2_X1 _13691_ (.A(net86),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][27] ),
    .S(_07723_),
    .Z(_00487_));
 BUF_X4 _13692_ (.A(_07721_),
    .Z(_07724_));
 MUX2_X1 _13693_ (.A(net87),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][28] ),
    .S(_07724_),
    .Z(_00488_));
 MUX2_X1 _13694_ (.A(net88),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][29] ),
    .S(_07724_),
    .Z(_00489_));
 MUX2_X1 _13695_ (.A(net89),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][2] ),
    .S(_07724_),
    .Z(_00490_));
 MUX2_X1 _13696_ (.A(net90),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][30] ),
    .S(_07724_),
    .Z(_00491_));
 MUX2_X1 _13697_ (.A(net91),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][31] ),
    .S(_07724_),
    .Z(_00492_));
 MUX2_X1 _13698_ (.A(net92),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][32] ),
    .S(_07724_),
    .Z(_00493_));
 MUX2_X1 _13699_ (.A(net93),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][33] ),
    .S(_07724_),
    .Z(_00494_));
 MUX2_X1 _13700_ (.A(net94),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][34] ),
    .S(_07724_),
    .Z(_00495_));
 MUX2_X1 _13701_ (.A(net95),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][35] ),
    .S(_07724_),
    .Z(_00496_));
 MUX2_X1 _13702_ (.A(net96),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][36] ),
    .S(_07724_),
    .Z(_00497_));
 BUF_X4 _13703_ (.A(_07721_),
    .Z(_07725_));
 MUX2_X1 _13704_ (.A(net97),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][37] ),
    .S(_07725_),
    .Z(_00498_));
 MUX2_X1 _13705_ (.A(net98),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][38] ),
    .S(_07725_),
    .Z(_00499_));
 MUX2_X1 _13706_ (.A(net99),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][39] ),
    .S(_07725_),
    .Z(_00500_));
 MUX2_X1 _13707_ (.A(net100),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][3] ),
    .S(_07725_),
    .Z(_00501_));
 MUX2_X1 _13708_ (.A(net101),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][40] ),
    .S(_07725_),
    .Z(_00502_));
 MUX2_X1 _13709_ (.A(net102),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][41] ),
    .S(_07725_),
    .Z(_00503_));
 MUX2_X1 _13710_ (.A(net103),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][42] ),
    .S(_07725_),
    .Z(_00504_));
 MUX2_X1 _13711_ (.A(net104),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][43] ),
    .S(_07725_),
    .Z(_00505_));
 MUX2_X1 _13712_ (.A(net105),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][44] ),
    .S(_07725_),
    .Z(_00506_));
 MUX2_X1 _13713_ (.A(net106),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][45] ),
    .S(_07725_),
    .Z(_00507_));
 CLKBUF_X3 _13714_ (.A(_07721_),
    .Z(_07726_));
 MUX2_X1 _13715_ (.A(net107),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][46] ),
    .S(_07726_),
    .Z(_00508_));
 MUX2_X1 _13716_ (.A(net108),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][47] ),
    .S(_07726_),
    .Z(_00509_));
 MUX2_X1 _13717_ (.A(net109),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][48] ),
    .S(_07726_),
    .Z(_00510_));
 MUX2_X1 _13718_ (.A(net110),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][49] ),
    .S(_07726_),
    .Z(_00511_));
 MUX2_X1 _13719_ (.A(net111),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][4] ),
    .S(_07726_),
    .Z(_00512_));
 MUX2_X1 _13720_ (.A(net112),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][50] ),
    .S(_07726_),
    .Z(_00513_));
 MUX2_X1 _13721_ (.A(net113),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][51] ),
    .S(_07726_),
    .Z(_00514_));
 MUX2_X1 _13722_ (.A(net114),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][52] ),
    .S(_07726_),
    .Z(_00515_));
 MUX2_X1 _13723_ (.A(net115),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][53] ),
    .S(_07726_),
    .Z(_00516_));
 MUX2_X1 _13724_ (.A(net116),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][54] ),
    .S(_07726_),
    .Z(_00517_));
 BUF_X4 _13725_ (.A(_07721_),
    .Z(_07727_));
 MUX2_X1 _13726_ (.A(net117),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][55] ),
    .S(_07727_),
    .Z(_00518_));
 MUX2_X1 _13727_ (.A(net118),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][56] ),
    .S(_07727_),
    .Z(_00519_));
 MUX2_X1 _13728_ (.A(net119),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][57] ),
    .S(_07727_),
    .Z(_00520_));
 MUX2_X1 _13729_ (.A(net120),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][58] ),
    .S(_07727_),
    .Z(_00521_));
 MUX2_X1 _13730_ (.A(net121),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][59] ),
    .S(_07727_),
    .Z(_00522_));
 MUX2_X1 _13731_ (.A(net122),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][5] ),
    .S(_07727_),
    .Z(_00523_));
 MUX2_X1 _13732_ (.A(net123),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][60] ),
    .S(_07727_),
    .Z(_00524_));
 MUX2_X1 _13733_ (.A(net124),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][61] ),
    .S(_07727_),
    .Z(_00525_));
 MUX2_X1 _13734_ (.A(net125),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][62] ),
    .S(_07727_),
    .Z(_00526_));
 MUX2_X1 _13735_ (.A(net126),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][63] ),
    .S(_07727_),
    .Z(_00527_));
 MUX2_X1 _13736_ (.A(net127),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][6] ),
    .S(_07721_),
    .Z(_00528_));
 MUX2_X1 _13737_ (.A(net128),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][7] ),
    .S(_07721_),
    .Z(_00529_));
 MUX2_X1 _13738_ (.A(net129),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][8] ),
    .S(_07721_),
    .Z(_00530_));
 MUX2_X1 _13739_ (.A(net130),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[1][9] ),
    .S(_07721_),
    .Z(_00531_));
 NAND2_X1 _13740_ (.A1(_10586_),
    .A2(_07711_),
    .ZN(_07728_));
 BUF_X4 _13741_ (.A(_07728_),
    .Z(_07729_));
 BUF_X4 _13742_ (.A(_07729_),
    .Z(_07730_));
 MUX2_X1 _13743_ (.A(net67),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][0] ),
    .S(_07730_),
    .Z(_00532_));
 MUX2_X1 _13744_ (.A(net68),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][10] ),
    .S(_07730_),
    .Z(_00533_));
 MUX2_X1 _13745_ (.A(net69),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][11] ),
    .S(_07730_),
    .Z(_00534_));
 MUX2_X1 _13746_ (.A(net70),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][12] ),
    .S(_07730_),
    .Z(_00535_));
 MUX2_X1 _13747_ (.A(net71),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][13] ),
    .S(_07730_),
    .Z(_00536_));
 MUX2_X1 _13748_ (.A(net72),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][14] ),
    .S(_07730_),
    .Z(_00537_));
 MUX2_X1 _13749_ (.A(net73),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][15] ),
    .S(_07730_),
    .Z(_00538_));
 MUX2_X1 _13750_ (.A(net74),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][16] ),
    .S(_07730_),
    .Z(_00539_));
 MUX2_X1 _13751_ (.A(net75),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][17] ),
    .S(_07730_),
    .Z(_00540_));
 MUX2_X1 _13752_ (.A(net76),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][18] ),
    .S(_07730_),
    .Z(_00541_));
 BUF_X4 _13753_ (.A(_07729_),
    .Z(_07731_));
 MUX2_X1 _13754_ (.A(net77),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][19] ),
    .S(_07731_),
    .Z(_00542_));
 MUX2_X1 _13755_ (.A(net78),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][1] ),
    .S(_07731_),
    .Z(_00543_));
 MUX2_X1 _13756_ (.A(net79),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][20] ),
    .S(_07731_),
    .Z(_00544_));
 MUX2_X1 _13757_ (.A(net80),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][21] ),
    .S(_07731_),
    .Z(_00545_));
 MUX2_X1 _13758_ (.A(net81),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][22] ),
    .S(_07731_),
    .Z(_00546_));
 MUX2_X1 _13759_ (.A(net82),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][23] ),
    .S(_07731_),
    .Z(_00547_));
 MUX2_X1 _13760_ (.A(net83),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][24] ),
    .S(_07731_),
    .Z(_00548_));
 MUX2_X1 _13761_ (.A(net84),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][25] ),
    .S(_07731_),
    .Z(_00549_));
 MUX2_X1 _13762_ (.A(net85),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][26] ),
    .S(_07731_),
    .Z(_00550_));
 MUX2_X1 _13763_ (.A(net86),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][27] ),
    .S(_07731_),
    .Z(_00551_));
 BUF_X4 _13764_ (.A(_07729_),
    .Z(_07732_));
 MUX2_X1 _13765_ (.A(net87),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][28] ),
    .S(_07732_),
    .Z(_00552_));
 MUX2_X1 _13766_ (.A(net88),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][29] ),
    .S(_07732_),
    .Z(_00553_));
 MUX2_X1 _13767_ (.A(net89),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][2] ),
    .S(_07732_),
    .Z(_00554_));
 MUX2_X1 _13768_ (.A(net90),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][30] ),
    .S(_07732_),
    .Z(_00555_));
 MUX2_X1 _13769_ (.A(net91),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][31] ),
    .S(_07732_),
    .Z(_00556_));
 MUX2_X1 _13770_ (.A(net92),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][32] ),
    .S(_07732_),
    .Z(_00557_));
 MUX2_X1 _13771_ (.A(net93),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][33] ),
    .S(_07732_),
    .Z(_00558_));
 MUX2_X1 _13772_ (.A(net94),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][34] ),
    .S(_07732_),
    .Z(_00559_));
 MUX2_X1 _13773_ (.A(net95),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][35] ),
    .S(_07732_),
    .Z(_00560_));
 MUX2_X1 _13774_ (.A(net96),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][36] ),
    .S(_07732_),
    .Z(_00561_));
 BUF_X4 _13775_ (.A(_07729_),
    .Z(_07733_));
 MUX2_X1 _13776_ (.A(net97),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][37] ),
    .S(_07733_),
    .Z(_00562_));
 MUX2_X1 _13777_ (.A(net98),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][38] ),
    .S(_07733_),
    .Z(_00563_));
 MUX2_X1 _13778_ (.A(net99),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][39] ),
    .S(_07733_),
    .Z(_00564_));
 MUX2_X1 _13779_ (.A(net100),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][3] ),
    .S(_07733_),
    .Z(_00565_));
 MUX2_X1 _13780_ (.A(net101),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][40] ),
    .S(_07733_),
    .Z(_00566_));
 MUX2_X1 _13781_ (.A(net102),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][41] ),
    .S(_07733_),
    .Z(_00567_));
 MUX2_X1 _13782_ (.A(net103),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][42] ),
    .S(_07733_),
    .Z(_00568_));
 MUX2_X1 _13783_ (.A(net104),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][43] ),
    .S(_07733_),
    .Z(_00569_));
 MUX2_X1 _13784_ (.A(net105),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][44] ),
    .S(_07733_),
    .Z(_00570_));
 MUX2_X1 _13785_ (.A(net106),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][45] ),
    .S(_07733_),
    .Z(_00571_));
 BUF_X4 _13786_ (.A(_07729_),
    .Z(_07734_));
 MUX2_X1 _13787_ (.A(net107),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][46] ),
    .S(_07734_),
    .Z(_00572_));
 MUX2_X1 _13788_ (.A(net108),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][47] ),
    .S(_07734_),
    .Z(_00573_));
 MUX2_X1 _13789_ (.A(net109),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][48] ),
    .S(_07734_),
    .Z(_00574_));
 MUX2_X1 _13790_ (.A(net110),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][49] ),
    .S(_07734_),
    .Z(_00575_));
 MUX2_X1 _13791_ (.A(net111),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][4] ),
    .S(_07734_),
    .Z(_00576_));
 MUX2_X1 _13792_ (.A(net112),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][50] ),
    .S(_07734_),
    .Z(_00577_));
 MUX2_X1 _13793_ (.A(net113),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][51] ),
    .S(_07734_),
    .Z(_00578_));
 MUX2_X1 _13794_ (.A(net114),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][52] ),
    .S(_07734_),
    .Z(_00579_));
 MUX2_X1 _13795_ (.A(net115),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][53] ),
    .S(_07734_),
    .Z(_00580_));
 MUX2_X1 _13796_ (.A(net116),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][54] ),
    .S(_07734_),
    .Z(_00581_));
 BUF_X4 _13797_ (.A(_07729_),
    .Z(_07735_));
 MUX2_X1 _13798_ (.A(net117),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][55] ),
    .S(_07735_),
    .Z(_00582_));
 MUX2_X1 _13799_ (.A(net118),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][56] ),
    .S(_07735_),
    .Z(_00583_));
 MUX2_X1 _13800_ (.A(net119),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][57] ),
    .S(_07735_),
    .Z(_00584_));
 MUX2_X1 _13801_ (.A(net120),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][58] ),
    .S(_07735_),
    .Z(_00585_));
 MUX2_X1 _13802_ (.A(net121),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][59] ),
    .S(_07735_),
    .Z(_00586_));
 MUX2_X1 _13803_ (.A(net122),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][5] ),
    .S(_07735_),
    .Z(_00587_));
 MUX2_X1 _13804_ (.A(net123),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][60] ),
    .S(_07735_),
    .Z(_00588_));
 MUX2_X1 _13805_ (.A(net124),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][61] ),
    .S(_07735_),
    .Z(_00589_));
 MUX2_X1 _13806_ (.A(net125),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][62] ),
    .S(_07735_),
    .Z(_00590_));
 MUX2_X1 _13807_ (.A(net126),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][63] ),
    .S(_07735_),
    .Z(_00591_));
 MUX2_X1 _13808_ (.A(net127),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][6] ),
    .S(_07729_),
    .Z(_00592_));
 MUX2_X1 _13809_ (.A(net128),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][7] ),
    .S(_07729_),
    .Z(_00593_));
 MUX2_X1 _13810_ (.A(net129),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][8] ),
    .S(_07729_),
    .Z(_00594_));
 MUX2_X1 _13811_ (.A(net130),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][9] ),
    .S(_07729_),
    .Z(_00595_));
 NAND2_X1 _13812_ (.A1(_10590_),
    .A2(_07711_),
    .ZN(_07736_));
 BUF_X4 _13813_ (.A(_07736_),
    .Z(_07737_));
 BUF_X4 _13814_ (.A(_07737_),
    .Z(_07738_));
 MUX2_X1 _13815_ (.A(net67),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][0] ),
    .S(_07738_),
    .Z(_00596_));
 MUX2_X1 _13816_ (.A(net68),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][10] ),
    .S(_07738_),
    .Z(_00597_));
 MUX2_X1 _13817_ (.A(net69),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][11] ),
    .S(_07738_),
    .Z(_00598_));
 MUX2_X1 _13818_ (.A(net70),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][12] ),
    .S(_07738_),
    .Z(_00599_));
 MUX2_X1 _13819_ (.A(net71),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][13] ),
    .S(_07738_),
    .Z(_00600_));
 MUX2_X1 _13820_ (.A(net72),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][14] ),
    .S(_07738_),
    .Z(_00601_));
 MUX2_X1 _13821_ (.A(net73),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][15] ),
    .S(_07738_),
    .Z(_00602_));
 MUX2_X1 _13822_ (.A(net74),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][16] ),
    .S(_07738_),
    .Z(_00603_));
 MUX2_X1 _13823_ (.A(net75),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][17] ),
    .S(_07738_),
    .Z(_00604_));
 MUX2_X1 _13824_ (.A(net76),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][18] ),
    .S(_07738_),
    .Z(_00605_));
 BUF_X4 _13825_ (.A(_07737_),
    .Z(_07739_));
 MUX2_X1 _13826_ (.A(net77),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][19] ),
    .S(_07739_),
    .Z(_00606_));
 MUX2_X1 _13827_ (.A(net78),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][1] ),
    .S(_07739_),
    .Z(_00607_));
 MUX2_X1 _13828_ (.A(net79),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][20] ),
    .S(_07739_),
    .Z(_00608_));
 MUX2_X1 _13829_ (.A(net80),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][21] ),
    .S(_07739_),
    .Z(_00609_));
 MUX2_X1 _13830_ (.A(net81),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][22] ),
    .S(_07739_),
    .Z(_00610_));
 MUX2_X1 _13831_ (.A(net82),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][23] ),
    .S(_07739_),
    .Z(_00611_));
 MUX2_X1 _13832_ (.A(net83),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][24] ),
    .S(_07739_),
    .Z(_00612_));
 MUX2_X1 _13833_ (.A(net84),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][25] ),
    .S(_07739_),
    .Z(_00613_));
 MUX2_X1 _13834_ (.A(net85),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][26] ),
    .S(_07739_),
    .Z(_00614_));
 MUX2_X1 _13835_ (.A(net86),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][27] ),
    .S(_07739_),
    .Z(_00615_));
 BUF_X4 _13836_ (.A(_07737_),
    .Z(_07740_));
 MUX2_X1 _13837_ (.A(net87),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][28] ),
    .S(_07740_),
    .Z(_00616_));
 MUX2_X1 _13838_ (.A(net88),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][29] ),
    .S(_07740_),
    .Z(_00617_));
 MUX2_X1 _13839_ (.A(net89),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][2] ),
    .S(_07740_),
    .Z(_00618_));
 MUX2_X1 _13840_ (.A(net90),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][30] ),
    .S(_07740_),
    .Z(_00619_));
 MUX2_X1 _13841_ (.A(net91),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][31] ),
    .S(_07740_),
    .Z(_00620_));
 MUX2_X1 _13842_ (.A(net92),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][32] ),
    .S(_07740_),
    .Z(_00621_));
 MUX2_X1 _13843_ (.A(net93),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][33] ),
    .S(_07740_),
    .Z(_00622_));
 MUX2_X1 _13844_ (.A(net94),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][34] ),
    .S(_07740_),
    .Z(_00623_));
 MUX2_X1 _13845_ (.A(net95),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][35] ),
    .S(_07740_),
    .Z(_00624_));
 MUX2_X1 _13846_ (.A(net96),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][36] ),
    .S(_07740_),
    .Z(_00625_));
 BUF_X4 _13847_ (.A(_07737_),
    .Z(_07741_));
 MUX2_X1 _13848_ (.A(net97),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][37] ),
    .S(_07741_),
    .Z(_00626_));
 MUX2_X1 _13849_ (.A(net98),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][38] ),
    .S(_07741_),
    .Z(_00627_));
 MUX2_X1 _13850_ (.A(net99),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][39] ),
    .S(_07741_),
    .Z(_00628_));
 MUX2_X1 _13851_ (.A(net100),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][3] ),
    .S(_07741_),
    .Z(_00629_));
 MUX2_X1 _13852_ (.A(net101),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][40] ),
    .S(_07741_),
    .Z(_00630_));
 MUX2_X1 _13853_ (.A(net102),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][41] ),
    .S(_07741_),
    .Z(_00631_));
 MUX2_X1 _13854_ (.A(net103),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][42] ),
    .S(_07741_),
    .Z(_00632_));
 MUX2_X1 _13855_ (.A(net104),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][43] ),
    .S(_07741_),
    .Z(_00633_));
 MUX2_X1 _13856_ (.A(net105),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][44] ),
    .S(_07741_),
    .Z(_00634_));
 MUX2_X1 _13857_ (.A(net106),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][45] ),
    .S(_07741_),
    .Z(_00635_));
 BUF_X4 _13858_ (.A(_07737_),
    .Z(_07742_));
 MUX2_X1 _13859_ (.A(net107),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][46] ),
    .S(_07742_),
    .Z(_00636_));
 MUX2_X1 _13860_ (.A(net108),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][47] ),
    .S(_07742_),
    .Z(_00637_));
 MUX2_X1 _13861_ (.A(net109),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][48] ),
    .S(_07742_),
    .Z(_00638_));
 MUX2_X1 _13862_ (.A(net110),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][49] ),
    .S(_07742_),
    .Z(_00639_));
 MUX2_X1 _13863_ (.A(net111),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][4] ),
    .S(_07742_),
    .Z(_00640_));
 MUX2_X1 _13864_ (.A(net112),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][50] ),
    .S(_07742_),
    .Z(_00641_));
 MUX2_X1 _13865_ (.A(net113),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][51] ),
    .S(_07742_),
    .Z(_00642_));
 MUX2_X1 _13866_ (.A(net114),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][52] ),
    .S(_07742_),
    .Z(_00643_));
 MUX2_X1 _13867_ (.A(net115),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][53] ),
    .S(_07742_),
    .Z(_00644_));
 MUX2_X1 _13868_ (.A(net116),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][54] ),
    .S(_07742_),
    .Z(_00645_));
 BUF_X4 _13869_ (.A(_07737_),
    .Z(_07743_));
 MUX2_X1 _13870_ (.A(net117),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][55] ),
    .S(_07743_),
    .Z(_00646_));
 MUX2_X1 _13871_ (.A(net118),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][56] ),
    .S(_07743_),
    .Z(_00647_));
 MUX2_X1 _13872_ (.A(net119),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][57] ),
    .S(_07743_),
    .Z(_00648_));
 MUX2_X1 _13873_ (.A(net120),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][58] ),
    .S(_07743_),
    .Z(_00649_));
 MUX2_X1 _13874_ (.A(net121),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][59] ),
    .S(_07743_),
    .Z(_00650_));
 MUX2_X1 _13875_ (.A(net122),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][5] ),
    .S(_07743_),
    .Z(_00651_));
 MUX2_X1 _13876_ (.A(net123),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][60] ),
    .S(_07743_),
    .Z(_00652_));
 MUX2_X1 _13877_ (.A(net124),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][61] ),
    .S(_07743_),
    .Z(_00653_));
 MUX2_X1 _13878_ (.A(net125),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][62] ),
    .S(_07743_),
    .Z(_00654_));
 MUX2_X1 _13879_ (.A(net126),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][63] ),
    .S(_07743_),
    .Z(_00655_));
 MUX2_X1 _13880_ (.A(net127),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][6] ),
    .S(_07737_),
    .Z(_00656_));
 MUX2_X1 _13881_ (.A(net128),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][7] ),
    .S(_07737_),
    .Z(_00657_));
 MUX2_X1 _13882_ (.A(net129),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][8] ),
    .S(_07737_),
    .Z(_00658_));
 MUX2_X1 _13883_ (.A(net130),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][9] ),
    .S(_07737_),
    .Z(_00659_));
 BUF_X1 _13884_ (.A(dataIn_P[0]),
    .Z(_07744_));
 BUF_X2 _13885_ (.A(_07744_),
    .Z(_07745_));
 BUF_X2 _13886_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_f[3] ),
    .Z(_07746_));
 BUF_X2 _13887_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_f[2] ),
    .Z(_07747_));
 NAND2_X1 _13888_ (.A1(_10594_),
    .A2(_07677_),
    .ZN(_07748_));
 NOR4_X2 _13889_ (.A1(_06540_),
    .A2(_07746_),
    .A3(_07747_),
    .A4(_07748_),
    .ZN(_07749_));
 BUF_X4 _13890_ (.A(_07749_),
    .Z(_07750_));
 CLKBUF_X3 _13891_ (.A(_07750_),
    .Z(_07751_));
 MUX2_X1 _13892_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][0] ),
    .B(_07745_),
    .S(_07751_),
    .Z(_00687_));
 CLKBUF_X2 _13893_ (.A(dataIn_P[10]),
    .Z(_07752_));
 BUF_X2 _13894_ (.A(_07752_),
    .Z(_07753_));
 MUX2_X1 _13895_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][10] ),
    .B(_07753_),
    .S(_07751_),
    .Z(_00688_));
 CLKBUF_X2 _13896_ (.A(dataIn_P[11]),
    .Z(_07754_));
 BUF_X2 _13897_ (.A(_07754_),
    .Z(_07755_));
 MUX2_X1 _13898_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][11] ),
    .B(_07755_),
    .S(_07751_),
    .Z(_00689_));
 CLKBUF_X2 _13899_ (.A(dataIn_P[12]),
    .Z(_07756_));
 BUF_X2 _13900_ (.A(_07756_),
    .Z(_07757_));
 MUX2_X1 _13901_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][12] ),
    .B(_07757_),
    .S(_07751_),
    .Z(_00690_));
 CLKBUF_X2 _13902_ (.A(dataIn_P[13]),
    .Z(_07758_));
 BUF_X2 _13903_ (.A(_07758_),
    .Z(_07759_));
 MUX2_X1 _13904_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][13] ),
    .B(_07759_),
    .S(_07751_),
    .Z(_00691_));
 CLKBUF_X2 _13905_ (.A(dataIn_P[14]),
    .Z(_07760_));
 BUF_X2 _13906_ (.A(_07760_),
    .Z(_07761_));
 MUX2_X1 _13907_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][14] ),
    .B(_07761_),
    .S(_07751_),
    .Z(_00692_));
 CLKBUF_X2 _13908_ (.A(dataIn_P[15]),
    .Z(_07762_));
 BUF_X2 _13909_ (.A(_07762_),
    .Z(_07763_));
 MUX2_X1 _13910_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][15] ),
    .B(_07763_),
    .S(_07751_),
    .Z(_00693_));
 CLKBUF_X2 _13911_ (.A(dataIn_P[16]),
    .Z(_07764_));
 BUF_X2 _13912_ (.A(_07764_),
    .Z(_07765_));
 MUX2_X1 _13913_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][16] ),
    .B(_07765_),
    .S(_07751_),
    .Z(_00694_));
 CLKBUF_X2 _13914_ (.A(dataIn_P[17]),
    .Z(_07766_));
 BUF_X2 _13915_ (.A(_07766_),
    .Z(_07767_));
 MUX2_X1 _13916_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][17] ),
    .B(_07767_),
    .S(_07751_),
    .Z(_00695_));
 CLKBUF_X2 _13917_ (.A(dataIn_P[18]),
    .Z(_07768_));
 BUF_X2 _13918_ (.A(_07768_),
    .Z(_07769_));
 MUX2_X1 _13919_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][18] ),
    .B(_07769_),
    .S(_07751_),
    .Z(_00696_));
 BUF_X1 _13920_ (.A(dataIn_P[19]),
    .Z(_07770_));
 CLKBUF_X2 _13921_ (.A(_07770_),
    .Z(_07771_));
 BUF_X4 _13922_ (.A(_07750_),
    .Z(_07772_));
 MUX2_X1 _13923_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][19] ),
    .B(_07771_),
    .S(_07772_),
    .Z(_00697_));
 BUF_X1 _13924_ (.A(dataIn_P[1]),
    .Z(_07773_));
 CLKBUF_X2 _13925_ (.A(_07773_),
    .Z(_07774_));
 MUX2_X1 _13926_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][1] ),
    .B(_07774_),
    .S(_07772_),
    .Z(_00698_));
 BUF_X1 _13927_ (.A(dataIn_P[20]),
    .Z(_07775_));
 BUF_X2 _13928_ (.A(_07775_),
    .Z(_07776_));
 MUX2_X1 _13929_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][20] ),
    .B(_07776_),
    .S(_07772_),
    .Z(_00699_));
 CLKBUF_X2 _13930_ (.A(dataIn_P[21]),
    .Z(_07777_));
 BUF_X2 _13931_ (.A(_07777_),
    .Z(_07778_));
 MUX2_X1 _13932_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][21] ),
    .B(_07778_),
    .S(_07772_),
    .Z(_00700_));
 BUF_X1 _13933_ (.A(dataIn_P[22]),
    .Z(_07779_));
 BUF_X2 _13934_ (.A(_07779_),
    .Z(_07780_));
 MUX2_X1 _13935_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][22] ),
    .B(_07780_),
    .S(_07772_),
    .Z(_00701_));
 CLKBUF_X2 _13936_ (.A(dataIn_P[23]),
    .Z(_07781_));
 CLKBUF_X2 _13937_ (.A(_07781_),
    .Z(_07782_));
 MUX2_X1 _13938_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][23] ),
    .B(_07782_),
    .S(_07772_),
    .Z(_00702_));
 BUF_X1 _13939_ (.A(dataIn_P[24]),
    .Z(_07783_));
 CLKBUF_X2 _13940_ (.A(_07783_),
    .Z(_07784_));
 MUX2_X1 _13941_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][24] ),
    .B(_07784_),
    .S(_07772_),
    .Z(_00703_));
 BUF_X1 _13942_ (.A(dataIn_P[25]),
    .Z(_07785_));
 BUF_X2 _13943_ (.A(_07785_),
    .Z(_07786_));
 MUX2_X1 _13944_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][25] ),
    .B(_07786_),
    .S(_07772_),
    .Z(_00704_));
 BUF_X1 _13945_ (.A(dataIn_P[26]),
    .Z(_07787_));
 BUF_X2 _13946_ (.A(_07787_),
    .Z(_07788_));
 MUX2_X1 _13947_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][26] ),
    .B(_07788_),
    .S(_07772_),
    .Z(_00705_));
 BUF_X1 _13948_ (.A(dataIn_P[27]),
    .Z(_07789_));
 BUF_X2 _13949_ (.A(_07789_),
    .Z(_07790_));
 MUX2_X1 _13950_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][27] ),
    .B(_07790_),
    .S(_07772_),
    .Z(_00706_));
 BUF_X1 _13951_ (.A(dataIn_P[28]),
    .Z(_07791_));
 CLKBUF_X2 _13952_ (.A(_07791_),
    .Z(_07792_));
 BUF_X4 _13953_ (.A(_07750_),
    .Z(_07793_));
 MUX2_X1 _13954_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][28] ),
    .B(_07792_),
    .S(_07793_),
    .Z(_00707_));
 BUF_X1 _13955_ (.A(dataIn_P[29]),
    .Z(_07794_));
 BUF_X2 _13956_ (.A(_07794_),
    .Z(_07795_));
 MUX2_X1 _13957_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][29] ),
    .B(_07795_),
    .S(_07793_),
    .Z(_00708_));
 BUF_X1 _13958_ (.A(dataIn_P[2]),
    .Z(_07796_));
 BUF_X2 _13959_ (.A(_07796_),
    .Z(_07797_));
 MUX2_X1 _13960_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][2] ),
    .B(_07797_),
    .S(_07793_),
    .Z(_00709_));
 BUF_X1 _13961_ (.A(dataIn_P[30]),
    .Z(_07798_));
 CLKBUF_X2 _13962_ (.A(_07798_),
    .Z(_07799_));
 MUX2_X1 _13963_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][30] ),
    .B(_07799_),
    .S(_07793_),
    .Z(_00710_));
 BUF_X1 _13964_ (.A(dataIn_P[31]),
    .Z(_07800_));
 BUF_X2 _13965_ (.A(_07800_),
    .Z(_07801_));
 MUX2_X1 _13966_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][31] ),
    .B(_07801_),
    .S(_07793_),
    .Z(_00711_));
 BUF_X1 _13967_ (.A(dataIn_P[32]),
    .Z(_07802_));
 CLKBUF_X2 _13968_ (.A(_07802_),
    .Z(_07803_));
 MUX2_X1 _13969_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][32] ),
    .B(_07803_),
    .S(_07793_),
    .Z(_00712_));
 BUF_X1 _13970_ (.A(dataIn_P[33]),
    .Z(_07804_));
 CLKBUF_X2 _13971_ (.A(_07804_),
    .Z(_07805_));
 MUX2_X1 _13972_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][33] ),
    .B(_07805_),
    .S(_07793_),
    .Z(_00713_));
 BUF_X1 _13973_ (.A(dataIn_P[34]),
    .Z(_07806_));
 BUF_X2 _13974_ (.A(_07806_),
    .Z(_07807_));
 MUX2_X1 _13975_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][34] ),
    .B(_07807_),
    .S(_07793_),
    .Z(_00714_));
 CLKBUF_X2 _13976_ (.A(dataIn_P[35]),
    .Z(_07808_));
 BUF_X2 _13977_ (.A(_07808_),
    .Z(_07809_));
 MUX2_X1 _13978_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][35] ),
    .B(_07809_),
    .S(_07793_),
    .Z(_00715_));
 BUF_X1 _13979_ (.A(dataIn_P[36]),
    .Z(_07810_));
 BUF_X2 _13980_ (.A(_07810_),
    .Z(_07811_));
 MUX2_X1 _13981_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][36] ),
    .B(_07811_),
    .S(_07793_),
    .Z(_00716_));
 BUF_X1 _13982_ (.A(dataIn_P[37]),
    .Z(_07812_));
 BUF_X2 _13983_ (.A(_07812_),
    .Z(_07813_));
 BUF_X4 _13984_ (.A(_07750_),
    .Z(_07814_));
 MUX2_X1 _13985_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][37] ),
    .B(_07813_),
    .S(_07814_),
    .Z(_00717_));
 BUF_X1 _13986_ (.A(dataIn_P[38]),
    .Z(_07815_));
 BUF_X2 _13987_ (.A(_07815_),
    .Z(_07816_));
 MUX2_X1 _13988_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][38] ),
    .B(_07816_),
    .S(_07814_),
    .Z(_00718_));
 BUF_X1 _13989_ (.A(dataIn_P[39]),
    .Z(_07817_));
 BUF_X2 _13990_ (.A(_07817_),
    .Z(_07818_));
 MUX2_X1 _13991_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][39] ),
    .B(_07818_),
    .S(_07814_),
    .Z(_00719_));
 BUF_X1 _13992_ (.A(dataIn_P[3]),
    .Z(_07819_));
 CLKBUF_X2 _13993_ (.A(_07819_),
    .Z(_07820_));
 MUX2_X1 _13994_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][3] ),
    .B(_07820_),
    .S(_07814_),
    .Z(_00720_));
 BUF_X1 _13995_ (.A(dataIn_P[40]),
    .Z(_07821_));
 BUF_X2 _13996_ (.A(_07821_),
    .Z(_07822_));
 MUX2_X1 _13997_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][40] ),
    .B(_07822_),
    .S(_07814_),
    .Z(_00721_));
 CLKBUF_X2 _13998_ (.A(dataIn_P[41]),
    .Z(_07823_));
 BUF_X2 _13999_ (.A(_07823_),
    .Z(_07824_));
 MUX2_X1 _14000_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][41] ),
    .B(_07824_),
    .S(_07814_),
    .Z(_00722_));
 CLKBUF_X2 _14001_ (.A(dataIn_P[42]),
    .Z(_07825_));
 BUF_X2 _14002_ (.A(_07825_),
    .Z(_07826_));
 MUX2_X1 _14003_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][42] ),
    .B(_07826_),
    .S(_07814_),
    .Z(_00723_));
 BUF_X1 _14004_ (.A(dataIn_P[43]),
    .Z(_07827_));
 BUF_X2 _14005_ (.A(_07827_),
    .Z(_07828_));
 MUX2_X1 _14006_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][43] ),
    .B(_07828_),
    .S(_07814_),
    .Z(_00724_));
 BUF_X1 _14007_ (.A(dataIn_P[44]),
    .Z(_07829_));
 BUF_X2 _14008_ (.A(_07829_),
    .Z(_07830_));
 MUX2_X1 _14009_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][44] ),
    .B(_07830_),
    .S(_07814_),
    .Z(_00725_));
 BUF_X1 _14010_ (.A(dataIn_P[45]),
    .Z(_07831_));
 BUF_X2 _14011_ (.A(_07831_),
    .Z(_07832_));
 MUX2_X1 _14012_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][45] ),
    .B(_07832_),
    .S(_07814_),
    .Z(_00726_));
 BUF_X1 _14013_ (.A(dataIn_P[46]),
    .Z(_07833_));
 CLKBUF_X2 _14014_ (.A(_07833_),
    .Z(_07834_));
 BUF_X4 _14015_ (.A(_07750_),
    .Z(_07835_));
 MUX2_X1 _14016_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][46] ),
    .B(_07834_),
    .S(_07835_),
    .Z(_00727_));
 CLKBUF_X2 _14017_ (.A(dataIn_P[47]),
    .Z(_07836_));
 BUF_X2 _14018_ (.A(_07836_),
    .Z(_07837_));
 MUX2_X1 _14019_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][47] ),
    .B(_07837_),
    .S(_07835_),
    .Z(_00728_));
 BUF_X1 _14020_ (.A(dataIn_P[48]),
    .Z(_07838_));
 BUF_X2 _14021_ (.A(_07838_),
    .Z(_07839_));
 MUX2_X1 _14022_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][48] ),
    .B(_07839_),
    .S(_07835_),
    .Z(_00729_));
 BUF_X1 _14023_ (.A(dataIn_P[49]),
    .Z(_07840_));
 BUF_X2 _14024_ (.A(_07840_),
    .Z(_07841_));
 MUX2_X1 _14025_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][49] ),
    .B(_07841_),
    .S(_07835_),
    .Z(_00730_));
 BUF_X1 _14026_ (.A(dataIn_P[4]),
    .Z(_07842_));
 BUF_X2 _14027_ (.A(_07842_),
    .Z(_07843_));
 MUX2_X1 _14028_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][4] ),
    .B(_07843_),
    .S(_07835_),
    .Z(_00731_));
 CLKBUF_X2 _14029_ (.A(dataIn_P[50]),
    .Z(_07844_));
 BUF_X2 _14030_ (.A(_07844_),
    .Z(_07845_));
 MUX2_X1 _14031_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][50] ),
    .B(_07845_),
    .S(_07835_),
    .Z(_00732_));
 CLKBUF_X2 _14032_ (.A(dataIn_P[51]),
    .Z(_07846_));
 BUF_X2 _14033_ (.A(_07846_),
    .Z(_07847_));
 MUX2_X1 _14034_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][51] ),
    .B(_07847_),
    .S(_07835_),
    .Z(_00733_));
 CLKBUF_X2 _14035_ (.A(dataIn_P[52]),
    .Z(_07848_));
 BUF_X2 _14036_ (.A(_07848_),
    .Z(_07849_));
 MUX2_X1 _14037_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][52] ),
    .B(_07849_),
    .S(_07835_),
    .Z(_00734_));
 CLKBUF_X2 _14038_ (.A(dataIn_P[53]),
    .Z(_07850_));
 BUF_X2 _14039_ (.A(_07850_),
    .Z(_07851_));
 MUX2_X1 _14040_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][53] ),
    .B(_07851_),
    .S(_07835_),
    .Z(_00735_));
 BUF_X1 _14041_ (.A(dataIn_P[54]),
    .Z(_07852_));
 BUF_X2 _14042_ (.A(_07852_),
    .Z(_07853_));
 MUX2_X1 _14043_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][54] ),
    .B(_07853_),
    .S(_07835_),
    .Z(_00736_));
 BUF_X1 _14044_ (.A(dataIn_P[55]),
    .Z(_07854_));
 BUF_X2 _14045_ (.A(_07854_),
    .Z(_07855_));
 BUF_X4 _14046_ (.A(_07750_),
    .Z(_07856_));
 MUX2_X1 _14047_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][55] ),
    .B(_07855_),
    .S(_07856_),
    .Z(_00737_));
 BUF_X1 _14048_ (.A(dataIn_P[56]),
    .Z(_07857_));
 BUF_X2 _14049_ (.A(_07857_),
    .Z(_07858_));
 MUX2_X1 _14050_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][56] ),
    .B(_07858_),
    .S(_07856_),
    .Z(_00738_));
 BUF_X1 _14051_ (.A(dataIn_P[57]),
    .Z(_07859_));
 BUF_X2 _14052_ (.A(_07859_),
    .Z(_07860_));
 MUX2_X1 _14053_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][57] ),
    .B(_07860_),
    .S(_07856_),
    .Z(_00739_));
 CLKBUF_X2 _14054_ (.A(dataIn_P[58]),
    .Z(_07861_));
 BUF_X2 _14055_ (.A(_07861_),
    .Z(_07862_));
 MUX2_X1 _14056_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][58] ),
    .B(_07862_),
    .S(_07856_),
    .Z(_00740_));
 CLKBUF_X2 _14057_ (.A(dataIn_P[59]),
    .Z(_07863_));
 BUF_X2 _14058_ (.A(_07863_),
    .Z(_07864_));
 MUX2_X1 _14059_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][59] ),
    .B(_07864_),
    .S(_07856_),
    .Z(_00741_));
 BUF_X1 _14060_ (.A(dataIn_P[5]),
    .Z(_07865_));
 BUF_X2 _14061_ (.A(_07865_),
    .Z(_07866_));
 MUX2_X1 _14062_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][5] ),
    .B(_07866_),
    .S(_07856_),
    .Z(_00742_));
 CLKBUF_X2 _14063_ (.A(dataIn_P[60]),
    .Z(_07867_));
 BUF_X2 _14064_ (.A(_07867_),
    .Z(_07868_));
 MUX2_X1 _14065_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][60] ),
    .B(_07868_),
    .S(_07856_),
    .Z(_00743_));
 BUF_X1 _14066_ (.A(dataIn_P[61]),
    .Z(_07869_));
 BUF_X2 _14067_ (.A(_07869_),
    .Z(_07870_));
 MUX2_X1 _14068_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][61] ),
    .B(_07870_),
    .S(_07856_),
    .Z(_00744_));
 BUF_X1 _14069_ (.A(dataIn_P[62]),
    .Z(_07871_));
 BUF_X2 _14070_ (.A(_07871_),
    .Z(_07872_));
 MUX2_X1 _14071_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][62] ),
    .B(_07872_),
    .S(_07856_),
    .Z(_00745_));
 BUF_X1 _14072_ (.A(dataIn_P[63]),
    .Z(_07873_));
 BUF_X2 _14073_ (.A(_07873_),
    .Z(_07874_));
 MUX2_X1 _14074_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][63] ),
    .B(_07874_),
    .S(_07856_),
    .Z(_00746_));
 BUF_X1 _14075_ (.A(dataIn_P[6]),
    .Z(_07875_));
 BUF_X2 _14076_ (.A(_07875_),
    .Z(_07876_));
 MUX2_X1 _14077_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][6] ),
    .B(_07876_),
    .S(_07750_),
    .Z(_00747_));
 BUF_X1 _14078_ (.A(dataIn_P[7]),
    .Z(_07877_));
 BUF_X2 _14079_ (.A(_07877_),
    .Z(_07878_));
 MUX2_X1 _14080_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][7] ),
    .B(_07878_),
    .S(_07750_),
    .Z(_00748_));
 BUF_X1 _14081_ (.A(dataIn_P[8]),
    .Z(_07879_));
 BUF_X2 _14082_ (.A(_07879_),
    .Z(_07880_));
 MUX2_X1 _14083_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][8] ),
    .B(_07880_),
    .S(_07750_),
    .Z(_00749_));
 CLKBUF_X2 _14084_ (.A(dataIn_P[9]),
    .Z(_07881_));
 BUF_X2 _14085_ (.A(_07881_),
    .Z(_07882_));
 MUX2_X1 _14086_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][9] ),
    .B(_07882_),
    .S(_07750_),
    .Z(_00750_));
 INV_X1 _14087_ (.A(_07747_),
    .ZN(_07883_));
 NAND2_X1 _14088_ (.A1(_07883_),
    .A2(_07677_),
    .ZN(_07884_));
 NAND2_X1 _14089_ (.A1(_06581_),
    .A2(_07746_),
    .ZN(_07885_));
 NOR2_X1 _14090_ (.A1(_07884_),
    .A2(_07885_),
    .ZN(_07886_));
 NAND2_X1 _14091_ (.A1(_10595_),
    .A2(_07886_),
    .ZN(_07887_));
 BUF_X4 _14092_ (.A(_07887_),
    .Z(_07888_));
 CLKBUF_X3 _14093_ (.A(_07888_),
    .Z(_07889_));
 MUX2_X1 _14094_ (.A(_07745_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][0] ),
    .S(_07889_),
    .Z(_00751_));
 MUX2_X1 _14095_ (.A(_07753_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][10] ),
    .S(_07889_),
    .Z(_00752_));
 MUX2_X1 _14096_ (.A(_07755_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][11] ),
    .S(_07889_),
    .Z(_00753_));
 MUX2_X1 _14097_ (.A(_07757_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][12] ),
    .S(_07889_),
    .Z(_00754_));
 MUX2_X1 _14098_ (.A(_07759_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][13] ),
    .S(_07889_),
    .Z(_00755_));
 MUX2_X1 _14099_ (.A(_07761_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][14] ),
    .S(_07889_),
    .Z(_00756_));
 MUX2_X1 _14100_ (.A(_07763_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][15] ),
    .S(_07889_),
    .Z(_00757_));
 MUX2_X1 _14101_ (.A(_07765_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][16] ),
    .S(_07889_),
    .Z(_00758_));
 MUX2_X1 _14102_ (.A(_07767_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][17] ),
    .S(_07889_),
    .Z(_00759_));
 MUX2_X1 _14103_ (.A(_07769_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][18] ),
    .S(_07889_),
    .Z(_00760_));
 BUF_X4 _14104_ (.A(_07888_),
    .Z(_07890_));
 MUX2_X1 _14105_ (.A(_07771_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][19] ),
    .S(_07890_),
    .Z(_00761_));
 MUX2_X1 _14106_ (.A(_07774_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][1] ),
    .S(_07890_),
    .Z(_00762_));
 MUX2_X1 _14107_ (.A(_07776_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][20] ),
    .S(_07890_),
    .Z(_00763_));
 MUX2_X1 _14108_ (.A(_07778_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][21] ),
    .S(_07890_),
    .Z(_00764_));
 MUX2_X1 _14109_ (.A(_07780_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][22] ),
    .S(_07890_),
    .Z(_00765_));
 MUX2_X1 _14110_ (.A(_07782_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][23] ),
    .S(_07890_),
    .Z(_00766_));
 MUX2_X1 _14111_ (.A(_07784_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][24] ),
    .S(_07890_),
    .Z(_00767_));
 MUX2_X1 _14112_ (.A(_07786_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][25] ),
    .S(_07890_),
    .Z(_00768_));
 MUX2_X1 _14113_ (.A(_07788_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][26] ),
    .S(_07890_),
    .Z(_00769_));
 MUX2_X1 _14114_ (.A(_07790_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][27] ),
    .S(_07890_),
    .Z(_00770_));
 BUF_X4 _14115_ (.A(_07888_),
    .Z(_07891_));
 MUX2_X1 _14116_ (.A(_07792_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][28] ),
    .S(_07891_),
    .Z(_00771_));
 MUX2_X1 _14117_ (.A(_07795_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][29] ),
    .S(_07891_),
    .Z(_00772_));
 MUX2_X1 _14118_ (.A(_07797_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][2] ),
    .S(_07891_),
    .Z(_00773_));
 MUX2_X1 _14119_ (.A(_07799_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][30] ),
    .S(_07891_),
    .Z(_00774_));
 MUX2_X1 _14120_ (.A(_07801_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][31] ),
    .S(_07891_),
    .Z(_00775_));
 MUX2_X1 _14121_ (.A(_07803_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][32] ),
    .S(_07891_),
    .Z(_00776_));
 MUX2_X1 _14122_ (.A(_07805_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][33] ),
    .S(_07891_),
    .Z(_00777_));
 MUX2_X1 _14123_ (.A(_07807_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][34] ),
    .S(_07891_),
    .Z(_00778_));
 MUX2_X1 _14124_ (.A(_07809_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][35] ),
    .S(_07891_),
    .Z(_00779_));
 MUX2_X1 _14125_ (.A(_07811_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][36] ),
    .S(_07891_),
    .Z(_00780_));
 BUF_X4 _14126_ (.A(_07888_),
    .Z(_07892_));
 MUX2_X1 _14127_ (.A(_07813_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][37] ),
    .S(_07892_),
    .Z(_00781_));
 MUX2_X1 _14128_ (.A(_07816_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][38] ),
    .S(_07892_),
    .Z(_00782_));
 MUX2_X1 _14129_ (.A(_07818_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][39] ),
    .S(_07892_),
    .Z(_00783_));
 MUX2_X1 _14130_ (.A(_07820_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][3] ),
    .S(_07892_),
    .Z(_00784_));
 MUX2_X1 _14131_ (.A(_07822_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][40] ),
    .S(_07892_),
    .Z(_00785_));
 MUX2_X1 _14132_ (.A(_07824_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][41] ),
    .S(_07892_),
    .Z(_00786_));
 MUX2_X1 _14133_ (.A(_07826_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][42] ),
    .S(_07892_),
    .Z(_00787_));
 MUX2_X1 _14134_ (.A(_07828_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][43] ),
    .S(_07892_),
    .Z(_00788_));
 MUX2_X1 _14135_ (.A(_07830_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][44] ),
    .S(_07892_),
    .Z(_00789_));
 MUX2_X1 _14136_ (.A(_07832_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][45] ),
    .S(_07892_),
    .Z(_00790_));
 BUF_X4 _14137_ (.A(_07888_),
    .Z(_07893_));
 MUX2_X1 _14138_ (.A(_07834_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][46] ),
    .S(_07893_),
    .Z(_00791_));
 MUX2_X1 _14139_ (.A(_07837_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][47] ),
    .S(_07893_),
    .Z(_00792_));
 MUX2_X1 _14140_ (.A(_07839_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][48] ),
    .S(_07893_),
    .Z(_00793_));
 MUX2_X1 _14141_ (.A(_07841_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][49] ),
    .S(_07893_),
    .Z(_00794_));
 MUX2_X1 _14142_ (.A(_07843_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][4] ),
    .S(_07893_),
    .Z(_00795_));
 MUX2_X1 _14143_ (.A(_07845_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][50] ),
    .S(_07893_),
    .Z(_00796_));
 MUX2_X1 _14144_ (.A(_07847_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][51] ),
    .S(_07893_),
    .Z(_00797_));
 MUX2_X1 _14145_ (.A(_07849_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][52] ),
    .S(_07893_),
    .Z(_00798_));
 MUX2_X1 _14146_ (.A(_07851_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][53] ),
    .S(_07893_),
    .Z(_00799_));
 MUX2_X1 _14147_ (.A(_07853_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][54] ),
    .S(_07893_),
    .Z(_00800_));
 BUF_X4 _14148_ (.A(_07888_),
    .Z(_07894_));
 MUX2_X1 _14149_ (.A(_07855_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][55] ),
    .S(_07894_),
    .Z(_00801_));
 MUX2_X1 _14150_ (.A(_07858_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][56] ),
    .S(_07894_),
    .Z(_00802_));
 MUX2_X1 _14151_ (.A(_07860_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][57] ),
    .S(_07894_),
    .Z(_00803_));
 MUX2_X1 _14152_ (.A(_07862_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][58] ),
    .S(_07894_),
    .Z(_00804_));
 MUX2_X1 _14153_ (.A(_07864_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][59] ),
    .S(_07894_),
    .Z(_00805_));
 MUX2_X1 _14154_ (.A(_07866_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][5] ),
    .S(_07894_),
    .Z(_00806_));
 MUX2_X1 _14155_ (.A(_07868_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][60] ),
    .S(_07894_),
    .Z(_00807_));
 MUX2_X1 _14156_ (.A(_07870_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][61] ),
    .S(_07894_),
    .Z(_00808_));
 MUX2_X1 _14157_ (.A(_07872_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][62] ),
    .S(_07894_),
    .Z(_00809_));
 MUX2_X1 _14158_ (.A(_07874_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][63] ),
    .S(_07894_),
    .Z(_00810_));
 MUX2_X1 _14159_ (.A(_07876_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][6] ),
    .S(_07888_),
    .Z(_00811_));
 MUX2_X1 _14160_ (.A(_07878_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][7] ),
    .S(_07888_),
    .Z(_00812_));
 MUX2_X1 _14161_ (.A(_07880_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][8] ),
    .S(_07888_),
    .Z(_00813_));
 MUX2_X1 _14162_ (.A(_07882_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][9] ),
    .S(_07888_),
    .Z(_00814_));
 BUF_X1 _14163_ (.A(_10599_),
    .Z(_07895_));
 NAND2_X1 _14164_ (.A1(_07895_),
    .A2(_07886_),
    .ZN(_07896_));
 BUF_X4 _14165_ (.A(_07896_),
    .Z(_07897_));
 CLKBUF_X3 _14166_ (.A(_07897_),
    .Z(_07898_));
 MUX2_X1 _14167_ (.A(_07745_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][0] ),
    .S(_07898_),
    .Z(_00815_));
 MUX2_X1 _14168_ (.A(_07753_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][10] ),
    .S(_07898_),
    .Z(_00816_));
 MUX2_X1 _14169_ (.A(_07755_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][11] ),
    .S(_07898_),
    .Z(_00817_));
 MUX2_X1 _14170_ (.A(_07757_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][12] ),
    .S(_07898_),
    .Z(_00818_));
 MUX2_X1 _14171_ (.A(_07759_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][13] ),
    .S(_07898_),
    .Z(_00819_));
 MUX2_X1 _14172_ (.A(_07761_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][14] ),
    .S(_07898_),
    .Z(_00820_));
 MUX2_X1 _14173_ (.A(_07763_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][15] ),
    .S(_07898_),
    .Z(_00821_));
 MUX2_X1 _14174_ (.A(_07765_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][16] ),
    .S(_07898_),
    .Z(_00822_));
 MUX2_X1 _14175_ (.A(_07767_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][17] ),
    .S(_07898_),
    .Z(_00823_));
 MUX2_X1 _14176_ (.A(_07769_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][18] ),
    .S(_07898_),
    .Z(_00824_));
 BUF_X4 _14177_ (.A(_07897_),
    .Z(_07899_));
 MUX2_X1 _14178_ (.A(_07771_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][19] ),
    .S(_07899_),
    .Z(_00825_));
 MUX2_X1 _14179_ (.A(_07774_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][1] ),
    .S(_07899_),
    .Z(_00826_));
 MUX2_X1 _14180_ (.A(_07776_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][20] ),
    .S(_07899_),
    .Z(_00827_));
 MUX2_X1 _14181_ (.A(_07778_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][21] ),
    .S(_07899_),
    .Z(_00828_));
 MUX2_X1 _14182_ (.A(_07780_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][22] ),
    .S(_07899_),
    .Z(_00829_));
 MUX2_X1 _14183_ (.A(_07782_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][23] ),
    .S(_07899_),
    .Z(_00830_));
 MUX2_X1 _14184_ (.A(_07784_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][24] ),
    .S(_07899_),
    .Z(_00831_));
 MUX2_X1 _14185_ (.A(_07786_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][25] ),
    .S(_07899_),
    .Z(_00832_));
 MUX2_X1 _14186_ (.A(_07788_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][26] ),
    .S(_07899_),
    .Z(_00833_));
 MUX2_X1 _14187_ (.A(_07790_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][27] ),
    .S(_07899_),
    .Z(_00834_));
 BUF_X4 _14188_ (.A(_07897_),
    .Z(_07900_));
 MUX2_X1 _14189_ (.A(_07792_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][28] ),
    .S(_07900_),
    .Z(_00835_));
 MUX2_X1 _14190_ (.A(_07795_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][29] ),
    .S(_07900_),
    .Z(_00836_));
 MUX2_X1 _14191_ (.A(_07797_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][2] ),
    .S(_07900_),
    .Z(_00837_));
 MUX2_X1 _14192_ (.A(_07799_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][30] ),
    .S(_07900_),
    .Z(_00838_));
 MUX2_X1 _14193_ (.A(_07801_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][31] ),
    .S(_07900_),
    .Z(_00839_));
 MUX2_X1 _14194_ (.A(_07803_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][32] ),
    .S(_07900_),
    .Z(_00840_));
 MUX2_X1 _14195_ (.A(_07805_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][33] ),
    .S(_07900_),
    .Z(_00841_));
 MUX2_X1 _14196_ (.A(_07807_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][34] ),
    .S(_07900_),
    .Z(_00842_));
 MUX2_X1 _14197_ (.A(_07809_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][35] ),
    .S(_07900_),
    .Z(_00843_));
 MUX2_X1 _14198_ (.A(_07811_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][36] ),
    .S(_07900_),
    .Z(_00844_));
 BUF_X4 _14199_ (.A(_07897_),
    .Z(_07901_));
 MUX2_X1 _14200_ (.A(_07813_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][37] ),
    .S(_07901_),
    .Z(_00845_));
 MUX2_X1 _14201_ (.A(_07816_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][38] ),
    .S(_07901_),
    .Z(_00846_));
 MUX2_X1 _14202_ (.A(_07818_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][39] ),
    .S(_07901_),
    .Z(_00847_));
 MUX2_X1 _14203_ (.A(_07820_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][3] ),
    .S(_07901_),
    .Z(_00848_));
 MUX2_X1 _14204_ (.A(_07822_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][40] ),
    .S(_07901_),
    .Z(_00849_));
 MUX2_X1 _14205_ (.A(_07824_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][41] ),
    .S(_07901_),
    .Z(_00850_));
 MUX2_X1 _14206_ (.A(_07826_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][42] ),
    .S(_07901_),
    .Z(_00851_));
 MUX2_X1 _14207_ (.A(_07828_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][43] ),
    .S(_07901_),
    .Z(_00852_));
 MUX2_X1 _14208_ (.A(_07830_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][44] ),
    .S(_07901_),
    .Z(_00853_));
 MUX2_X1 _14209_ (.A(_07832_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][45] ),
    .S(_07901_),
    .Z(_00854_));
 BUF_X4 _14210_ (.A(_07897_),
    .Z(_07902_));
 MUX2_X1 _14211_ (.A(_07834_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][46] ),
    .S(_07902_),
    .Z(_00855_));
 MUX2_X1 _14212_ (.A(_07837_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][47] ),
    .S(_07902_),
    .Z(_00856_));
 MUX2_X1 _14213_ (.A(_07839_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][48] ),
    .S(_07902_),
    .Z(_00857_));
 MUX2_X1 _14214_ (.A(_07841_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][49] ),
    .S(_07902_),
    .Z(_00858_));
 MUX2_X1 _14215_ (.A(_07843_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][4] ),
    .S(_07902_),
    .Z(_00859_));
 MUX2_X1 _14216_ (.A(_07845_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][50] ),
    .S(_07902_),
    .Z(_00860_));
 MUX2_X1 _14217_ (.A(_07847_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][51] ),
    .S(_07902_),
    .Z(_00861_));
 MUX2_X1 _14218_ (.A(_07849_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][52] ),
    .S(_07902_),
    .Z(_00862_));
 MUX2_X1 _14219_ (.A(_07851_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][53] ),
    .S(_07902_),
    .Z(_00863_));
 MUX2_X1 _14220_ (.A(_07853_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][54] ),
    .S(_07902_),
    .Z(_00864_));
 BUF_X4 _14221_ (.A(_07897_),
    .Z(_07903_));
 MUX2_X1 _14222_ (.A(_07855_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][55] ),
    .S(_07903_),
    .Z(_00865_));
 MUX2_X1 _14223_ (.A(_07858_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][56] ),
    .S(_07903_),
    .Z(_00866_));
 MUX2_X1 _14224_ (.A(_07860_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][57] ),
    .S(_07903_),
    .Z(_00867_));
 MUX2_X1 _14225_ (.A(_07862_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][58] ),
    .S(_07903_),
    .Z(_00868_));
 MUX2_X1 _14226_ (.A(_07864_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][59] ),
    .S(_07903_),
    .Z(_00869_));
 MUX2_X1 _14227_ (.A(_07866_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][5] ),
    .S(_07903_),
    .Z(_00870_));
 MUX2_X1 _14228_ (.A(_07868_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][60] ),
    .S(_07903_),
    .Z(_00871_));
 MUX2_X1 _14229_ (.A(_07870_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][61] ),
    .S(_07903_),
    .Z(_00872_));
 MUX2_X1 _14230_ (.A(_07872_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][62] ),
    .S(_07903_),
    .Z(_00873_));
 MUX2_X1 _14231_ (.A(_07874_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][63] ),
    .S(_07903_),
    .Z(_00874_));
 MUX2_X1 _14232_ (.A(_07876_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][6] ),
    .S(_07897_),
    .Z(_00875_));
 MUX2_X1 _14233_ (.A(_07878_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][7] ),
    .S(_07897_),
    .Z(_00876_));
 MUX2_X1 _14234_ (.A(_07880_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][8] ),
    .S(_07897_),
    .Z(_00877_));
 MUX2_X1 _14235_ (.A(_07882_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][9] ),
    .S(_07897_),
    .Z(_00878_));
 NAND3_X1 _14236_ (.A1(_07747_),
    .A2(_10594_),
    .A3(_07677_),
    .ZN(_07904_));
 NOR2_X1 _14237_ (.A1(_07885_),
    .A2(_07904_),
    .ZN(_07905_));
 BUF_X4 _14238_ (.A(_07905_),
    .Z(_07906_));
 BUF_X4 _14239_ (.A(_07906_),
    .Z(_07907_));
 MUX2_X1 _14240_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][0] ),
    .B(_07745_),
    .S(_07907_),
    .Z(_00879_));
 MUX2_X1 _14241_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][10] ),
    .B(_07753_),
    .S(_07907_),
    .Z(_00880_));
 MUX2_X1 _14242_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][11] ),
    .B(_07755_),
    .S(_07907_),
    .Z(_00881_));
 MUX2_X1 _14243_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][12] ),
    .B(_07757_),
    .S(_07907_),
    .Z(_00882_));
 MUX2_X1 _14244_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][13] ),
    .B(_07759_),
    .S(_07907_),
    .Z(_00883_));
 MUX2_X1 _14245_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][14] ),
    .B(_07761_),
    .S(_07907_),
    .Z(_00884_));
 MUX2_X1 _14246_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][15] ),
    .B(_07763_),
    .S(_07907_),
    .Z(_00885_));
 MUX2_X1 _14247_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][16] ),
    .B(_07765_),
    .S(_07907_),
    .Z(_00886_));
 MUX2_X1 _14248_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][17] ),
    .B(_07767_),
    .S(_07907_),
    .Z(_00887_));
 MUX2_X1 _14249_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][18] ),
    .B(_07769_),
    .S(_07907_),
    .Z(_00888_));
 BUF_X4 _14250_ (.A(_07906_),
    .Z(_07908_));
 MUX2_X1 _14251_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][19] ),
    .B(_07771_),
    .S(_07908_),
    .Z(_00889_));
 MUX2_X1 _14252_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][1] ),
    .B(_07774_),
    .S(_07908_),
    .Z(_00890_));
 MUX2_X1 _14253_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][20] ),
    .B(_07776_),
    .S(_07908_),
    .Z(_00891_));
 MUX2_X1 _14254_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][21] ),
    .B(_07778_),
    .S(_07908_),
    .Z(_00892_));
 MUX2_X1 _14255_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][22] ),
    .B(_07780_),
    .S(_07908_),
    .Z(_00893_));
 MUX2_X1 _14256_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][23] ),
    .B(_07782_),
    .S(_07908_),
    .Z(_00894_));
 MUX2_X1 _14257_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][24] ),
    .B(_07784_),
    .S(_07908_),
    .Z(_00895_));
 MUX2_X1 _14258_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][25] ),
    .B(_07786_),
    .S(_07908_),
    .Z(_00896_));
 MUX2_X1 _14259_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][26] ),
    .B(_07788_),
    .S(_07908_),
    .Z(_00897_));
 MUX2_X1 _14260_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][27] ),
    .B(_07790_),
    .S(_07908_),
    .Z(_00898_));
 BUF_X4 _14261_ (.A(_07906_),
    .Z(_07909_));
 MUX2_X1 _14262_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][28] ),
    .B(_07792_),
    .S(_07909_),
    .Z(_00899_));
 MUX2_X1 _14263_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][29] ),
    .B(_07795_),
    .S(_07909_),
    .Z(_00900_));
 MUX2_X1 _14264_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][2] ),
    .B(_07797_),
    .S(_07909_),
    .Z(_00901_));
 MUX2_X1 _14265_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][30] ),
    .B(_07799_),
    .S(_07909_),
    .Z(_00902_));
 MUX2_X1 _14266_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][31] ),
    .B(_07801_),
    .S(_07909_),
    .Z(_00903_));
 MUX2_X1 _14267_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][32] ),
    .B(_07803_),
    .S(_07909_),
    .Z(_00904_));
 MUX2_X1 _14268_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][33] ),
    .B(_07805_),
    .S(_07909_),
    .Z(_00905_));
 MUX2_X1 _14269_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][34] ),
    .B(_07807_),
    .S(_07909_),
    .Z(_00906_));
 MUX2_X1 _14270_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][35] ),
    .B(_07809_),
    .S(_07909_),
    .Z(_00907_));
 MUX2_X1 _14271_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][36] ),
    .B(_07811_),
    .S(_07909_),
    .Z(_00908_));
 BUF_X4 _14272_ (.A(_07906_),
    .Z(_07910_));
 MUX2_X1 _14273_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][37] ),
    .B(_07813_),
    .S(_07910_),
    .Z(_00909_));
 MUX2_X1 _14274_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][38] ),
    .B(_07816_),
    .S(_07910_),
    .Z(_00910_));
 MUX2_X1 _14275_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][39] ),
    .B(_07818_),
    .S(_07910_),
    .Z(_00911_));
 MUX2_X1 _14276_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][3] ),
    .B(_07820_),
    .S(_07910_),
    .Z(_00912_));
 MUX2_X1 _14277_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][40] ),
    .B(_07822_),
    .S(_07910_),
    .Z(_00913_));
 MUX2_X1 _14278_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][41] ),
    .B(_07824_),
    .S(_07910_),
    .Z(_00914_));
 MUX2_X1 _14279_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][42] ),
    .B(_07826_),
    .S(_07910_),
    .Z(_00915_));
 MUX2_X1 _14280_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][43] ),
    .B(_07828_),
    .S(_07910_),
    .Z(_00916_));
 MUX2_X1 _14281_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][44] ),
    .B(_07830_),
    .S(_07910_),
    .Z(_00917_));
 MUX2_X1 _14282_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][45] ),
    .B(_07832_),
    .S(_07910_),
    .Z(_00918_));
 BUF_X4 _14283_ (.A(_07906_),
    .Z(_07911_));
 MUX2_X1 _14284_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][46] ),
    .B(_07834_),
    .S(_07911_),
    .Z(_00919_));
 MUX2_X1 _14285_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][47] ),
    .B(_07837_),
    .S(_07911_),
    .Z(_00920_));
 MUX2_X1 _14286_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][48] ),
    .B(_07839_),
    .S(_07911_),
    .Z(_00921_));
 MUX2_X1 _14287_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][49] ),
    .B(_07841_),
    .S(_07911_),
    .Z(_00922_));
 MUX2_X1 _14288_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][4] ),
    .B(_07843_),
    .S(_07911_),
    .Z(_00923_));
 MUX2_X1 _14289_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][50] ),
    .B(_07845_),
    .S(_07911_),
    .Z(_00924_));
 MUX2_X1 _14290_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][51] ),
    .B(_07847_),
    .S(_07911_),
    .Z(_00925_));
 MUX2_X1 _14291_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][52] ),
    .B(_07849_),
    .S(_07911_),
    .Z(_00926_));
 MUX2_X1 _14292_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][53] ),
    .B(_07851_),
    .S(_07911_),
    .Z(_00927_));
 MUX2_X1 _14293_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][54] ),
    .B(_07853_),
    .S(_07911_),
    .Z(_00928_));
 BUF_X4 _14294_ (.A(_07906_),
    .Z(_07912_));
 MUX2_X1 _14295_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][55] ),
    .B(_07855_),
    .S(_07912_),
    .Z(_00929_));
 MUX2_X1 _14296_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][56] ),
    .B(_07858_),
    .S(_07912_),
    .Z(_00930_));
 MUX2_X1 _14297_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][57] ),
    .B(_07860_),
    .S(_07912_),
    .Z(_00931_));
 MUX2_X1 _14298_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][58] ),
    .B(_07862_),
    .S(_07912_),
    .Z(_00932_));
 MUX2_X1 _14299_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][59] ),
    .B(_07864_),
    .S(_07912_),
    .Z(_00933_));
 MUX2_X1 _14300_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][5] ),
    .B(_07866_),
    .S(_07912_),
    .Z(_00934_));
 MUX2_X1 _14301_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][60] ),
    .B(_07868_),
    .S(_07912_),
    .Z(_00935_));
 MUX2_X1 _14302_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][61] ),
    .B(_07870_),
    .S(_07912_),
    .Z(_00936_));
 MUX2_X1 _14303_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][62] ),
    .B(_07872_),
    .S(_07912_),
    .Z(_00937_));
 MUX2_X1 _14304_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][63] ),
    .B(_07874_),
    .S(_07912_),
    .Z(_00938_));
 MUX2_X1 _14305_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][6] ),
    .B(_07876_),
    .S(_07906_),
    .Z(_00939_));
 MUX2_X1 _14306_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][7] ),
    .B(_07878_),
    .S(_07906_),
    .Z(_00940_));
 MUX2_X1 _14307_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][8] ),
    .B(_07880_),
    .S(_07906_),
    .Z(_00941_));
 MUX2_X1 _14308_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][9] ),
    .B(_07882_),
    .S(_07906_),
    .Z(_00942_));
 NAND2_X1 _14309_ (.A1(_07747_),
    .A2(_07677_),
    .ZN(_07913_));
 NOR2_X1 _14310_ (.A1(_07885_),
    .A2(_07913_),
    .ZN(_07914_));
 NAND2_X1 _14311_ (.A1(_10597_),
    .A2(_07914_),
    .ZN(_07915_));
 BUF_X4 _14312_ (.A(_07915_),
    .Z(_07916_));
 BUF_X4 _14313_ (.A(_07916_),
    .Z(_07917_));
 MUX2_X1 _14314_ (.A(_07745_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][0] ),
    .S(_07917_),
    .Z(_00943_));
 MUX2_X1 _14315_ (.A(_07753_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][10] ),
    .S(_07917_),
    .Z(_00944_));
 MUX2_X1 _14316_ (.A(_07755_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][11] ),
    .S(_07917_),
    .Z(_00945_));
 MUX2_X1 _14317_ (.A(_07757_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][12] ),
    .S(_07917_),
    .Z(_00946_));
 MUX2_X1 _14318_ (.A(_07759_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][13] ),
    .S(_07917_),
    .Z(_00947_));
 MUX2_X1 _14319_ (.A(_07761_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][14] ),
    .S(_07917_),
    .Z(_00948_));
 MUX2_X1 _14320_ (.A(_07763_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][15] ),
    .S(_07917_),
    .Z(_00949_));
 MUX2_X1 _14321_ (.A(_07765_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][16] ),
    .S(_07917_),
    .Z(_00950_));
 MUX2_X1 _14322_ (.A(_07767_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][17] ),
    .S(_07917_),
    .Z(_00951_));
 MUX2_X1 _14323_ (.A(_07769_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][18] ),
    .S(_07917_),
    .Z(_00952_));
 BUF_X4 _14324_ (.A(_07916_),
    .Z(_07918_));
 MUX2_X1 _14325_ (.A(_07771_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][19] ),
    .S(_07918_),
    .Z(_00953_));
 MUX2_X1 _14326_ (.A(_07774_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][1] ),
    .S(_07918_),
    .Z(_00954_));
 MUX2_X1 _14327_ (.A(_07776_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][20] ),
    .S(_07918_),
    .Z(_00955_));
 MUX2_X1 _14328_ (.A(_07778_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][21] ),
    .S(_07918_),
    .Z(_00956_));
 MUX2_X1 _14329_ (.A(_07780_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][22] ),
    .S(_07918_),
    .Z(_00957_));
 MUX2_X1 _14330_ (.A(_07782_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][23] ),
    .S(_07918_),
    .Z(_00958_));
 MUX2_X1 _14331_ (.A(_07784_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][24] ),
    .S(_07918_),
    .Z(_00959_));
 MUX2_X1 _14332_ (.A(_07786_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][25] ),
    .S(_07918_),
    .Z(_00960_));
 MUX2_X1 _14333_ (.A(_07788_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][26] ),
    .S(_07918_),
    .Z(_00961_));
 MUX2_X1 _14334_ (.A(_07790_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][27] ),
    .S(_07918_),
    .Z(_00962_));
 BUF_X4 _14335_ (.A(_07916_),
    .Z(_07919_));
 MUX2_X1 _14336_ (.A(_07792_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][28] ),
    .S(_07919_),
    .Z(_00963_));
 MUX2_X1 _14337_ (.A(_07795_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][29] ),
    .S(_07919_),
    .Z(_00964_));
 MUX2_X1 _14338_ (.A(_07797_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][2] ),
    .S(_07919_),
    .Z(_00965_));
 MUX2_X1 _14339_ (.A(_07799_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][30] ),
    .S(_07919_),
    .Z(_00966_));
 MUX2_X1 _14340_ (.A(_07801_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][31] ),
    .S(_07919_),
    .Z(_00967_));
 MUX2_X1 _14341_ (.A(_07803_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][32] ),
    .S(_07919_),
    .Z(_00968_));
 MUX2_X1 _14342_ (.A(_07805_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][33] ),
    .S(_07919_),
    .Z(_00969_));
 MUX2_X1 _14343_ (.A(_07807_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][34] ),
    .S(_07919_),
    .Z(_00970_));
 MUX2_X1 _14344_ (.A(_07809_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][35] ),
    .S(_07919_),
    .Z(_00971_));
 MUX2_X1 _14345_ (.A(_07811_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][36] ),
    .S(_07919_),
    .Z(_00972_));
 BUF_X4 _14346_ (.A(_07916_),
    .Z(_07920_));
 MUX2_X1 _14347_ (.A(_07813_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][37] ),
    .S(_07920_),
    .Z(_00973_));
 MUX2_X1 _14348_ (.A(_07816_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][38] ),
    .S(_07920_),
    .Z(_00974_));
 MUX2_X1 _14349_ (.A(_07818_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][39] ),
    .S(_07920_),
    .Z(_00975_));
 MUX2_X1 _14350_ (.A(_07820_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][3] ),
    .S(_07920_),
    .Z(_00976_));
 MUX2_X1 _14351_ (.A(_07822_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][40] ),
    .S(_07920_),
    .Z(_00977_));
 MUX2_X1 _14352_ (.A(_07824_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][41] ),
    .S(_07920_),
    .Z(_00978_));
 MUX2_X1 _14353_ (.A(_07826_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][42] ),
    .S(_07920_),
    .Z(_00979_));
 MUX2_X1 _14354_ (.A(_07828_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][43] ),
    .S(_07920_),
    .Z(_00980_));
 MUX2_X1 _14355_ (.A(_07830_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][44] ),
    .S(_07920_),
    .Z(_00981_));
 MUX2_X1 _14356_ (.A(_07832_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][45] ),
    .S(_07920_),
    .Z(_00982_));
 BUF_X4 _14357_ (.A(_07916_),
    .Z(_07921_));
 MUX2_X1 _14358_ (.A(_07834_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][46] ),
    .S(_07921_),
    .Z(_00983_));
 MUX2_X1 _14359_ (.A(_07837_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][47] ),
    .S(_07921_),
    .Z(_00984_));
 MUX2_X1 _14360_ (.A(_07839_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][48] ),
    .S(_07921_),
    .Z(_00985_));
 MUX2_X1 _14361_ (.A(_07841_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][49] ),
    .S(_07921_),
    .Z(_00986_));
 MUX2_X1 _14362_ (.A(_07843_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][4] ),
    .S(_07921_),
    .Z(_00987_));
 MUX2_X1 _14363_ (.A(_07845_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][50] ),
    .S(_07921_),
    .Z(_00988_));
 MUX2_X1 _14364_ (.A(_07847_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][51] ),
    .S(_07921_),
    .Z(_00989_));
 MUX2_X1 _14365_ (.A(_07849_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][52] ),
    .S(_07921_),
    .Z(_00990_));
 MUX2_X1 _14366_ (.A(_07851_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][53] ),
    .S(_07921_),
    .Z(_00991_));
 MUX2_X1 _14367_ (.A(_07853_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][54] ),
    .S(_07921_),
    .Z(_00992_));
 BUF_X4 _14368_ (.A(_07916_),
    .Z(_07922_));
 MUX2_X1 _14369_ (.A(_07855_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][55] ),
    .S(_07922_),
    .Z(_00993_));
 MUX2_X1 _14370_ (.A(_07858_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][56] ),
    .S(_07922_),
    .Z(_00994_));
 MUX2_X1 _14371_ (.A(_07860_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][57] ),
    .S(_07922_),
    .Z(_00995_));
 MUX2_X1 _14372_ (.A(_07862_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][58] ),
    .S(_07922_),
    .Z(_00996_));
 MUX2_X1 _14373_ (.A(_07864_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][59] ),
    .S(_07922_),
    .Z(_00997_));
 MUX2_X1 _14374_ (.A(_07866_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][5] ),
    .S(_07922_),
    .Z(_00998_));
 MUX2_X1 _14375_ (.A(_07868_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][60] ),
    .S(_07922_),
    .Z(_00999_));
 MUX2_X1 _14376_ (.A(_07870_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][61] ),
    .S(_07922_),
    .Z(_01000_));
 MUX2_X1 _14377_ (.A(_07872_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][62] ),
    .S(_07922_),
    .Z(_01001_));
 MUX2_X1 _14378_ (.A(_07874_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][63] ),
    .S(_07922_),
    .Z(_01002_));
 MUX2_X1 _14379_ (.A(_07876_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][6] ),
    .S(_07916_),
    .Z(_01003_));
 MUX2_X1 _14380_ (.A(_07878_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][7] ),
    .S(_07916_),
    .Z(_01004_));
 MUX2_X1 _14381_ (.A(_07880_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][8] ),
    .S(_07916_),
    .Z(_01005_));
 MUX2_X1 _14382_ (.A(_07882_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[13][9] ),
    .S(_07916_),
    .Z(_01006_));
 NAND2_X1 _14383_ (.A1(_10595_),
    .A2(_07914_),
    .ZN(_07923_));
 BUF_X4 _14384_ (.A(_07923_),
    .Z(_07924_));
 BUF_X4 _14385_ (.A(_07924_),
    .Z(_07925_));
 MUX2_X1 _14386_ (.A(_07745_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][0] ),
    .S(_07925_),
    .Z(_01007_));
 MUX2_X1 _14387_ (.A(_07753_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][10] ),
    .S(_07925_),
    .Z(_01008_));
 MUX2_X1 _14388_ (.A(_07755_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][11] ),
    .S(_07925_),
    .Z(_01009_));
 MUX2_X1 _14389_ (.A(_07757_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][12] ),
    .S(_07925_),
    .Z(_01010_));
 MUX2_X1 _14390_ (.A(_07759_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][13] ),
    .S(_07925_),
    .Z(_01011_));
 MUX2_X1 _14391_ (.A(_07761_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][14] ),
    .S(_07925_),
    .Z(_01012_));
 MUX2_X1 _14392_ (.A(_07763_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][15] ),
    .S(_07925_),
    .Z(_01013_));
 MUX2_X1 _14393_ (.A(_07765_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][16] ),
    .S(_07925_),
    .Z(_01014_));
 MUX2_X1 _14394_ (.A(_07767_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][17] ),
    .S(_07925_),
    .Z(_01015_));
 MUX2_X1 _14395_ (.A(_07769_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][18] ),
    .S(_07925_),
    .Z(_01016_));
 BUF_X4 _14396_ (.A(_07924_),
    .Z(_07926_));
 MUX2_X1 _14397_ (.A(_07771_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][19] ),
    .S(_07926_),
    .Z(_01017_));
 MUX2_X1 _14398_ (.A(_07774_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][1] ),
    .S(_07926_),
    .Z(_01018_));
 MUX2_X1 _14399_ (.A(_07776_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][20] ),
    .S(_07926_),
    .Z(_01019_));
 MUX2_X1 _14400_ (.A(_07778_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][21] ),
    .S(_07926_),
    .Z(_01020_));
 MUX2_X1 _14401_ (.A(_07780_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][22] ),
    .S(_07926_),
    .Z(_01021_));
 MUX2_X1 _14402_ (.A(_07782_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][23] ),
    .S(_07926_),
    .Z(_01022_));
 MUX2_X1 _14403_ (.A(_07784_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][24] ),
    .S(_07926_),
    .Z(_01023_));
 MUX2_X1 _14404_ (.A(_07786_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][25] ),
    .S(_07926_),
    .Z(_01024_));
 MUX2_X1 _14405_ (.A(_07788_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][26] ),
    .S(_07926_),
    .Z(_01025_));
 MUX2_X1 _14406_ (.A(_07790_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][27] ),
    .S(_07926_),
    .Z(_01026_));
 BUF_X4 _14407_ (.A(_07924_),
    .Z(_07927_));
 MUX2_X1 _14408_ (.A(_07792_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][28] ),
    .S(_07927_),
    .Z(_01027_));
 MUX2_X1 _14409_ (.A(_07795_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][29] ),
    .S(_07927_),
    .Z(_01028_));
 MUX2_X1 _14410_ (.A(_07797_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][2] ),
    .S(_07927_),
    .Z(_01029_));
 MUX2_X1 _14411_ (.A(_07799_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][30] ),
    .S(_07927_),
    .Z(_01030_));
 MUX2_X1 _14412_ (.A(_07801_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][31] ),
    .S(_07927_),
    .Z(_01031_));
 MUX2_X1 _14413_ (.A(_07803_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][32] ),
    .S(_07927_),
    .Z(_01032_));
 MUX2_X1 _14414_ (.A(_07805_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][33] ),
    .S(_07927_),
    .Z(_01033_));
 MUX2_X1 _14415_ (.A(_07807_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][34] ),
    .S(_07927_),
    .Z(_01034_));
 MUX2_X1 _14416_ (.A(_07809_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][35] ),
    .S(_07927_),
    .Z(_01035_));
 MUX2_X1 _14417_ (.A(_07811_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][36] ),
    .S(_07927_),
    .Z(_01036_));
 BUF_X4 _14418_ (.A(_07924_),
    .Z(_07928_));
 MUX2_X1 _14419_ (.A(_07813_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][37] ),
    .S(_07928_),
    .Z(_01037_));
 MUX2_X1 _14420_ (.A(_07816_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][38] ),
    .S(_07928_),
    .Z(_01038_));
 MUX2_X1 _14421_ (.A(_07818_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][39] ),
    .S(_07928_),
    .Z(_01039_));
 MUX2_X1 _14422_ (.A(_07820_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][3] ),
    .S(_07928_),
    .Z(_01040_));
 MUX2_X1 _14423_ (.A(_07822_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][40] ),
    .S(_07928_),
    .Z(_01041_));
 MUX2_X1 _14424_ (.A(_07824_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][41] ),
    .S(_07928_),
    .Z(_01042_));
 MUX2_X1 _14425_ (.A(_07826_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][42] ),
    .S(_07928_),
    .Z(_01043_));
 MUX2_X1 _14426_ (.A(_07828_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][43] ),
    .S(_07928_),
    .Z(_01044_));
 MUX2_X1 _14427_ (.A(_07830_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][44] ),
    .S(_07928_),
    .Z(_01045_));
 MUX2_X1 _14428_ (.A(_07832_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][45] ),
    .S(_07928_),
    .Z(_01046_));
 BUF_X4 _14429_ (.A(_07924_),
    .Z(_07929_));
 MUX2_X1 _14430_ (.A(_07834_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][46] ),
    .S(_07929_),
    .Z(_01047_));
 MUX2_X1 _14431_ (.A(_07837_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][47] ),
    .S(_07929_),
    .Z(_01048_));
 MUX2_X1 _14432_ (.A(_07839_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][48] ),
    .S(_07929_),
    .Z(_01049_));
 MUX2_X1 _14433_ (.A(_07841_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][49] ),
    .S(_07929_),
    .Z(_01050_));
 MUX2_X1 _14434_ (.A(_07843_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][4] ),
    .S(_07929_),
    .Z(_01051_));
 MUX2_X1 _14435_ (.A(_07845_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][50] ),
    .S(_07929_),
    .Z(_01052_));
 MUX2_X1 _14436_ (.A(_07847_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][51] ),
    .S(_07929_),
    .Z(_01053_));
 MUX2_X1 _14437_ (.A(_07849_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][52] ),
    .S(_07929_),
    .Z(_01054_));
 MUX2_X1 _14438_ (.A(_07851_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][53] ),
    .S(_07929_),
    .Z(_01055_));
 MUX2_X1 _14439_ (.A(_07853_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][54] ),
    .S(_07929_),
    .Z(_01056_));
 BUF_X4 _14440_ (.A(_07924_),
    .Z(_07930_));
 MUX2_X1 _14441_ (.A(_07855_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][55] ),
    .S(_07930_),
    .Z(_01057_));
 MUX2_X1 _14442_ (.A(_07858_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][56] ),
    .S(_07930_),
    .Z(_01058_));
 MUX2_X1 _14443_ (.A(_07860_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][57] ),
    .S(_07930_),
    .Z(_01059_));
 MUX2_X1 _14444_ (.A(_07862_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][58] ),
    .S(_07930_),
    .Z(_01060_));
 MUX2_X1 _14445_ (.A(_07864_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][59] ),
    .S(_07930_),
    .Z(_01061_));
 MUX2_X1 _14446_ (.A(_07866_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][5] ),
    .S(_07930_),
    .Z(_01062_));
 MUX2_X1 _14447_ (.A(_07868_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][60] ),
    .S(_07930_),
    .Z(_01063_));
 MUX2_X1 _14448_ (.A(_07870_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][61] ),
    .S(_07930_),
    .Z(_01064_));
 MUX2_X1 _14449_ (.A(_07872_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][62] ),
    .S(_07930_),
    .Z(_01065_));
 MUX2_X1 _14450_ (.A(_07874_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][63] ),
    .S(_07930_),
    .Z(_01066_));
 MUX2_X1 _14451_ (.A(_07876_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][6] ),
    .S(_07924_),
    .Z(_01067_));
 MUX2_X1 _14452_ (.A(_07878_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][7] ),
    .S(_07924_),
    .Z(_01068_));
 MUX2_X1 _14453_ (.A(_07880_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][8] ),
    .S(_07924_),
    .Z(_01069_));
 MUX2_X1 _14454_ (.A(_07882_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][9] ),
    .S(_07924_),
    .Z(_01070_));
 NAND2_X1 _14455_ (.A1(_07895_),
    .A2(_07914_),
    .ZN(_07931_));
 BUF_X4 _14456_ (.A(_07931_),
    .Z(_07932_));
 BUF_X4 _14457_ (.A(_07932_),
    .Z(_07933_));
 MUX2_X1 _14458_ (.A(_07745_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][0] ),
    .S(_07933_),
    .Z(_01071_));
 MUX2_X1 _14459_ (.A(_07753_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][10] ),
    .S(_07933_),
    .Z(_01072_));
 MUX2_X1 _14460_ (.A(_07755_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][11] ),
    .S(_07933_),
    .Z(_01073_));
 MUX2_X1 _14461_ (.A(_07757_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][12] ),
    .S(_07933_),
    .Z(_01074_));
 MUX2_X1 _14462_ (.A(_07759_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][13] ),
    .S(_07933_),
    .Z(_01075_));
 MUX2_X1 _14463_ (.A(_07761_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][14] ),
    .S(_07933_),
    .Z(_01076_));
 MUX2_X1 _14464_ (.A(_07763_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][15] ),
    .S(_07933_),
    .Z(_01077_));
 MUX2_X1 _14465_ (.A(_07765_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][16] ),
    .S(_07933_),
    .Z(_01078_));
 MUX2_X1 _14466_ (.A(_07767_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][17] ),
    .S(_07933_),
    .Z(_01079_));
 MUX2_X1 _14467_ (.A(_07769_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][18] ),
    .S(_07933_),
    .Z(_01080_));
 BUF_X4 _14468_ (.A(_07932_),
    .Z(_07934_));
 MUX2_X1 _14469_ (.A(_07771_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][19] ),
    .S(_07934_),
    .Z(_01081_));
 MUX2_X1 _14470_ (.A(_07774_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][1] ),
    .S(_07934_),
    .Z(_01082_));
 MUX2_X1 _14471_ (.A(_07776_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][20] ),
    .S(_07934_),
    .Z(_01083_));
 MUX2_X1 _14472_ (.A(_07778_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][21] ),
    .S(_07934_),
    .Z(_01084_));
 MUX2_X1 _14473_ (.A(_07780_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][22] ),
    .S(_07934_),
    .Z(_01085_));
 MUX2_X1 _14474_ (.A(_07782_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][23] ),
    .S(_07934_),
    .Z(_01086_));
 MUX2_X1 _14475_ (.A(_07784_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][24] ),
    .S(_07934_),
    .Z(_01087_));
 MUX2_X1 _14476_ (.A(_07786_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][25] ),
    .S(_07934_),
    .Z(_01088_));
 MUX2_X1 _14477_ (.A(_07788_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][26] ),
    .S(_07934_),
    .Z(_01089_));
 MUX2_X1 _14478_ (.A(_07790_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][27] ),
    .S(_07934_),
    .Z(_01090_));
 BUF_X4 _14479_ (.A(_07932_),
    .Z(_07935_));
 MUX2_X1 _14480_ (.A(_07792_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][28] ),
    .S(_07935_),
    .Z(_01091_));
 MUX2_X1 _14481_ (.A(_07795_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][29] ),
    .S(_07935_),
    .Z(_01092_));
 MUX2_X1 _14482_ (.A(_07797_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][2] ),
    .S(_07935_),
    .Z(_01093_));
 MUX2_X1 _14483_ (.A(_07799_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][30] ),
    .S(_07935_),
    .Z(_01094_));
 MUX2_X1 _14484_ (.A(_07801_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][31] ),
    .S(_07935_),
    .Z(_01095_));
 MUX2_X1 _14485_ (.A(_07803_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][32] ),
    .S(_07935_),
    .Z(_01096_));
 MUX2_X1 _14486_ (.A(_07805_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][33] ),
    .S(_07935_),
    .Z(_01097_));
 MUX2_X1 _14487_ (.A(_07807_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][34] ),
    .S(_07935_),
    .Z(_01098_));
 MUX2_X1 _14488_ (.A(_07809_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][35] ),
    .S(_07935_),
    .Z(_01099_));
 MUX2_X1 _14489_ (.A(_07811_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][36] ),
    .S(_07935_),
    .Z(_01100_));
 BUF_X4 _14490_ (.A(_07932_),
    .Z(_07936_));
 MUX2_X1 _14491_ (.A(_07813_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][37] ),
    .S(_07936_),
    .Z(_01101_));
 MUX2_X1 _14492_ (.A(_07816_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][38] ),
    .S(_07936_),
    .Z(_01102_));
 MUX2_X1 _14493_ (.A(_07818_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][39] ),
    .S(_07936_),
    .Z(_01103_));
 MUX2_X1 _14494_ (.A(_07820_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][3] ),
    .S(_07936_),
    .Z(_01104_));
 MUX2_X1 _14495_ (.A(_07822_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][40] ),
    .S(_07936_),
    .Z(_01105_));
 MUX2_X1 _14496_ (.A(_07824_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][41] ),
    .S(_07936_),
    .Z(_01106_));
 MUX2_X1 _14497_ (.A(_07826_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][42] ),
    .S(_07936_),
    .Z(_01107_));
 MUX2_X1 _14498_ (.A(_07828_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][43] ),
    .S(_07936_),
    .Z(_01108_));
 MUX2_X1 _14499_ (.A(_07830_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][44] ),
    .S(_07936_),
    .Z(_01109_));
 MUX2_X1 _14500_ (.A(_07832_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][45] ),
    .S(_07936_),
    .Z(_01110_));
 BUF_X4 _14501_ (.A(_07932_),
    .Z(_07937_));
 MUX2_X1 _14502_ (.A(_07834_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][46] ),
    .S(_07937_),
    .Z(_01111_));
 MUX2_X1 _14503_ (.A(_07837_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][47] ),
    .S(_07937_),
    .Z(_01112_));
 MUX2_X1 _14504_ (.A(_07839_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][48] ),
    .S(_07937_),
    .Z(_01113_));
 MUX2_X1 _14505_ (.A(_07841_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][49] ),
    .S(_07937_),
    .Z(_01114_));
 MUX2_X1 _14506_ (.A(_07843_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][4] ),
    .S(_07937_),
    .Z(_01115_));
 MUX2_X1 _14507_ (.A(_07845_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][50] ),
    .S(_07937_),
    .Z(_01116_));
 MUX2_X1 _14508_ (.A(_07847_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][51] ),
    .S(_07937_),
    .Z(_01117_));
 MUX2_X1 _14509_ (.A(_07849_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][52] ),
    .S(_07937_),
    .Z(_01118_));
 MUX2_X1 _14510_ (.A(_07851_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][53] ),
    .S(_07937_),
    .Z(_01119_));
 MUX2_X1 _14511_ (.A(_07853_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][54] ),
    .S(_07937_),
    .Z(_01120_));
 BUF_X4 _14512_ (.A(_07932_),
    .Z(_07938_));
 MUX2_X1 _14513_ (.A(_07855_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][55] ),
    .S(_07938_),
    .Z(_01121_));
 MUX2_X1 _14514_ (.A(_07858_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][56] ),
    .S(_07938_),
    .Z(_01122_));
 MUX2_X1 _14515_ (.A(_07860_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][57] ),
    .S(_07938_),
    .Z(_01123_));
 MUX2_X1 _14516_ (.A(_07862_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][58] ),
    .S(_07938_),
    .Z(_01124_));
 MUX2_X1 _14517_ (.A(_07864_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][59] ),
    .S(_07938_),
    .Z(_01125_));
 MUX2_X1 _14518_ (.A(_07866_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][5] ),
    .S(_07938_),
    .Z(_01126_));
 MUX2_X1 _14519_ (.A(_07868_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][60] ),
    .S(_07938_),
    .Z(_01127_));
 MUX2_X1 _14520_ (.A(_07870_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][61] ),
    .S(_07938_),
    .Z(_01128_));
 MUX2_X1 _14521_ (.A(_07872_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][62] ),
    .S(_07938_),
    .Z(_01129_));
 MUX2_X1 _14522_ (.A(_07874_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][63] ),
    .S(_07938_),
    .Z(_01130_));
 MUX2_X1 _14523_ (.A(_07876_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][6] ),
    .S(_07932_),
    .Z(_01131_));
 MUX2_X1 _14524_ (.A(_07878_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][7] ),
    .S(_07932_),
    .Z(_01132_));
 MUX2_X1 _14525_ (.A(_07880_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][8] ),
    .S(_07932_),
    .Z(_01133_));
 MUX2_X1 _14526_ (.A(_07882_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][9] ),
    .S(_07932_),
    .Z(_01134_));
 NOR3_X2 _14527_ (.A1(_06540_),
    .A2(_07746_),
    .A3(_07884_),
    .ZN(_07939_));
 NAND2_X1 _14528_ (.A1(_10597_),
    .A2(_07939_),
    .ZN(_07940_));
 BUF_X4 _14529_ (.A(_07940_),
    .Z(_07941_));
 CLKBUF_X3 _14530_ (.A(_07941_),
    .Z(_07942_));
 MUX2_X1 _14531_ (.A(_07745_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][0] ),
    .S(_07942_),
    .Z(_01135_));
 MUX2_X1 _14532_ (.A(_07753_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][10] ),
    .S(_07942_),
    .Z(_01136_));
 MUX2_X1 _14533_ (.A(_07755_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][11] ),
    .S(_07942_),
    .Z(_01137_));
 MUX2_X1 _14534_ (.A(_07757_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][12] ),
    .S(_07942_),
    .Z(_01138_));
 MUX2_X1 _14535_ (.A(_07759_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][13] ),
    .S(_07942_),
    .Z(_01139_));
 MUX2_X1 _14536_ (.A(_07761_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][14] ),
    .S(_07942_),
    .Z(_01140_));
 MUX2_X1 _14537_ (.A(_07763_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][15] ),
    .S(_07942_),
    .Z(_01141_));
 MUX2_X1 _14538_ (.A(_07765_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][16] ),
    .S(_07942_),
    .Z(_01142_));
 MUX2_X1 _14539_ (.A(_07767_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][17] ),
    .S(_07942_),
    .Z(_01143_));
 MUX2_X1 _14540_ (.A(_07769_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][18] ),
    .S(_07942_),
    .Z(_01144_));
 BUF_X4 _14541_ (.A(_07941_),
    .Z(_07943_));
 MUX2_X1 _14542_ (.A(_07771_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][19] ),
    .S(_07943_),
    .Z(_01145_));
 MUX2_X1 _14543_ (.A(_07774_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][1] ),
    .S(_07943_),
    .Z(_01146_));
 MUX2_X1 _14544_ (.A(_07776_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][20] ),
    .S(_07943_),
    .Z(_01147_));
 MUX2_X1 _14545_ (.A(_07778_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][21] ),
    .S(_07943_),
    .Z(_01148_));
 MUX2_X1 _14546_ (.A(_07780_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][22] ),
    .S(_07943_),
    .Z(_01149_));
 MUX2_X1 _14547_ (.A(_07782_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][23] ),
    .S(_07943_),
    .Z(_01150_));
 MUX2_X1 _14548_ (.A(_07784_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][24] ),
    .S(_07943_),
    .Z(_01151_));
 MUX2_X1 _14549_ (.A(_07786_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][25] ),
    .S(_07943_),
    .Z(_01152_));
 MUX2_X1 _14550_ (.A(_07788_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][26] ),
    .S(_07943_),
    .Z(_01153_));
 MUX2_X1 _14551_ (.A(_07790_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][27] ),
    .S(_07943_),
    .Z(_01154_));
 BUF_X4 _14552_ (.A(_07941_),
    .Z(_07944_));
 MUX2_X1 _14553_ (.A(_07792_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][28] ),
    .S(_07944_),
    .Z(_01155_));
 MUX2_X1 _14554_ (.A(_07795_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][29] ),
    .S(_07944_),
    .Z(_01156_));
 MUX2_X1 _14555_ (.A(_07797_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][2] ),
    .S(_07944_),
    .Z(_01157_));
 MUX2_X1 _14556_ (.A(_07799_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][30] ),
    .S(_07944_),
    .Z(_01158_));
 MUX2_X1 _14557_ (.A(_07801_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][31] ),
    .S(_07944_),
    .Z(_01159_));
 MUX2_X1 _14558_ (.A(_07803_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][32] ),
    .S(_07944_),
    .Z(_01160_));
 MUX2_X1 _14559_ (.A(_07805_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][33] ),
    .S(_07944_),
    .Z(_01161_));
 MUX2_X1 _14560_ (.A(_07807_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][34] ),
    .S(_07944_),
    .Z(_01162_));
 MUX2_X1 _14561_ (.A(_07809_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][35] ),
    .S(_07944_),
    .Z(_01163_));
 MUX2_X1 _14562_ (.A(_07811_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][36] ),
    .S(_07944_),
    .Z(_01164_));
 BUF_X4 _14563_ (.A(_07941_),
    .Z(_07945_));
 MUX2_X1 _14564_ (.A(_07813_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][37] ),
    .S(_07945_),
    .Z(_01165_));
 MUX2_X1 _14565_ (.A(_07816_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][38] ),
    .S(_07945_),
    .Z(_01166_));
 MUX2_X1 _14566_ (.A(_07818_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][39] ),
    .S(_07945_),
    .Z(_01167_));
 MUX2_X1 _14567_ (.A(_07820_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][3] ),
    .S(_07945_),
    .Z(_01168_));
 MUX2_X1 _14568_ (.A(_07822_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][40] ),
    .S(_07945_),
    .Z(_01169_));
 MUX2_X1 _14569_ (.A(_07824_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][41] ),
    .S(_07945_),
    .Z(_01170_));
 MUX2_X1 _14570_ (.A(_07826_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][42] ),
    .S(_07945_),
    .Z(_01171_));
 MUX2_X1 _14571_ (.A(_07828_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][43] ),
    .S(_07945_),
    .Z(_01172_));
 MUX2_X1 _14572_ (.A(_07830_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][44] ),
    .S(_07945_),
    .Z(_01173_));
 MUX2_X1 _14573_ (.A(_07832_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][45] ),
    .S(_07945_),
    .Z(_01174_));
 BUF_X4 _14574_ (.A(_07941_),
    .Z(_07946_));
 MUX2_X1 _14575_ (.A(_07834_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][46] ),
    .S(_07946_),
    .Z(_01175_));
 MUX2_X1 _14576_ (.A(_07837_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][47] ),
    .S(_07946_),
    .Z(_01176_));
 MUX2_X1 _14577_ (.A(_07839_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][48] ),
    .S(_07946_),
    .Z(_01177_));
 MUX2_X1 _14578_ (.A(_07841_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][49] ),
    .S(_07946_),
    .Z(_01178_));
 MUX2_X1 _14579_ (.A(_07843_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][4] ),
    .S(_07946_),
    .Z(_01179_));
 MUX2_X1 _14580_ (.A(_07845_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][50] ),
    .S(_07946_),
    .Z(_01180_));
 MUX2_X1 _14581_ (.A(_07847_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][51] ),
    .S(_07946_),
    .Z(_01181_));
 MUX2_X1 _14582_ (.A(_07849_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][52] ),
    .S(_07946_),
    .Z(_01182_));
 MUX2_X1 _14583_ (.A(_07851_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][53] ),
    .S(_07946_),
    .Z(_01183_));
 MUX2_X1 _14584_ (.A(_07853_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][54] ),
    .S(_07946_),
    .Z(_01184_));
 BUF_X4 _14585_ (.A(_07941_),
    .Z(_07947_));
 MUX2_X1 _14586_ (.A(_07855_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][55] ),
    .S(_07947_),
    .Z(_01185_));
 MUX2_X1 _14587_ (.A(_07858_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][56] ),
    .S(_07947_),
    .Z(_01186_));
 MUX2_X1 _14588_ (.A(_07860_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][57] ),
    .S(_07947_),
    .Z(_01187_));
 MUX2_X1 _14589_ (.A(_07862_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][58] ),
    .S(_07947_),
    .Z(_01188_));
 MUX2_X1 _14590_ (.A(_07864_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][59] ),
    .S(_07947_),
    .Z(_01189_));
 MUX2_X1 _14591_ (.A(_07866_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][5] ),
    .S(_07947_),
    .Z(_01190_));
 MUX2_X1 _14592_ (.A(_07868_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][60] ),
    .S(_07947_),
    .Z(_01191_));
 MUX2_X1 _14593_ (.A(_07870_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][61] ),
    .S(_07947_),
    .Z(_01192_));
 MUX2_X1 _14594_ (.A(_07872_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][62] ),
    .S(_07947_),
    .Z(_01193_));
 MUX2_X1 _14595_ (.A(_07874_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][63] ),
    .S(_07947_),
    .Z(_01194_));
 MUX2_X1 _14596_ (.A(_07876_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][6] ),
    .S(_07941_),
    .Z(_01195_));
 MUX2_X1 _14597_ (.A(_07878_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][7] ),
    .S(_07941_),
    .Z(_01196_));
 MUX2_X1 _14598_ (.A(_07880_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][8] ),
    .S(_07941_),
    .Z(_01197_));
 MUX2_X1 _14599_ (.A(_07882_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[1][9] ),
    .S(_07941_),
    .Z(_01198_));
 NAND2_X1 _14600_ (.A1(_10595_),
    .A2(_07939_),
    .ZN(_07948_));
 BUF_X4 _14601_ (.A(_07948_),
    .Z(_07949_));
 CLKBUF_X3 _14602_ (.A(_07949_),
    .Z(_07950_));
 MUX2_X1 _14603_ (.A(_07744_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][0] ),
    .S(_07950_),
    .Z(_01199_));
 MUX2_X1 _14604_ (.A(_07752_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][10] ),
    .S(_07950_),
    .Z(_01200_));
 MUX2_X1 _14605_ (.A(_07754_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][11] ),
    .S(_07950_),
    .Z(_01201_));
 MUX2_X1 _14606_ (.A(_07756_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][12] ),
    .S(_07950_),
    .Z(_01202_));
 MUX2_X1 _14607_ (.A(_07758_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][13] ),
    .S(_07950_),
    .Z(_01203_));
 MUX2_X1 _14608_ (.A(_07760_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][14] ),
    .S(_07950_),
    .Z(_01204_));
 MUX2_X1 _14609_ (.A(_07762_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][15] ),
    .S(_07950_),
    .Z(_01205_));
 MUX2_X1 _14610_ (.A(_07764_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][16] ),
    .S(_07950_),
    .Z(_01206_));
 MUX2_X1 _14611_ (.A(_07766_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][17] ),
    .S(_07950_),
    .Z(_01207_));
 MUX2_X1 _14612_ (.A(_07768_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][18] ),
    .S(_07950_),
    .Z(_01208_));
 BUF_X4 _14613_ (.A(_07949_),
    .Z(_07951_));
 MUX2_X1 _14614_ (.A(_07770_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][19] ),
    .S(_07951_),
    .Z(_01209_));
 MUX2_X1 _14615_ (.A(_07773_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][1] ),
    .S(_07951_),
    .Z(_01210_));
 MUX2_X1 _14616_ (.A(_07775_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][20] ),
    .S(_07951_),
    .Z(_01211_));
 MUX2_X1 _14617_ (.A(_07777_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][21] ),
    .S(_07951_),
    .Z(_01212_));
 MUX2_X1 _14618_ (.A(_07779_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][22] ),
    .S(_07951_),
    .Z(_01213_));
 MUX2_X1 _14619_ (.A(_07781_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][23] ),
    .S(_07951_),
    .Z(_01214_));
 MUX2_X1 _14620_ (.A(_07783_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][24] ),
    .S(_07951_),
    .Z(_01215_));
 MUX2_X1 _14621_ (.A(_07785_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][25] ),
    .S(_07951_),
    .Z(_01216_));
 MUX2_X1 _14622_ (.A(_07787_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][26] ),
    .S(_07951_),
    .Z(_01217_));
 MUX2_X1 _14623_ (.A(_07789_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][27] ),
    .S(_07951_),
    .Z(_01218_));
 BUF_X4 _14624_ (.A(_07949_),
    .Z(_07952_));
 MUX2_X1 _14625_ (.A(_07791_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][28] ),
    .S(_07952_),
    .Z(_01219_));
 MUX2_X1 _14626_ (.A(_07794_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][29] ),
    .S(_07952_),
    .Z(_01220_));
 MUX2_X1 _14627_ (.A(_07796_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][2] ),
    .S(_07952_),
    .Z(_01221_));
 MUX2_X1 _14628_ (.A(_07798_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][30] ),
    .S(_07952_),
    .Z(_01222_));
 MUX2_X1 _14629_ (.A(_07800_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][31] ),
    .S(_07952_),
    .Z(_01223_));
 MUX2_X1 _14630_ (.A(_07802_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][32] ),
    .S(_07952_),
    .Z(_01224_));
 MUX2_X1 _14631_ (.A(_07804_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][33] ),
    .S(_07952_),
    .Z(_01225_));
 MUX2_X1 _14632_ (.A(_07806_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][34] ),
    .S(_07952_),
    .Z(_01226_));
 MUX2_X1 _14633_ (.A(_07808_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][35] ),
    .S(_07952_),
    .Z(_01227_));
 MUX2_X1 _14634_ (.A(_07810_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][36] ),
    .S(_07952_),
    .Z(_01228_));
 BUF_X4 _14635_ (.A(_07949_),
    .Z(_07953_));
 MUX2_X1 _14636_ (.A(_07812_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][37] ),
    .S(_07953_),
    .Z(_01229_));
 MUX2_X1 _14637_ (.A(_07815_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][38] ),
    .S(_07953_),
    .Z(_01230_));
 MUX2_X1 _14638_ (.A(_07817_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][39] ),
    .S(_07953_),
    .Z(_01231_));
 MUX2_X1 _14639_ (.A(_07819_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][3] ),
    .S(_07953_),
    .Z(_01232_));
 MUX2_X1 _14640_ (.A(_07821_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][40] ),
    .S(_07953_),
    .Z(_01233_));
 MUX2_X1 _14641_ (.A(_07823_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][41] ),
    .S(_07953_),
    .Z(_01234_));
 MUX2_X1 _14642_ (.A(_07825_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][42] ),
    .S(_07953_),
    .Z(_01235_));
 MUX2_X1 _14643_ (.A(_07827_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][43] ),
    .S(_07953_),
    .Z(_01236_));
 MUX2_X1 _14644_ (.A(_07829_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][44] ),
    .S(_07953_),
    .Z(_01237_));
 MUX2_X1 _14645_ (.A(_07831_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][45] ),
    .S(_07953_),
    .Z(_01238_));
 BUF_X4 _14646_ (.A(_07949_),
    .Z(_07954_));
 MUX2_X1 _14647_ (.A(_07833_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][46] ),
    .S(_07954_),
    .Z(_01239_));
 MUX2_X1 _14648_ (.A(_07836_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][47] ),
    .S(_07954_),
    .Z(_01240_));
 MUX2_X1 _14649_ (.A(_07838_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][48] ),
    .S(_07954_),
    .Z(_01241_));
 MUX2_X1 _14650_ (.A(_07840_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][49] ),
    .S(_07954_),
    .Z(_01242_));
 MUX2_X1 _14651_ (.A(_07842_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][4] ),
    .S(_07954_),
    .Z(_01243_));
 MUX2_X1 _14652_ (.A(_07844_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][50] ),
    .S(_07954_),
    .Z(_01244_));
 MUX2_X1 _14653_ (.A(_07846_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][51] ),
    .S(_07954_),
    .Z(_01245_));
 MUX2_X1 _14654_ (.A(_07848_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][52] ),
    .S(_07954_),
    .Z(_01246_));
 MUX2_X1 _14655_ (.A(_07850_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][53] ),
    .S(_07954_),
    .Z(_01247_));
 MUX2_X1 _14656_ (.A(_07852_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][54] ),
    .S(_07954_),
    .Z(_01248_));
 BUF_X4 _14657_ (.A(_07949_),
    .Z(_07955_));
 MUX2_X1 _14658_ (.A(_07854_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][55] ),
    .S(_07955_),
    .Z(_01249_));
 MUX2_X1 _14659_ (.A(_07857_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][56] ),
    .S(_07955_),
    .Z(_01250_));
 MUX2_X1 _14660_ (.A(_07859_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][57] ),
    .S(_07955_),
    .Z(_01251_));
 MUX2_X1 _14661_ (.A(_07861_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][58] ),
    .S(_07955_),
    .Z(_01252_));
 MUX2_X1 _14662_ (.A(_07863_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][59] ),
    .S(_07955_),
    .Z(_01253_));
 MUX2_X1 _14663_ (.A(_07865_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][5] ),
    .S(_07955_),
    .Z(_01254_));
 MUX2_X1 _14664_ (.A(_07867_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][60] ),
    .S(_07955_),
    .Z(_01255_));
 MUX2_X1 _14665_ (.A(_07869_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][61] ),
    .S(_07955_),
    .Z(_01256_));
 MUX2_X1 _14666_ (.A(_07871_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][62] ),
    .S(_07955_),
    .Z(_01257_));
 MUX2_X1 _14667_ (.A(_07873_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][63] ),
    .S(_07955_),
    .Z(_01258_));
 MUX2_X1 _14668_ (.A(_07875_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][6] ),
    .S(_07949_),
    .Z(_01259_));
 MUX2_X1 _14669_ (.A(_07877_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][7] ),
    .S(_07949_),
    .Z(_01260_));
 MUX2_X1 _14670_ (.A(_07879_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][8] ),
    .S(_07949_),
    .Z(_01261_));
 MUX2_X1 _14671_ (.A(_07881_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][9] ),
    .S(_07949_),
    .Z(_01262_));
 NAND2_X1 _14672_ (.A1(_07895_),
    .A2(_07939_),
    .ZN(_07956_));
 BUF_X4 _14673_ (.A(_07956_),
    .Z(_07957_));
 CLKBUF_X3 _14674_ (.A(_07957_),
    .Z(_07958_));
 MUX2_X1 _14675_ (.A(_07744_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][0] ),
    .S(_07958_),
    .Z(_01263_));
 MUX2_X1 _14676_ (.A(_07752_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][10] ),
    .S(_07958_),
    .Z(_01264_));
 MUX2_X1 _14677_ (.A(_07754_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][11] ),
    .S(_07958_),
    .Z(_01265_));
 MUX2_X1 _14678_ (.A(_07756_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][12] ),
    .S(_07958_),
    .Z(_01266_));
 MUX2_X1 _14679_ (.A(_07758_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][13] ),
    .S(_07958_),
    .Z(_01267_));
 MUX2_X1 _14680_ (.A(_07760_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][14] ),
    .S(_07958_),
    .Z(_01268_));
 MUX2_X1 _14681_ (.A(_07762_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][15] ),
    .S(_07958_),
    .Z(_01269_));
 MUX2_X1 _14682_ (.A(_07764_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][16] ),
    .S(_07958_),
    .Z(_01270_));
 MUX2_X1 _14683_ (.A(_07766_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][17] ),
    .S(_07958_),
    .Z(_01271_));
 MUX2_X1 _14684_ (.A(_07768_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][18] ),
    .S(_07958_),
    .Z(_01272_));
 BUF_X4 _14685_ (.A(_07957_),
    .Z(_07959_));
 MUX2_X1 _14686_ (.A(_07770_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][19] ),
    .S(_07959_),
    .Z(_01273_));
 MUX2_X1 _14687_ (.A(_07773_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][1] ),
    .S(_07959_),
    .Z(_01274_));
 MUX2_X1 _14688_ (.A(_07775_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][20] ),
    .S(_07959_),
    .Z(_01275_));
 MUX2_X1 _14689_ (.A(_07777_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][21] ),
    .S(_07959_),
    .Z(_01276_));
 MUX2_X1 _14690_ (.A(_07779_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][22] ),
    .S(_07959_),
    .Z(_01277_));
 MUX2_X1 _14691_ (.A(_07781_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][23] ),
    .S(_07959_),
    .Z(_01278_));
 MUX2_X1 _14692_ (.A(_07783_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][24] ),
    .S(_07959_),
    .Z(_01279_));
 MUX2_X1 _14693_ (.A(_07785_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][25] ),
    .S(_07959_),
    .Z(_01280_));
 MUX2_X1 _14694_ (.A(_07787_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][26] ),
    .S(_07959_),
    .Z(_01281_));
 MUX2_X1 _14695_ (.A(_07789_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][27] ),
    .S(_07959_),
    .Z(_01282_));
 BUF_X4 _14696_ (.A(_07957_),
    .Z(_07960_));
 MUX2_X1 _14697_ (.A(_07791_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][28] ),
    .S(_07960_),
    .Z(_01283_));
 MUX2_X1 _14698_ (.A(_07794_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][29] ),
    .S(_07960_),
    .Z(_01284_));
 MUX2_X1 _14699_ (.A(_07796_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][2] ),
    .S(_07960_),
    .Z(_01285_));
 MUX2_X1 _14700_ (.A(_07798_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][30] ),
    .S(_07960_),
    .Z(_01286_));
 MUX2_X1 _14701_ (.A(_07800_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][31] ),
    .S(_07960_),
    .Z(_01287_));
 MUX2_X1 _14702_ (.A(_07802_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][32] ),
    .S(_07960_),
    .Z(_01288_));
 MUX2_X1 _14703_ (.A(_07804_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][33] ),
    .S(_07960_),
    .Z(_01289_));
 MUX2_X1 _14704_ (.A(_07806_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][34] ),
    .S(_07960_),
    .Z(_01290_));
 MUX2_X1 _14705_ (.A(_07808_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][35] ),
    .S(_07960_),
    .Z(_01291_));
 MUX2_X1 _14706_ (.A(_07810_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][36] ),
    .S(_07960_),
    .Z(_01292_));
 BUF_X4 _14707_ (.A(_07957_),
    .Z(_07961_));
 MUX2_X1 _14708_ (.A(_07812_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][37] ),
    .S(_07961_),
    .Z(_01293_));
 MUX2_X1 _14709_ (.A(_07815_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][38] ),
    .S(_07961_),
    .Z(_01294_));
 MUX2_X1 _14710_ (.A(_07817_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][39] ),
    .S(_07961_),
    .Z(_01295_));
 MUX2_X1 _14711_ (.A(_07819_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][3] ),
    .S(_07961_),
    .Z(_01296_));
 MUX2_X1 _14712_ (.A(_07821_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][40] ),
    .S(_07961_),
    .Z(_01297_));
 MUX2_X1 _14713_ (.A(_07823_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][41] ),
    .S(_07961_),
    .Z(_01298_));
 MUX2_X1 _14714_ (.A(_07825_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][42] ),
    .S(_07961_),
    .Z(_01299_));
 MUX2_X1 _14715_ (.A(_07827_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][43] ),
    .S(_07961_),
    .Z(_01300_));
 MUX2_X1 _14716_ (.A(_07829_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][44] ),
    .S(_07961_),
    .Z(_01301_));
 MUX2_X1 _14717_ (.A(_07831_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][45] ),
    .S(_07961_),
    .Z(_01302_));
 BUF_X4 _14718_ (.A(_07957_),
    .Z(_07962_));
 MUX2_X1 _14719_ (.A(_07833_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][46] ),
    .S(_07962_),
    .Z(_01303_));
 MUX2_X1 _14720_ (.A(_07836_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][47] ),
    .S(_07962_),
    .Z(_01304_));
 MUX2_X1 _14721_ (.A(_07838_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][48] ),
    .S(_07962_),
    .Z(_01305_));
 MUX2_X1 _14722_ (.A(_07840_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][49] ),
    .S(_07962_),
    .Z(_01306_));
 MUX2_X1 _14723_ (.A(_07842_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][4] ),
    .S(_07962_),
    .Z(_01307_));
 MUX2_X1 _14724_ (.A(_07844_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][50] ),
    .S(_07962_),
    .Z(_01308_));
 MUX2_X1 _14725_ (.A(_07846_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][51] ),
    .S(_07962_),
    .Z(_01309_));
 MUX2_X1 _14726_ (.A(_07848_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][52] ),
    .S(_07962_),
    .Z(_01310_));
 MUX2_X1 _14727_ (.A(_07850_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][53] ),
    .S(_07962_),
    .Z(_01311_));
 MUX2_X1 _14728_ (.A(_07852_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][54] ),
    .S(_07962_),
    .Z(_01312_));
 BUF_X4 _14729_ (.A(_07957_),
    .Z(_07963_));
 MUX2_X1 _14730_ (.A(_07854_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][55] ),
    .S(_07963_),
    .Z(_01313_));
 MUX2_X1 _14731_ (.A(_07857_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][56] ),
    .S(_07963_),
    .Z(_01314_));
 MUX2_X1 _14732_ (.A(_07859_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][57] ),
    .S(_07963_),
    .Z(_01315_));
 MUX2_X1 _14733_ (.A(_07861_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][58] ),
    .S(_07963_),
    .Z(_01316_));
 MUX2_X1 _14734_ (.A(_07863_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][59] ),
    .S(_07963_),
    .Z(_01317_));
 MUX2_X1 _14735_ (.A(_07865_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][5] ),
    .S(_07963_),
    .Z(_01318_));
 MUX2_X1 _14736_ (.A(_07867_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][60] ),
    .S(_07963_),
    .Z(_01319_));
 MUX2_X1 _14737_ (.A(_07869_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][61] ),
    .S(_07963_),
    .Z(_01320_));
 MUX2_X1 _14738_ (.A(_07871_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][62] ),
    .S(_07963_),
    .Z(_01321_));
 MUX2_X1 _14739_ (.A(_07873_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][63] ),
    .S(_07963_),
    .Z(_01322_));
 MUX2_X1 _14740_ (.A(_07875_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][6] ),
    .S(_07957_),
    .Z(_01323_));
 MUX2_X1 _14741_ (.A(_07877_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][7] ),
    .S(_07957_),
    .Z(_01324_));
 MUX2_X1 _14742_ (.A(_07879_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][8] ),
    .S(_07957_),
    .Z(_01325_));
 MUX2_X1 _14743_ (.A(_07881_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][9] ),
    .S(_07957_),
    .Z(_01326_));
 NOR3_X1 _14744_ (.A1(_06540_),
    .A2(_07746_),
    .A3(_07904_),
    .ZN(_07964_));
 BUF_X4 _14745_ (.A(_07964_),
    .Z(_07965_));
 CLKBUF_X3 _14746_ (.A(_07965_),
    .Z(_07966_));
 MUX2_X1 _14747_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][0] ),
    .B(_07745_),
    .S(_07966_),
    .Z(_01327_));
 MUX2_X1 _14748_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][10] ),
    .B(_07753_),
    .S(_07966_),
    .Z(_01328_));
 MUX2_X1 _14749_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][11] ),
    .B(_07755_),
    .S(_07966_),
    .Z(_01329_));
 MUX2_X1 _14750_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][12] ),
    .B(_07757_),
    .S(_07966_),
    .Z(_01330_));
 MUX2_X1 _14751_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][13] ),
    .B(_07759_),
    .S(_07966_),
    .Z(_01331_));
 MUX2_X1 _14752_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][14] ),
    .B(_07761_),
    .S(_07966_),
    .Z(_01332_));
 MUX2_X1 _14753_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][15] ),
    .B(_07763_),
    .S(_07966_),
    .Z(_01333_));
 MUX2_X1 _14754_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][16] ),
    .B(_07765_),
    .S(_07966_),
    .Z(_01334_));
 MUX2_X1 _14755_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][17] ),
    .B(_07767_),
    .S(_07966_),
    .Z(_01335_));
 MUX2_X1 _14756_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][18] ),
    .B(_07769_),
    .S(_07966_),
    .Z(_01336_));
 BUF_X4 _14757_ (.A(_07965_),
    .Z(_07967_));
 MUX2_X1 _14758_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][19] ),
    .B(_07771_),
    .S(_07967_),
    .Z(_01337_));
 MUX2_X1 _14759_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][1] ),
    .B(_07774_),
    .S(_07967_),
    .Z(_01338_));
 MUX2_X1 _14760_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][20] ),
    .B(_07776_),
    .S(_07967_),
    .Z(_01339_));
 MUX2_X1 _14761_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][21] ),
    .B(_07778_),
    .S(_07967_),
    .Z(_01340_));
 MUX2_X1 _14762_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][22] ),
    .B(_07780_),
    .S(_07967_),
    .Z(_01341_));
 MUX2_X1 _14763_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][23] ),
    .B(_07782_),
    .S(_07967_),
    .Z(_01342_));
 MUX2_X1 _14764_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][24] ),
    .B(_07784_),
    .S(_07967_),
    .Z(_01343_));
 MUX2_X1 _14765_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][25] ),
    .B(_07786_),
    .S(_07967_),
    .Z(_01344_));
 MUX2_X1 _14766_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][26] ),
    .B(_07788_),
    .S(_07967_),
    .Z(_01345_));
 MUX2_X1 _14767_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][27] ),
    .B(_07790_),
    .S(_07967_),
    .Z(_01346_));
 BUF_X4 _14768_ (.A(_07965_),
    .Z(_07968_));
 MUX2_X1 _14769_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][28] ),
    .B(_07792_),
    .S(_07968_),
    .Z(_01347_));
 MUX2_X1 _14770_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][29] ),
    .B(_07795_),
    .S(_07968_),
    .Z(_01348_));
 MUX2_X1 _14771_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][2] ),
    .B(_07797_),
    .S(_07968_),
    .Z(_01349_));
 MUX2_X1 _14772_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][30] ),
    .B(_07799_),
    .S(_07968_),
    .Z(_01350_));
 MUX2_X1 _14773_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][31] ),
    .B(_07801_),
    .S(_07968_),
    .Z(_01351_));
 MUX2_X1 _14774_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][32] ),
    .B(_07803_),
    .S(_07968_),
    .Z(_01352_));
 MUX2_X1 _14775_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][33] ),
    .B(_07805_),
    .S(_07968_),
    .Z(_01353_));
 MUX2_X1 _14776_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][34] ),
    .B(_07807_),
    .S(_07968_),
    .Z(_01354_));
 MUX2_X1 _14777_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][35] ),
    .B(_07809_),
    .S(_07968_),
    .Z(_01355_));
 MUX2_X1 _14778_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][36] ),
    .B(_07811_),
    .S(_07968_),
    .Z(_01356_));
 BUF_X4 _14779_ (.A(_07965_),
    .Z(_07969_));
 MUX2_X1 _14780_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][37] ),
    .B(_07813_),
    .S(_07969_),
    .Z(_01357_));
 MUX2_X1 _14781_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][38] ),
    .B(_07816_),
    .S(_07969_),
    .Z(_01358_));
 MUX2_X1 _14782_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][39] ),
    .B(_07818_),
    .S(_07969_),
    .Z(_01359_));
 MUX2_X1 _14783_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][3] ),
    .B(_07820_),
    .S(_07969_),
    .Z(_01360_));
 MUX2_X1 _14784_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][40] ),
    .B(_07822_),
    .S(_07969_),
    .Z(_01361_));
 MUX2_X1 _14785_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][41] ),
    .B(_07824_),
    .S(_07969_),
    .Z(_01362_));
 MUX2_X1 _14786_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][42] ),
    .B(_07826_),
    .S(_07969_),
    .Z(_01363_));
 MUX2_X1 _14787_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][43] ),
    .B(_07828_),
    .S(_07969_),
    .Z(_01364_));
 MUX2_X1 _14788_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][44] ),
    .B(_07830_),
    .S(_07969_),
    .Z(_01365_));
 MUX2_X1 _14789_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][45] ),
    .B(_07832_),
    .S(_07969_),
    .Z(_01366_));
 BUF_X4 _14790_ (.A(_07965_),
    .Z(_07970_));
 MUX2_X1 _14791_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][46] ),
    .B(_07834_),
    .S(_07970_),
    .Z(_01367_));
 MUX2_X1 _14792_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][47] ),
    .B(_07837_),
    .S(_07970_),
    .Z(_01368_));
 MUX2_X1 _14793_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][48] ),
    .B(_07839_),
    .S(_07970_),
    .Z(_01369_));
 MUX2_X1 _14794_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][49] ),
    .B(_07841_),
    .S(_07970_),
    .Z(_01370_));
 MUX2_X1 _14795_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][4] ),
    .B(_07843_),
    .S(_07970_),
    .Z(_01371_));
 MUX2_X1 _14796_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][50] ),
    .B(_07845_),
    .S(_07970_),
    .Z(_01372_));
 MUX2_X1 _14797_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][51] ),
    .B(_07847_),
    .S(_07970_),
    .Z(_01373_));
 MUX2_X1 _14798_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][52] ),
    .B(_07849_),
    .S(_07970_),
    .Z(_01374_));
 MUX2_X1 _14799_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][53] ),
    .B(_07851_),
    .S(_07970_),
    .Z(_01375_));
 MUX2_X1 _14800_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][54] ),
    .B(_07853_),
    .S(_07970_),
    .Z(_01376_));
 BUF_X4 _14801_ (.A(_07965_),
    .Z(_07971_));
 MUX2_X1 _14802_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][55] ),
    .B(_07855_),
    .S(_07971_),
    .Z(_01377_));
 MUX2_X1 _14803_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][56] ),
    .B(_07858_),
    .S(_07971_),
    .Z(_01378_));
 MUX2_X1 _14804_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][57] ),
    .B(_07860_),
    .S(_07971_),
    .Z(_01379_));
 MUX2_X1 _14805_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][58] ),
    .B(_07862_),
    .S(_07971_),
    .Z(_01380_));
 MUX2_X1 _14806_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][59] ),
    .B(_07864_),
    .S(_07971_),
    .Z(_01381_));
 MUX2_X1 _14807_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][5] ),
    .B(_07866_),
    .S(_07971_),
    .Z(_01382_));
 MUX2_X1 _14808_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][60] ),
    .B(_07868_),
    .S(_07971_),
    .Z(_01383_));
 MUX2_X1 _14809_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][61] ),
    .B(_07870_),
    .S(_07971_),
    .Z(_01384_));
 MUX2_X1 _14810_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][62] ),
    .B(_07872_),
    .S(_07971_),
    .Z(_01385_));
 MUX2_X1 _14811_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][63] ),
    .B(_07874_),
    .S(_07971_),
    .Z(_01386_));
 MUX2_X1 _14812_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][6] ),
    .B(_07876_),
    .S(_07965_),
    .Z(_01387_));
 MUX2_X1 _14813_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][7] ),
    .B(_07878_),
    .S(_07965_),
    .Z(_01388_));
 MUX2_X1 _14814_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][8] ),
    .B(_07880_),
    .S(_07965_),
    .Z(_01389_));
 MUX2_X1 _14815_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][9] ),
    .B(_07882_),
    .S(_07965_),
    .Z(_01390_));
 NOR3_X2 _14816_ (.A1(_06539_),
    .A2(_07746_),
    .A3(_07913_),
    .ZN(_07972_));
 NAND2_X1 _14817_ (.A1(_10597_),
    .A2(_07972_),
    .ZN(_07973_));
 BUF_X4 _14818_ (.A(_07973_),
    .Z(_07974_));
 CLKBUF_X3 _14819_ (.A(_07974_),
    .Z(_07975_));
 MUX2_X1 _14820_ (.A(_07744_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][0] ),
    .S(_07975_),
    .Z(_01391_));
 MUX2_X1 _14821_ (.A(_07752_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][10] ),
    .S(_07975_),
    .Z(_01392_));
 MUX2_X1 _14822_ (.A(_07754_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][11] ),
    .S(_07975_),
    .Z(_01393_));
 MUX2_X1 _14823_ (.A(_07756_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][12] ),
    .S(_07975_),
    .Z(_01394_));
 MUX2_X1 _14824_ (.A(_07758_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][13] ),
    .S(_07975_),
    .Z(_01395_));
 MUX2_X1 _14825_ (.A(_07760_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][14] ),
    .S(_07975_),
    .Z(_01396_));
 MUX2_X1 _14826_ (.A(_07762_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][15] ),
    .S(_07975_),
    .Z(_01397_));
 MUX2_X1 _14827_ (.A(_07764_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][16] ),
    .S(_07975_),
    .Z(_01398_));
 MUX2_X1 _14828_ (.A(_07766_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][17] ),
    .S(_07975_),
    .Z(_01399_));
 MUX2_X1 _14829_ (.A(_07768_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][18] ),
    .S(_07975_),
    .Z(_01400_));
 BUF_X4 _14830_ (.A(_07974_),
    .Z(_07976_));
 MUX2_X1 _14831_ (.A(_07770_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][19] ),
    .S(_07976_),
    .Z(_01401_));
 MUX2_X1 _14832_ (.A(_07773_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][1] ),
    .S(_07976_),
    .Z(_01402_));
 MUX2_X1 _14833_ (.A(_07775_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][20] ),
    .S(_07976_),
    .Z(_01403_));
 MUX2_X1 _14834_ (.A(_07777_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][21] ),
    .S(_07976_),
    .Z(_01404_));
 MUX2_X1 _14835_ (.A(_07779_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][22] ),
    .S(_07976_),
    .Z(_01405_));
 MUX2_X1 _14836_ (.A(_07781_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][23] ),
    .S(_07976_),
    .Z(_01406_));
 MUX2_X1 _14837_ (.A(_07783_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][24] ),
    .S(_07976_),
    .Z(_01407_));
 MUX2_X1 _14838_ (.A(_07785_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][25] ),
    .S(_07976_),
    .Z(_01408_));
 MUX2_X1 _14839_ (.A(_07787_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][26] ),
    .S(_07976_),
    .Z(_01409_));
 MUX2_X1 _14840_ (.A(_07789_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][27] ),
    .S(_07976_),
    .Z(_01410_));
 BUF_X4 _14841_ (.A(_07974_),
    .Z(_07977_));
 MUX2_X1 _14842_ (.A(_07791_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][28] ),
    .S(_07977_),
    .Z(_01411_));
 MUX2_X1 _14843_ (.A(_07794_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][29] ),
    .S(_07977_),
    .Z(_01412_));
 MUX2_X1 _14844_ (.A(_07796_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][2] ),
    .S(_07977_),
    .Z(_01413_));
 MUX2_X1 _14845_ (.A(_07798_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][30] ),
    .S(_07977_),
    .Z(_01414_));
 MUX2_X1 _14846_ (.A(_07800_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][31] ),
    .S(_07977_),
    .Z(_01415_));
 MUX2_X1 _14847_ (.A(_07802_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][32] ),
    .S(_07977_),
    .Z(_01416_));
 MUX2_X1 _14848_ (.A(_07804_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][33] ),
    .S(_07977_),
    .Z(_01417_));
 MUX2_X1 _14849_ (.A(_07806_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][34] ),
    .S(_07977_),
    .Z(_01418_));
 MUX2_X1 _14850_ (.A(_07808_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][35] ),
    .S(_07977_),
    .Z(_01419_));
 MUX2_X1 _14851_ (.A(_07810_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][36] ),
    .S(_07977_),
    .Z(_01420_));
 BUF_X4 _14852_ (.A(_07974_),
    .Z(_07978_));
 MUX2_X1 _14853_ (.A(_07812_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][37] ),
    .S(_07978_),
    .Z(_01421_));
 MUX2_X1 _14854_ (.A(_07815_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][38] ),
    .S(_07978_),
    .Z(_01422_));
 MUX2_X1 _14855_ (.A(_07817_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][39] ),
    .S(_07978_),
    .Z(_01423_));
 MUX2_X1 _14856_ (.A(_07819_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][3] ),
    .S(_07978_),
    .Z(_01424_));
 MUX2_X1 _14857_ (.A(_07821_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][40] ),
    .S(_07978_),
    .Z(_01425_));
 MUX2_X1 _14858_ (.A(_07823_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][41] ),
    .S(_07978_),
    .Z(_01426_));
 MUX2_X1 _14859_ (.A(_07825_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][42] ),
    .S(_07978_),
    .Z(_01427_));
 MUX2_X1 _14860_ (.A(_07827_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][43] ),
    .S(_07978_),
    .Z(_01428_));
 MUX2_X1 _14861_ (.A(_07829_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][44] ),
    .S(_07978_),
    .Z(_01429_));
 MUX2_X1 _14862_ (.A(_07831_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][45] ),
    .S(_07978_),
    .Z(_01430_));
 BUF_X4 _14863_ (.A(_07974_),
    .Z(_07979_));
 MUX2_X1 _14864_ (.A(_07833_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][46] ),
    .S(_07979_),
    .Z(_01431_));
 MUX2_X1 _14865_ (.A(_07836_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][47] ),
    .S(_07979_),
    .Z(_01432_));
 MUX2_X1 _14866_ (.A(_07838_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][48] ),
    .S(_07979_),
    .Z(_01433_));
 MUX2_X1 _14867_ (.A(_07840_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][49] ),
    .S(_07979_),
    .Z(_01434_));
 MUX2_X1 _14868_ (.A(_07842_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][4] ),
    .S(_07979_),
    .Z(_01435_));
 MUX2_X1 _14869_ (.A(_07844_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][50] ),
    .S(_07979_),
    .Z(_01436_));
 MUX2_X1 _14870_ (.A(_07846_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][51] ),
    .S(_07979_),
    .Z(_01437_));
 MUX2_X1 _14871_ (.A(_07848_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][52] ),
    .S(_07979_),
    .Z(_01438_));
 MUX2_X1 _14872_ (.A(_07850_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][53] ),
    .S(_07979_),
    .Z(_01439_));
 MUX2_X1 _14873_ (.A(_07852_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][54] ),
    .S(_07979_),
    .Z(_01440_));
 BUF_X4 _14874_ (.A(_07974_),
    .Z(_07980_));
 MUX2_X1 _14875_ (.A(_07854_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][55] ),
    .S(_07980_),
    .Z(_01441_));
 MUX2_X1 _14876_ (.A(_07857_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][56] ),
    .S(_07980_),
    .Z(_01442_));
 MUX2_X1 _14877_ (.A(_07859_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][57] ),
    .S(_07980_),
    .Z(_01443_));
 MUX2_X1 _14878_ (.A(_07861_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][58] ),
    .S(_07980_),
    .Z(_01444_));
 MUX2_X1 _14879_ (.A(_07863_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][59] ),
    .S(_07980_),
    .Z(_01445_));
 MUX2_X1 _14880_ (.A(_07865_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][5] ),
    .S(_07980_),
    .Z(_01446_));
 MUX2_X1 _14881_ (.A(_07867_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][60] ),
    .S(_07980_),
    .Z(_01447_));
 MUX2_X1 _14882_ (.A(_07869_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][61] ),
    .S(_07980_),
    .Z(_01448_));
 MUX2_X1 _14883_ (.A(_07871_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][62] ),
    .S(_07980_),
    .Z(_01449_));
 MUX2_X1 _14884_ (.A(_07873_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][63] ),
    .S(_07980_),
    .Z(_01450_));
 MUX2_X1 _14885_ (.A(_07875_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][6] ),
    .S(_07974_),
    .Z(_01451_));
 MUX2_X1 _14886_ (.A(_07877_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][7] ),
    .S(_07974_),
    .Z(_01452_));
 MUX2_X1 _14887_ (.A(_07879_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][8] ),
    .S(_07974_),
    .Z(_01453_));
 MUX2_X1 _14888_ (.A(_07881_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[5][9] ),
    .S(_07974_),
    .Z(_01454_));
 NAND2_X1 _14889_ (.A1(_10595_),
    .A2(_07972_),
    .ZN(_07981_));
 BUF_X4 _14890_ (.A(_07981_),
    .Z(_07982_));
 CLKBUF_X3 _14891_ (.A(_07982_),
    .Z(_07983_));
 MUX2_X1 _14892_ (.A(_07744_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][0] ),
    .S(_07983_),
    .Z(_01455_));
 MUX2_X1 _14893_ (.A(_07752_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][10] ),
    .S(_07983_),
    .Z(_01456_));
 MUX2_X1 _14894_ (.A(_07754_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][11] ),
    .S(_07983_),
    .Z(_01457_));
 MUX2_X1 _14895_ (.A(_07756_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][12] ),
    .S(_07983_),
    .Z(_01458_));
 MUX2_X1 _14896_ (.A(_07758_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][13] ),
    .S(_07983_),
    .Z(_01459_));
 MUX2_X1 _14897_ (.A(_07760_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][14] ),
    .S(_07983_),
    .Z(_01460_));
 MUX2_X1 _14898_ (.A(_07762_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][15] ),
    .S(_07983_),
    .Z(_01461_));
 MUX2_X1 _14899_ (.A(_07764_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][16] ),
    .S(_07983_),
    .Z(_01462_));
 MUX2_X1 _14900_ (.A(_07766_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][17] ),
    .S(_07983_),
    .Z(_01463_));
 MUX2_X1 _14901_ (.A(_07768_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][18] ),
    .S(_07983_),
    .Z(_01464_));
 BUF_X4 _14902_ (.A(_07982_),
    .Z(_07984_));
 MUX2_X1 _14903_ (.A(_07770_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][19] ),
    .S(_07984_),
    .Z(_01465_));
 MUX2_X1 _14904_ (.A(_07773_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][1] ),
    .S(_07984_),
    .Z(_01466_));
 MUX2_X1 _14905_ (.A(_07775_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][20] ),
    .S(_07984_),
    .Z(_01467_));
 MUX2_X1 _14906_ (.A(_07777_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][21] ),
    .S(_07984_),
    .Z(_01468_));
 MUX2_X1 _14907_ (.A(_07779_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][22] ),
    .S(_07984_),
    .Z(_01469_));
 MUX2_X1 _14908_ (.A(_07781_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][23] ),
    .S(_07984_),
    .Z(_01470_));
 MUX2_X1 _14909_ (.A(_07783_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][24] ),
    .S(_07984_),
    .Z(_01471_));
 MUX2_X1 _14910_ (.A(_07785_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][25] ),
    .S(_07984_),
    .Z(_01472_));
 MUX2_X1 _14911_ (.A(_07787_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][26] ),
    .S(_07984_),
    .Z(_01473_));
 MUX2_X1 _14912_ (.A(_07789_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][27] ),
    .S(_07984_),
    .Z(_01474_));
 BUF_X4 _14913_ (.A(_07982_),
    .Z(_07985_));
 MUX2_X1 _14914_ (.A(_07791_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][28] ),
    .S(_07985_),
    .Z(_01475_));
 MUX2_X1 _14915_ (.A(_07794_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][29] ),
    .S(_07985_),
    .Z(_01476_));
 MUX2_X1 _14916_ (.A(_07796_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][2] ),
    .S(_07985_),
    .Z(_01477_));
 MUX2_X1 _14917_ (.A(_07798_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][30] ),
    .S(_07985_),
    .Z(_01478_));
 MUX2_X1 _14918_ (.A(_07800_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][31] ),
    .S(_07985_),
    .Z(_01479_));
 MUX2_X1 _14919_ (.A(_07802_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][32] ),
    .S(_07985_),
    .Z(_01480_));
 MUX2_X1 _14920_ (.A(_07804_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][33] ),
    .S(_07985_),
    .Z(_01481_));
 MUX2_X1 _14921_ (.A(_07806_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][34] ),
    .S(_07985_),
    .Z(_01482_));
 MUX2_X1 _14922_ (.A(_07808_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][35] ),
    .S(_07985_),
    .Z(_01483_));
 MUX2_X1 _14923_ (.A(_07810_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][36] ),
    .S(_07985_),
    .Z(_01484_));
 BUF_X4 _14924_ (.A(_07982_),
    .Z(_07986_));
 MUX2_X1 _14925_ (.A(_07812_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][37] ),
    .S(_07986_),
    .Z(_01485_));
 MUX2_X1 _14926_ (.A(_07815_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][38] ),
    .S(_07986_),
    .Z(_01486_));
 MUX2_X1 _14927_ (.A(_07817_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][39] ),
    .S(_07986_),
    .Z(_01487_));
 MUX2_X1 _14928_ (.A(_07819_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][3] ),
    .S(_07986_),
    .Z(_01488_));
 MUX2_X1 _14929_ (.A(_07821_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][40] ),
    .S(_07986_),
    .Z(_01489_));
 MUX2_X1 _14930_ (.A(_07823_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][41] ),
    .S(_07986_),
    .Z(_01490_));
 MUX2_X1 _14931_ (.A(_07825_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][42] ),
    .S(_07986_),
    .Z(_01491_));
 MUX2_X1 _14932_ (.A(_07827_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][43] ),
    .S(_07986_),
    .Z(_01492_));
 MUX2_X1 _14933_ (.A(_07829_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][44] ),
    .S(_07986_),
    .Z(_01493_));
 MUX2_X1 _14934_ (.A(_07831_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][45] ),
    .S(_07986_),
    .Z(_01494_));
 BUF_X4 _14935_ (.A(_07982_),
    .Z(_07987_));
 MUX2_X1 _14936_ (.A(_07833_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][46] ),
    .S(_07987_),
    .Z(_01495_));
 MUX2_X1 _14937_ (.A(_07836_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][47] ),
    .S(_07987_),
    .Z(_01496_));
 MUX2_X1 _14938_ (.A(_07838_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][48] ),
    .S(_07987_),
    .Z(_01497_));
 MUX2_X1 _14939_ (.A(_07840_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][49] ),
    .S(_07987_),
    .Z(_01498_));
 MUX2_X1 _14940_ (.A(_07842_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][4] ),
    .S(_07987_),
    .Z(_01499_));
 MUX2_X1 _14941_ (.A(_07844_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][50] ),
    .S(_07987_),
    .Z(_01500_));
 MUX2_X1 _14942_ (.A(_07846_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][51] ),
    .S(_07987_),
    .Z(_01501_));
 MUX2_X1 _14943_ (.A(_07848_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][52] ),
    .S(_07987_),
    .Z(_01502_));
 MUX2_X1 _14944_ (.A(_07850_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][53] ),
    .S(_07987_),
    .Z(_01503_));
 MUX2_X1 _14945_ (.A(_07852_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][54] ),
    .S(_07987_),
    .Z(_01504_));
 BUF_X4 _14946_ (.A(_07982_),
    .Z(_07988_));
 MUX2_X1 _14947_ (.A(_07854_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][55] ),
    .S(_07988_),
    .Z(_01505_));
 MUX2_X1 _14948_ (.A(_07857_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][56] ),
    .S(_07988_),
    .Z(_01506_));
 MUX2_X1 _14949_ (.A(_07859_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][57] ),
    .S(_07988_),
    .Z(_01507_));
 MUX2_X1 _14950_ (.A(_07861_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][58] ),
    .S(_07988_),
    .Z(_01508_));
 MUX2_X1 _14951_ (.A(_07863_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][59] ),
    .S(_07988_),
    .Z(_01509_));
 MUX2_X1 _14952_ (.A(_07865_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][5] ),
    .S(_07988_),
    .Z(_01510_));
 MUX2_X1 _14953_ (.A(_07867_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][60] ),
    .S(_07988_),
    .Z(_01511_));
 MUX2_X1 _14954_ (.A(_07869_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][61] ),
    .S(_07988_),
    .Z(_01512_));
 MUX2_X1 _14955_ (.A(_07871_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][62] ),
    .S(_07988_),
    .Z(_01513_));
 MUX2_X1 _14956_ (.A(_07873_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][63] ),
    .S(_07988_),
    .Z(_01514_));
 MUX2_X1 _14957_ (.A(_07875_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][6] ),
    .S(_07982_),
    .Z(_01515_));
 MUX2_X1 _14958_ (.A(_07877_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][7] ),
    .S(_07982_),
    .Z(_01516_));
 MUX2_X1 _14959_ (.A(_07879_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][8] ),
    .S(_07982_),
    .Z(_01517_));
 MUX2_X1 _14960_ (.A(_07881_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][9] ),
    .S(_07982_),
    .Z(_01518_));
 NAND2_X1 _14961_ (.A1(_07895_),
    .A2(_07972_),
    .ZN(_07989_));
 BUF_X4 _14962_ (.A(_07989_),
    .Z(_07990_));
 CLKBUF_X3 _14963_ (.A(_07990_),
    .Z(_07991_));
 MUX2_X1 _14964_ (.A(_07744_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][0] ),
    .S(_07991_),
    .Z(_01519_));
 MUX2_X1 _14965_ (.A(_07752_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][10] ),
    .S(_07991_),
    .Z(_01520_));
 MUX2_X1 _14966_ (.A(_07754_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][11] ),
    .S(_07991_),
    .Z(_01521_));
 MUX2_X1 _14967_ (.A(_07756_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][12] ),
    .S(_07991_),
    .Z(_01522_));
 MUX2_X1 _14968_ (.A(_07758_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][13] ),
    .S(_07991_),
    .Z(_01523_));
 MUX2_X1 _14969_ (.A(_07760_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][14] ),
    .S(_07991_),
    .Z(_01524_));
 MUX2_X1 _14970_ (.A(_07762_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][15] ),
    .S(_07991_),
    .Z(_01525_));
 MUX2_X1 _14971_ (.A(_07764_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][16] ),
    .S(_07991_),
    .Z(_01526_));
 MUX2_X1 _14972_ (.A(_07766_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][17] ),
    .S(_07991_),
    .Z(_01527_));
 MUX2_X1 _14973_ (.A(_07768_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][18] ),
    .S(_07991_),
    .Z(_01528_));
 BUF_X4 _14974_ (.A(_07990_),
    .Z(_07992_));
 MUX2_X1 _14975_ (.A(_07770_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][19] ),
    .S(_07992_),
    .Z(_01529_));
 MUX2_X1 _14976_ (.A(_07773_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][1] ),
    .S(_07992_),
    .Z(_01530_));
 MUX2_X1 _14977_ (.A(_07775_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][20] ),
    .S(_07992_),
    .Z(_01531_));
 MUX2_X1 _14978_ (.A(_07777_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][21] ),
    .S(_07992_),
    .Z(_01532_));
 MUX2_X1 _14979_ (.A(_07779_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][22] ),
    .S(_07992_),
    .Z(_01533_));
 MUX2_X1 _14980_ (.A(_07781_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][23] ),
    .S(_07992_),
    .Z(_01534_));
 MUX2_X1 _14981_ (.A(_07783_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][24] ),
    .S(_07992_),
    .Z(_01535_));
 MUX2_X1 _14982_ (.A(_07785_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][25] ),
    .S(_07992_),
    .Z(_01536_));
 MUX2_X1 _14983_ (.A(_07787_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][26] ),
    .S(_07992_),
    .Z(_01537_));
 MUX2_X1 _14984_ (.A(_07789_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][27] ),
    .S(_07992_),
    .Z(_01538_));
 BUF_X4 _14985_ (.A(_07990_),
    .Z(_02296_));
 MUX2_X1 _14986_ (.A(_07791_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][28] ),
    .S(_02296_),
    .Z(_01539_));
 MUX2_X1 _14987_ (.A(_07794_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][29] ),
    .S(_02296_),
    .Z(_01540_));
 MUX2_X1 _14988_ (.A(_07796_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][2] ),
    .S(_02296_),
    .Z(_01541_));
 MUX2_X1 _14989_ (.A(_07798_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][30] ),
    .S(_02296_),
    .Z(_01542_));
 MUX2_X1 _14990_ (.A(_07800_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][31] ),
    .S(_02296_),
    .Z(_01543_));
 MUX2_X1 _14991_ (.A(_07802_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][32] ),
    .S(_02296_),
    .Z(_01544_));
 MUX2_X1 _14992_ (.A(_07804_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][33] ),
    .S(_02296_),
    .Z(_01545_));
 MUX2_X1 _14993_ (.A(_07806_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][34] ),
    .S(_02296_),
    .Z(_01546_));
 MUX2_X1 _14994_ (.A(_07808_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][35] ),
    .S(_02296_),
    .Z(_01547_));
 MUX2_X1 _14995_ (.A(_07810_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][36] ),
    .S(_02296_),
    .Z(_01548_));
 BUF_X4 _14996_ (.A(_07990_),
    .Z(_02297_));
 MUX2_X1 _14997_ (.A(_07812_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][37] ),
    .S(_02297_),
    .Z(_01549_));
 MUX2_X1 _14998_ (.A(_07815_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][38] ),
    .S(_02297_),
    .Z(_01550_));
 MUX2_X1 _14999_ (.A(_07817_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][39] ),
    .S(_02297_),
    .Z(_01551_));
 MUX2_X1 _15000_ (.A(_07819_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][3] ),
    .S(_02297_),
    .Z(_01552_));
 MUX2_X1 _15001_ (.A(_07821_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][40] ),
    .S(_02297_),
    .Z(_01553_));
 MUX2_X1 _15002_ (.A(_07823_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][41] ),
    .S(_02297_),
    .Z(_01554_));
 MUX2_X1 _15003_ (.A(_07825_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][42] ),
    .S(_02297_),
    .Z(_01555_));
 MUX2_X1 _15004_ (.A(_07827_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][43] ),
    .S(_02297_),
    .Z(_01556_));
 MUX2_X1 _15005_ (.A(_07829_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][44] ),
    .S(_02297_),
    .Z(_01557_));
 MUX2_X1 _15006_ (.A(_07831_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][45] ),
    .S(_02297_),
    .Z(_01558_));
 BUF_X4 _15007_ (.A(_07990_),
    .Z(_02298_));
 MUX2_X1 _15008_ (.A(_07833_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][46] ),
    .S(_02298_),
    .Z(_01559_));
 MUX2_X1 _15009_ (.A(_07836_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][47] ),
    .S(_02298_),
    .Z(_01560_));
 MUX2_X1 _15010_ (.A(_07838_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][48] ),
    .S(_02298_),
    .Z(_01561_));
 MUX2_X1 _15011_ (.A(_07840_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][49] ),
    .S(_02298_),
    .Z(_01562_));
 MUX2_X1 _15012_ (.A(_07842_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][4] ),
    .S(_02298_),
    .Z(_01563_));
 MUX2_X1 _15013_ (.A(_07844_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][50] ),
    .S(_02298_),
    .Z(_01564_));
 MUX2_X1 _15014_ (.A(_07846_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][51] ),
    .S(_02298_),
    .Z(_01565_));
 MUX2_X1 _15015_ (.A(_07848_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][52] ),
    .S(_02298_),
    .Z(_01566_));
 MUX2_X1 _15016_ (.A(_07850_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][53] ),
    .S(_02298_),
    .Z(_01567_));
 MUX2_X1 _15017_ (.A(_07852_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][54] ),
    .S(_02298_),
    .Z(_01568_));
 BUF_X4 _15018_ (.A(_07990_),
    .Z(_02299_));
 MUX2_X1 _15019_ (.A(_07854_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][55] ),
    .S(_02299_),
    .Z(_01569_));
 MUX2_X1 _15020_ (.A(_07857_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][56] ),
    .S(_02299_),
    .Z(_01570_));
 MUX2_X1 _15021_ (.A(_07859_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][57] ),
    .S(_02299_),
    .Z(_01571_));
 MUX2_X1 _15022_ (.A(_07861_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][58] ),
    .S(_02299_),
    .Z(_01572_));
 MUX2_X1 _15023_ (.A(_07863_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][59] ),
    .S(_02299_),
    .Z(_01573_));
 MUX2_X1 _15024_ (.A(_07865_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][5] ),
    .S(_02299_),
    .Z(_01574_));
 MUX2_X1 _15025_ (.A(_07867_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][60] ),
    .S(_02299_),
    .Z(_01575_));
 MUX2_X1 _15026_ (.A(_07869_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][61] ),
    .S(_02299_),
    .Z(_01576_));
 MUX2_X1 _15027_ (.A(_07871_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][62] ),
    .S(_02299_),
    .Z(_01577_));
 MUX2_X1 _15028_ (.A(_07873_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][63] ),
    .S(_02299_),
    .Z(_01578_));
 MUX2_X1 _15029_ (.A(_07875_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][6] ),
    .S(_07990_),
    .Z(_01579_));
 MUX2_X1 _15030_ (.A(_07877_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][7] ),
    .S(_07990_),
    .Z(_01580_));
 MUX2_X1 _15031_ (.A(_07879_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][8] ),
    .S(_07990_),
    .Z(_01581_));
 MUX2_X1 _15032_ (.A(_07881_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][9] ),
    .S(_07990_),
    .Z(_01582_));
 NOR3_X1 _15033_ (.A1(_07747_),
    .A2(_07748_),
    .A3(_07885_),
    .ZN(_02300_));
 BUF_X4 _15034_ (.A(_02300_),
    .Z(_02301_));
 CLKBUF_X3 _15035_ (.A(_02301_),
    .Z(_02302_));
 MUX2_X1 _15036_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][0] ),
    .B(_07745_),
    .S(_02302_),
    .Z(_01583_));
 MUX2_X1 _15037_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][10] ),
    .B(_07753_),
    .S(_02302_),
    .Z(_01584_));
 MUX2_X1 _15038_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][11] ),
    .B(_07755_),
    .S(_02302_),
    .Z(_01585_));
 MUX2_X1 _15039_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][12] ),
    .B(_07757_),
    .S(_02302_),
    .Z(_01586_));
 MUX2_X1 _15040_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][13] ),
    .B(_07759_),
    .S(_02302_),
    .Z(_01587_));
 MUX2_X1 _15041_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][14] ),
    .B(_07761_),
    .S(_02302_),
    .Z(_01588_));
 MUX2_X1 _15042_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][15] ),
    .B(_07763_),
    .S(_02302_),
    .Z(_01589_));
 MUX2_X1 _15043_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][16] ),
    .B(_07765_),
    .S(_02302_),
    .Z(_01590_));
 MUX2_X1 _15044_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][17] ),
    .B(_07767_),
    .S(_02302_),
    .Z(_01591_));
 MUX2_X1 _15045_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][18] ),
    .B(_07769_),
    .S(_02302_),
    .Z(_01592_));
 BUF_X4 _15046_ (.A(_02301_),
    .Z(_02303_));
 MUX2_X1 _15047_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][19] ),
    .B(_07771_),
    .S(_02303_),
    .Z(_01593_));
 MUX2_X1 _15048_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][1] ),
    .B(_07774_),
    .S(_02303_),
    .Z(_01594_));
 MUX2_X1 _15049_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][20] ),
    .B(_07776_),
    .S(_02303_),
    .Z(_01595_));
 MUX2_X1 _15050_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][21] ),
    .B(_07778_),
    .S(_02303_),
    .Z(_01596_));
 MUX2_X1 _15051_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][22] ),
    .B(_07780_),
    .S(_02303_),
    .Z(_01597_));
 MUX2_X1 _15052_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][23] ),
    .B(_07782_),
    .S(_02303_),
    .Z(_01598_));
 MUX2_X1 _15053_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][24] ),
    .B(_07784_),
    .S(_02303_),
    .Z(_01599_));
 MUX2_X1 _15054_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][25] ),
    .B(_07786_),
    .S(_02303_),
    .Z(_01600_));
 MUX2_X1 _15055_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][26] ),
    .B(_07788_),
    .S(_02303_),
    .Z(_01601_));
 MUX2_X1 _15056_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][27] ),
    .B(_07790_),
    .S(_02303_),
    .Z(_01602_));
 BUF_X4 _15057_ (.A(_02301_),
    .Z(_02304_));
 MUX2_X1 _15058_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][28] ),
    .B(_07792_),
    .S(_02304_),
    .Z(_01603_));
 MUX2_X1 _15059_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][29] ),
    .B(_07795_),
    .S(_02304_),
    .Z(_01604_));
 MUX2_X1 _15060_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][2] ),
    .B(_07797_),
    .S(_02304_),
    .Z(_01605_));
 MUX2_X1 _15061_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][30] ),
    .B(_07799_),
    .S(_02304_),
    .Z(_01606_));
 MUX2_X1 _15062_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][31] ),
    .B(_07801_),
    .S(_02304_),
    .Z(_01607_));
 MUX2_X1 _15063_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][32] ),
    .B(_07803_),
    .S(_02304_),
    .Z(_01608_));
 MUX2_X1 _15064_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][33] ),
    .B(_07805_),
    .S(_02304_),
    .Z(_01609_));
 MUX2_X1 _15065_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][34] ),
    .B(_07807_),
    .S(_02304_),
    .Z(_01610_));
 MUX2_X1 _15066_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][35] ),
    .B(_07809_),
    .S(_02304_),
    .Z(_01611_));
 MUX2_X1 _15067_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][36] ),
    .B(_07811_),
    .S(_02304_),
    .Z(_01612_));
 BUF_X4 _15068_ (.A(_02301_),
    .Z(_02305_));
 MUX2_X1 _15069_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][37] ),
    .B(_07813_),
    .S(_02305_),
    .Z(_01613_));
 MUX2_X1 _15070_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][38] ),
    .B(_07816_),
    .S(_02305_),
    .Z(_01614_));
 MUX2_X1 _15071_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][39] ),
    .B(_07818_),
    .S(_02305_),
    .Z(_01615_));
 MUX2_X1 _15072_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][3] ),
    .B(_07820_),
    .S(_02305_),
    .Z(_01616_));
 MUX2_X1 _15073_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][40] ),
    .B(_07822_),
    .S(_02305_),
    .Z(_01617_));
 MUX2_X1 _15074_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][41] ),
    .B(_07824_),
    .S(_02305_),
    .Z(_01618_));
 MUX2_X1 _15075_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][42] ),
    .B(_07826_),
    .S(_02305_),
    .Z(_01619_));
 MUX2_X1 _15076_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][43] ),
    .B(_07828_),
    .S(_02305_),
    .Z(_01620_));
 MUX2_X1 _15077_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][44] ),
    .B(_07830_),
    .S(_02305_),
    .Z(_01621_));
 MUX2_X1 _15078_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][45] ),
    .B(_07832_),
    .S(_02305_),
    .Z(_01622_));
 BUF_X4 _15079_ (.A(_02301_),
    .Z(_02306_));
 MUX2_X1 _15080_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][46] ),
    .B(_07834_),
    .S(_02306_),
    .Z(_01623_));
 MUX2_X1 _15081_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][47] ),
    .B(_07837_),
    .S(_02306_),
    .Z(_01624_));
 MUX2_X1 _15082_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][48] ),
    .B(_07839_),
    .S(_02306_),
    .Z(_01625_));
 MUX2_X1 _15083_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][49] ),
    .B(_07841_),
    .S(_02306_),
    .Z(_01626_));
 MUX2_X1 _15084_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][4] ),
    .B(_07843_),
    .S(_02306_),
    .Z(_01627_));
 MUX2_X1 _15085_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][50] ),
    .B(_07845_),
    .S(_02306_),
    .Z(_01628_));
 MUX2_X1 _15086_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][51] ),
    .B(_07847_),
    .S(_02306_),
    .Z(_01629_));
 MUX2_X1 _15087_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][52] ),
    .B(_07849_),
    .S(_02306_),
    .Z(_01630_));
 MUX2_X1 _15088_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][53] ),
    .B(_07851_),
    .S(_02306_),
    .Z(_01631_));
 MUX2_X1 _15089_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][54] ),
    .B(_07853_),
    .S(_02306_),
    .Z(_01632_));
 BUF_X4 _15090_ (.A(_02301_),
    .Z(_02307_));
 MUX2_X1 _15091_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][55] ),
    .B(_07855_),
    .S(_02307_),
    .Z(_01633_));
 MUX2_X1 _15092_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][56] ),
    .B(_07858_),
    .S(_02307_),
    .Z(_01634_));
 MUX2_X1 _15093_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][57] ),
    .B(_07860_),
    .S(_02307_),
    .Z(_01635_));
 MUX2_X1 _15094_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][58] ),
    .B(_07862_),
    .S(_02307_),
    .Z(_01636_));
 MUX2_X1 _15095_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][59] ),
    .B(_07864_),
    .S(_02307_),
    .Z(_01637_));
 MUX2_X1 _15096_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][5] ),
    .B(_07866_),
    .S(_02307_),
    .Z(_01638_));
 MUX2_X1 _15097_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][60] ),
    .B(_07868_),
    .S(_02307_),
    .Z(_01639_));
 MUX2_X1 _15098_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][61] ),
    .B(_07870_),
    .S(_02307_),
    .Z(_01640_));
 MUX2_X1 _15099_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][62] ),
    .B(_07872_),
    .S(_02307_),
    .Z(_01641_));
 MUX2_X1 _15100_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][63] ),
    .B(_07874_),
    .S(_02307_),
    .Z(_01642_));
 MUX2_X1 _15101_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][6] ),
    .B(_07876_),
    .S(_02301_),
    .Z(_01643_));
 MUX2_X1 _15102_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][7] ),
    .B(_07878_),
    .S(_02301_),
    .Z(_01644_));
 MUX2_X1 _15103_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][8] ),
    .B(_07880_),
    .S(_02301_),
    .Z(_01645_));
 MUX2_X1 _15104_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][9] ),
    .B(_07882_),
    .S(_02301_),
    .Z(_01646_));
 NAND2_X1 _15105_ (.A1(_10597_),
    .A2(_07886_),
    .ZN(_02308_));
 BUF_X4 _15106_ (.A(_02308_),
    .Z(_02309_));
 CLKBUF_X3 _15107_ (.A(_02309_),
    .Z(_02310_));
 MUX2_X1 _15108_ (.A(_07744_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][0] ),
    .S(_02310_),
    .Z(_01647_));
 MUX2_X1 _15109_ (.A(_07752_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][10] ),
    .S(_02310_),
    .Z(_01648_));
 MUX2_X1 _15110_ (.A(_07754_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][11] ),
    .S(_02310_),
    .Z(_01649_));
 MUX2_X1 _15111_ (.A(_07756_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][12] ),
    .S(_02310_),
    .Z(_01650_));
 MUX2_X1 _15112_ (.A(_07758_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][13] ),
    .S(_02310_),
    .Z(_01651_));
 MUX2_X1 _15113_ (.A(_07760_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][14] ),
    .S(_02310_),
    .Z(_01652_));
 MUX2_X1 _15114_ (.A(_07762_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][15] ),
    .S(_02310_),
    .Z(_01653_));
 MUX2_X1 _15115_ (.A(_07764_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][16] ),
    .S(_02310_),
    .Z(_01654_));
 MUX2_X1 _15116_ (.A(_07766_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][17] ),
    .S(_02310_),
    .Z(_01655_));
 MUX2_X1 _15117_ (.A(_07768_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][18] ),
    .S(_02310_),
    .Z(_01656_));
 BUF_X4 _15118_ (.A(_02309_),
    .Z(_02311_));
 MUX2_X1 _15119_ (.A(_07770_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][19] ),
    .S(_02311_),
    .Z(_01657_));
 MUX2_X1 _15120_ (.A(_07773_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][1] ),
    .S(_02311_),
    .Z(_01658_));
 MUX2_X1 _15121_ (.A(_07775_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][20] ),
    .S(_02311_),
    .Z(_01659_));
 MUX2_X1 _15122_ (.A(_07777_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][21] ),
    .S(_02311_),
    .Z(_01660_));
 MUX2_X1 _15123_ (.A(_07779_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][22] ),
    .S(_02311_),
    .Z(_01661_));
 MUX2_X1 _15124_ (.A(_07781_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][23] ),
    .S(_02311_),
    .Z(_01662_));
 MUX2_X1 _15125_ (.A(_07783_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][24] ),
    .S(_02311_),
    .Z(_01663_));
 MUX2_X1 _15126_ (.A(_07785_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][25] ),
    .S(_02311_),
    .Z(_01664_));
 MUX2_X1 _15127_ (.A(_07787_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][26] ),
    .S(_02311_),
    .Z(_01665_));
 MUX2_X1 _15128_ (.A(_07789_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][27] ),
    .S(_02311_),
    .Z(_01666_));
 BUF_X4 _15129_ (.A(_02309_),
    .Z(_02312_));
 MUX2_X1 _15130_ (.A(_07791_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][28] ),
    .S(_02312_),
    .Z(_01667_));
 MUX2_X1 _15131_ (.A(_07794_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][29] ),
    .S(_02312_),
    .Z(_01668_));
 MUX2_X1 _15132_ (.A(_07796_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][2] ),
    .S(_02312_),
    .Z(_01669_));
 MUX2_X1 _15133_ (.A(_07798_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][30] ),
    .S(_02312_),
    .Z(_01670_));
 MUX2_X1 _15134_ (.A(_07800_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][31] ),
    .S(_02312_),
    .Z(_01671_));
 MUX2_X1 _15135_ (.A(_07802_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][32] ),
    .S(_02312_),
    .Z(_01672_));
 MUX2_X1 _15136_ (.A(_07804_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][33] ),
    .S(_02312_),
    .Z(_01673_));
 MUX2_X1 _15137_ (.A(_07806_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][34] ),
    .S(_02312_),
    .Z(_01674_));
 MUX2_X1 _15138_ (.A(_07808_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][35] ),
    .S(_02312_),
    .Z(_01675_));
 MUX2_X1 _15139_ (.A(_07810_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][36] ),
    .S(_02312_),
    .Z(_01676_));
 BUF_X4 _15140_ (.A(_02309_),
    .Z(_02313_));
 MUX2_X1 _15141_ (.A(_07812_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][37] ),
    .S(_02313_),
    .Z(_01677_));
 MUX2_X1 _15142_ (.A(_07815_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][38] ),
    .S(_02313_),
    .Z(_01678_));
 MUX2_X1 _15143_ (.A(_07817_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][39] ),
    .S(_02313_),
    .Z(_01679_));
 MUX2_X1 _15144_ (.A(_07819_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][3] ),
    .S(_02313_),
    .Z(_01680_));
 MUX2_X1 _15145_ (.A(_07821_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][40] ),
    .S(_02313_),
    .Z(_01681_));
 MUX2_X1 _15146_ (.A(_07823_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][41] ),
    .S(_02313_),
    .Z(_01682_));
 MUX2_X1 _15147_ (.A(_07825_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][42] ),
    .S(_02313_),
    .Z(_01683_));
 MUX2_X1 _15148_ (.A(_07827_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][43] ),
    .S(_02313_),
    .Z(_01684_));
 MUX2_X1 _15149_ (.A(_07829_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][44] ),
    .S(_02313_),
    .Z(_01685_));
 MUX2_X1 _15150_ (.A(_07831_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][45] ),
    .S(_02313_),
    .Z(_01686_));
 BUF_X4 _15151_ (.A(_02309_),
    .Z(_02314_));
 MUX2_X1 _15152_ (.A(_07833_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][46] ),
    .S(_02314_),
    .Z(_01687_));
 MUX2_X1 _15153_ (.A(_07836_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][47] ),
    .S(_02314_),
    .Z(_01688_));
 MUX2_X1 _15154_ (.A(_07838_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][48] ),
    .S(_02314_),
    .Z(_01689_));
 MUX2_X1 _15155_ (.A(_07840_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][49] ),
    .S(_02314_),
    .Z(_01690_));
 MUX2_X1 _15156_ (.A(_07842_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][4] ),
    .S(_02314_),
    .Z(_01691_));
 MUX2_X1 _15157_ (.A(_07844_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][50] ),
    .S(_02314_),
    .Z(_01692_));
 MUX2_X1 _15158_ (.A(_07846_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][51] ),
    .S(_02314_),
    .Z(_01693_));
 MUX2_X1 _15159_ (.A(_07848_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][52] ),
    .S(_02314_),
    .Z(_01694_));
 MUX2_X1 _15160_ (.A(_07850_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][53] ),
    .S(_02314_),
    .Z(_01695_));
 MUX2_X1 _15161_ (.A(_07852_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][54] ),
    .S(_02314_),
    .Z(_01696_));
 BUF_X4 _15162_ (.A(_02309_),
    .Z(_02315_));
 MUX2_X1 _15163_ (.A(_07854_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][55] ),
    .S(_02315_),
    .Z(_01697_));
 MUX2_X1 _15164_ (.A(_07857_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][56] ),
    .S(_02315_),
    .Z(_01698_));
 MUX2_X1 _15165_ (.A(_07859_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][57] ),
    .S(_02315_),
    .Z(_01699_));
 MUX2_X1 _15166_ (.A(_07861_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][58] ),
    .S(_02315_),
    .Z(_01700_));
 MUX2_X1 _15167_ (.A(_07863_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][59] ),
    .S(_02315_),
    .Z(_01701_));
 MUX2_X1 _15168_ (.A(_07865_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][5] ),
    .S(_02315_),
    .Z(_01702_));
 MUX2_X1 _15169_ (.A(_07867_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][60] ),
    .S(_02315_),
    .Z(_01703_));
 MUX2_X1 _15170_ (.A(_07869_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][61] ),
    .S(_02315_),
    .Z(_01704_));
 MUX2_X1 _15171_ (.A(_07871_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][62] ),
    .S(_02315_),
    .Z(_01705_));
 MUX2_X1 _15172_ (.A(_07873_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][63] ),
    .S(_02315_),
    .Z(_01706_));
 MUX2_X1 _15173_ (.A(_07875_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][6] ),
    .S(_02309_),
    .Z(_01707_));
 MUX2_X1 _15174_ (.A(_07877_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][7] ),
    .S(_02309_),
    .Z(_01708_));
 MUX2_X1 _15175_ (.A(_07879_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][8] ),
    .S(_02309_),
    .Z(_01709_));
 MUX2_X1 _15176_ (.A(_07881_),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[9][9] ),
    .S(_02309_),
    .Z(_01710_));
 NOR2_X4 _15177_ (.A1(_06540_),
    .A2(_10463_),
    .ZN(_02316_));
 NAND2_X1 _15178_ (.A1(_10602_),
    .A2(_02316_),
    .ZN(_02317_));
 BUF_X4 _15179_ (.A(_02317_),
    .Z(_02318_));
 CLKBUF_X3 _15180_ (.A(_02318_),
    .Z(_02319_));
 MUX2_X1 _15181_ (.A(net131),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][0] ),
    .S(_02319_),
    .Z(_01738_));
 MUX2_X1 _15182_ (.A(net132),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][10] ),
    .S(_02319_),
    .Z(_01739_));
 MUX2_X1 _15183_ (.A(net133),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][11] ),
    .S(_02319_),
    .Z(_01740_));
 MUX2_X1 _15184_ (.A(net134),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][12] ),
    .S(_02319_),
    .Z(_01741_));
 MUX2_X1 _15185_ (.A(net135),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][13] ),
    .S(_02319_),
    .Z(_01742_));
 MUX2_X1 _15186_ (.A(net136),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][14] ),
    .S(_02319_),
    .Z(_01743_));
 MUX2_X1 _15187_ (.A(net137),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][15] ),
    .S(_02319_),
    .Z(_01744_));
 MUX2_X1 _15188_ (.A(net138),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][16] ),
    .S(_02319_),
    .Z(_01745_));
 MUX2_X1 _15189_ (.A(net139),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][17] ),
    .S(_02319_),
    .Z(_01746_));
 MUX2_X1 _15190_ (.A(net140),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][18] ),
    .S(_02319_),
    .Z(_01747_));
 BUF_X4 _15191_ (.A(_02318_),
    .Z(_02320_));
 MUX2_X1 _15192_ (.A(net141),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][19] ),
    .S(_02320_),
    .Z(_01748_));
 MUX2_X1 _15193_ (.A(net142),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][1] ),
    .S(_02320_),
    .Z(_01749_));
 MUX2_X1 _15194_ (.A(net143),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][20] ),
    .S(_02320_),
    .Z(_01750_));
 MUX2_X1 _15195_ (.A(net144),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][21] ),
    .S(_02320_),
    .Z(_01751_));
 MUX2_X1 _15196_ (.A(net145),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][22] ),
    .S(_02320_),
    .Z(_01752_));
 MUX2_X1 _15197_ (.A(net146),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][23] ),
    .S(_02320_),
    .Z(_01753_));
 MUX2_X1 _15198_ (.A(net147),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][24] ),
    .S(_02320_),
    .Z(_01754_));
 MUX2_X1 _15199_ (.A(net148),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][25] ),
    .S(_02320_),
    .Z(_01755_));
 MUX2_X1 _15200_ (.A(net149),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][26] ),
    .S(_02320_),
    .Z(_01756_));
 MUX2_X1 _15201_ (.A(net150),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][27] ),
    .S(_02320_),
    .Z(_01757_));
 BUF_X4 _15202_ (.A(_02318_),
    .Z(_02321_));
 MUX2_X1 _15203_ (.A(net151),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][28] ),
    .S(_02321_),
    .Z(_01758_));
 MUX2_X1 _15204_ (.A(net152),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][29] ),
    .S(_02321_),
    .Z(_01759_));
 MUX2_X1 _15205_ (.A(net153),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][2] ),
    .S(_02321_),
    .Z(_01760_));
 MUX2_X1 _15206_ (.A(net154),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][30] ),
    .S(_02321_),
    .Z(_01761_));
 MUX2_X1 _15207_ (.A(net155),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][31] ),
    .S(_02321_),
    .Z(_01762_));
 MUX2_X1 _15208_ (.A(net156),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][32] ),
    .S(_02321_),
    .Z(_01763_));
 MUX2_X1 _15209_ (.A(net157),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][33] ),
    .S(_02321_),
    .Z(_01764_));
 MUX2_X1 _15210_ (.A(net158),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][34] ),
    .S(_02321_),
    .Z(_01765_));
 MUX2_X1 _15211_ (.A(net159),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][35] ),
    .S(_02321_),
    .Z(_01766_));
 MUX2_X1 _15212_ (.A(net160),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][36] ),
    .S(_02321_),
    .Z(_01767_));
 BUF_X4 _15213_ (.A(_02318_),
    .Z(_02322_));
 MUX2_X1 _15214_ (.A(net161),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][37] ),
    .S(_02322_),
    .Z(_01768_));
 MUX2_X1 _15215_ (.A(net162),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][38] ),
    .S(_02322_),
    .Z(_01769_));
 MUX2_X1 _15216_ (.A(net163),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][39] ),
    .S(_02322_),
    .Z(_01770_));
 MUX2_X1 _15217_ (.A(net164),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][3] ),
    .S(_02322_),
    .Z(_01771_));
 MUX2_X1 _15218_ (.A(net165),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][40] ),
    .S(_02322_),
    .Z(_01772_));
 MUX2_X1 _15219_ (.A(net166),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][41] ),
    .S(_02322_),
    .Z(_01773_));
 MUX2_X1 _15220_ (.A(net167),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][42] ),
    .S(_02322_),
    .Z(_01774_));
 MUX2_X1 _15221_ (.A(net168),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][43] ),
    .S(_02322_),
    .Z(_01775_));
 MUX2_X1 _15222_ (.A(net169),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][44] ),
    .S(_02322_),
    .Z(_01776_));
 MUX2_X1 _15223_ (.A(net170),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][45] ),
    .S(_02322_),
    .Z(_01777_));
 BUF_X4 _15224_ (.A(_02318_),
    .Z(_02323_));
 MUX2_X1 _15225_ (.A(net171),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][46] ),
    .S(_02323_),
    .Z(_01778_));
 MUX2_X1 _15226_ (.A(net172),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][47] ),
    .S(_02323_),
    .Z(_01779_));
 MUX2_X1 _15227_ (.A(net173),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][48] ),
    .S(_02323_),
    .Z(_01780_));
 MUX2_X1 _15228_ (.A(net174),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][49] ),
    .S(_02323_),
    .Z(_01781_));
 MUX2_X1 _15229_ (.A(net175),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][4] ),
    .S(_02323_),
    .Z(_01782_));
 MUX2_X1 _15230_ (.A(net176),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][50] ),
    .S(_02323_),
    .Z(_01783_));
 MUX2_X1 _15231_ (.A(net177),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][51] ),
    .S(_02323_),
    .Z(_01784_));
 MUX2_X1 _15232_ (.A(net178),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][52] ),
    .S(_02323_),
    .Z(_01785_));
 MUX2_X1 _15233_ (.A(net179),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][53] ),
    .S(_02323_),
    .Z(_01786_));
 MUX2_X1 _15234_ (.A(net180),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][54] ),
    .S(_02323_),
    .Z(_01787_));
 BUF_X4 _15235_ (.A(_02318_),
    .Z(_02324_));
 MUX2_X1 _15236_ (.A(net181),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][55] ),
    .S(_02324_),
    .Z(_01788_));
 MUX2_X1 _15237_ (.A(net182),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][56] ),
    .S(_02324_),
    .Z(_01789_));
 MUX2_X1 _15238_ (.A(net183),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][57] ),
    .S(_02324_),
    .Z(_01790_));
 MUX2_X1 _15239_ (.A(net184),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][58] ),
    .S(_02324_),
    .Z(_01791_));
 MUX2_X1 _15240_ (.A(net185),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][59] ),
    .S(_02324_),
    .Z(_01792_));
 MUX2_X1 _15241_ (.A(net186),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][5] ),
    .S(_02324_),
    .Z(_01793_));
 MUX2_X1 _15242_ (.A(net187),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][60] ),
    .S(_02324_),
    .Z(_01794_));
 MUX2_X1 _15243_ (.A(net188),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][61] ),
    .S(_02324_),
    .Z(_01795_));
 MUX2_X1 _15244_ (.A(net189),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][62] ),
    .S(_02324_),
    .Z(_01796_));
 MUX2_X1 _15245_ (.A(net190),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][63] ),
    .S(_02324_),
    .Z(_01797_));
 MUX2_X1 _15246_ (.A(net191),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][6] ),
    .S(_02318_),
    .Z(_01798_));
 MUX2_X1 _15247_ (.A(net192),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][7] ),
    .S(_02318_),
    .Z(_01799_));
 MUX2_X1 _15248_ (.A(net193),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][8] ),
    .S(_02318_),
    .Z(_01800_));
 MUX2_X1 _15249_ (.A(net194),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[0][9] ),
    .S(_02318_),
    .Z(_01801_));
 NAND2_X1 _15250_ (.A1(_10605_),
    .A2(_02316_),
    .ZN(_02325_));
 BUF_X4 _15251_ (.A(_02325_),
    .Z(_02326_));
 CLKBUF_X3 _15252_ (.A(_02326_),
    .Z(_02327_));
 MUX2_X1 _15253_ (.A(net131),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][0] ),
    .S(_02327_),
    .Z(_01802_));
 MUX2_X1 _15254_ (.A(net132),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][10] ),
    .S(_02327_),
    .Z(_01803_));
 MUX2_X1 _15255_ (.A(net133),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][11] ),
    .S(_02327_),
    .Z(_01804_));
 MUX2_X1 _15256_ (.A(net134),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][12] ),
    .S(_02327_),
    .Z(_01805_));
 MUX2_X1 _15257_ (.A(net135),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][13] ),
    .S(_02327_),
    .Z(_01806_));
 MUX2_X1 _15258_ (.A(net136),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][14] ),
    .S(_02327_),
    .Z(_01807_));
 MUX2_X1 _15259_ (.A(net137),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][15] ),
    .S(_02327_),
    .Z(_01808_));
 MUX2_X1 _15260_ (.A(net138),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][16] ),
    .S(_02327_),
    .Z(_01809_));
 MUX2_X1 _15261_ (.A(net139),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][17] ),
    .S(_02327_),
    .Z(_01810_));
 MUX2_X1 _15262_ (.A(net140),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][18] ),
    .S(_02327_),
    .Z(_01811_));
 CLKBUF_X3 _15263_ (.A(_02326_),
    .Z(_02328_));
 MUX2_X1 _15264_ (.A(net141),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][19] ),
    .S(_02328_),
    .Z(_01812_));
 MUX2_X1 _15265_ (.A(net142),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][1] ),
    .S(_02328_),
    .Z(_01813_));
 MUX2_X1 _15266_ (.A(net143),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][20] ),
    .S(_02328_),
    .Z(_01814_));
 MUX2_X1 _15267_ (.A(net144),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][21] ),
    .S(_02328_),
    .Z(_01815_));
 MUX2_X1 _15268_ (.A(net145),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][22] ),
    .S(_02328_),
    .Z(_01816_));
 MUX2_X1 _15269_ (.A(net146),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][23] ),
    .S(_02328_),
    .Z(_01817_));
 MUX2_X1 _15270_ (.A(net147),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][24] ),
    .S(_02328_),
    .Z(_01818_));
 MUX2_X1 _15271_ (.A(net148),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][25] ),
    .S(_02328_),
    .Z(_01819_));
 MUX2_X1 _15272_ (.A(net149),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][26] ),
    .S(_02328_),
    .Z(_01820_));
 MUX2_X1 _15273_ (.A(net150),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][27] ),
    .S(_02328_),
    .Z(_01821_));
 BUF_X4 _15274_ (.A(_02326_),
    .Z(_02329_));
 MUX2_X1 _15275_ (.A(net151),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][28] ),
    .S(_02329_),
    .Z(_01822_));
 MUX2_X1 _15276_ (.A(net152),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][29] ),
    .S(_02329_),
    .Z(_01823_));
 MUX2_X1 _15277_ (.A(net153),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][2] ),
    .S(_02329_),
    .Z(_01824_));
 MUX2_X1 _15278_ (.A(net154),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][30] ),
    .S(_02329_),
    .Z(_01825_));
 MUX2_X1 _15279_ (.A(net155),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][31] ),
    .S(_02329_),
    .Z(_01826_));
 MUX2_X1 _15280_ (.A(net156),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][32] ),
    .S(_02329_),
    .Z(_01827_));
 MUX2_X1 _15281_ (.A(net157),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][33] ),
    .S(_02329_),
    .Z(_01828_));
 MUX2_X1 _15282_ (.A(net158),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][34] ),
    .S(_02329_),
    .Z(_01829_));
 MUX2_X1 _15283_ (.A(net159),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][35] ),
    .S(_02329_),
    .Z(_01830_));
 MUX2_X1 _15284_ (.A(net160),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][36] ),
    .S(_02329_),
    .Z(_01831_));
 BUF_X4 _15285_ (.A(_02326_),
    .Z(_02330_));
 MUX2_X1 _15286_ (.A(net161),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][37] ),
    .S(_02330_),
    .Z(_01832_));
 MUX2_X1 _15287_ (.A(net162),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][38] ),
    .S(_02330_),
    .Z(_01833_));
 MUX2_X1 _15288_ (.A(net163),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][39] ),
    .S(_02330_),
    .Z(_01834_));
 MUX2_X1 _15289_ (.A(net164),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][3] ),
    .S(_02330_),
    .Z(_01835_));
 MUX2_X1 _15290_ (.A(net165),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][40] ),
    .S(_02330_),
    .Z(_01836_));
 MUX2_X1 _15291_ (.A(net166),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][41] ),
    .S(_02330_),
    .Z(_01837_));
 MUX2_X1 _15292_ (.A(net167),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][42] ),
    .S(_02330_),
    .Z(_01838_));
 MUX2_X1 _15293_ (.A(net168),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][43] ),
    .S(_02330_),
    .Z(_01839_));
 MUX2_X1 _15294_ (.A(net169),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][44] ),
    .S(_02330_),
    .Z(_01840_));
 MUX2_X1 _15295_ (.A(net170),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][45] ),
    .S(_02330_),
    .Z(_01841_));
 BUF_X4 _15296_ (.A(_02326_),
    .Z(_02331_));
 MUX2_X1 _15297_ (.A(net171),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][46] ),
    .S(_02331_),
    .Z(_01842_));
 MUX2_X1 _15298_ (.A(net172),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][47] ),
    .S(_02331_),
    .Z(_01843_));
 MUX2_X1 _15299_ (.A(net173),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][48] ),
    .S(_02331_),
    .Z(_01844_));
 MUX2_X1 _15300_ (.A(net174),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][49] ),
    .S(_02331_),
    .Z(_01845_));
 MUX2_X1 _15301_ (.A(net175),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][4] ),
    .S(_02331_),
    .Z(_01846_));
 MUX2_X1 _15302_ (.A(net176),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][50] ),
    .S(_02331_),
    .Z(_01847_));
 MUX2_X1 _15303_ (.A(net177),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][51] ),
    .S(_02331_),
    .Z(_01848_));
 MUX2_X1 _15304_ (.A(net178),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][52] ),
    .S(_02331_),
    .Z(_01849_));
 MUX2_X1 _15305_ (.A(net179),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][53] ),
    .S(_02331_),
    .Z(_01850_));
 MUX2_X1 _15306_ (.A(net180),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][54] ),
    .S(_02331_),
    .Z(_01851_));
 BUF_X4 _15307_ (.A(_02326_),
    .Z(_02332_));
 MUX2_X1 _15308_ (.A(net181),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][55] ),
    .S(_02332_),
    .Z(_01852_));
 MUX2_X1 _15309_ (.A(net182),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][56] ),
    .S(_02332_),
    .Z(_01853_));
 MUX2_X1 _15310_ (.A(net183),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][57] ),
    .S(_02332_),
    .Z(_01854_));
 MUX2_X1 _15311_ (.A(net184),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][58] ),
    .S(_02332_),
    .Z(_01855_));
 MUX2_X1 _15312_ (.A(net185),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][59] ),
    .S(_02332_),
    .Z(_01856_));
 MUX2_X1 _15313_ (.A(net186),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][5] ),
    .S(_02332_),
    .Z(_01857_));
 MUX2_X1 _15314_ (.A(net187),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][60] ),
    .S(_02332_),
    .Z(_01858_));
 MUX2_X1 _15315_ (.A(net188),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][61] ),
    .S(_02332_),
    .Z(_01859_));
 MUX2_X1 _15316_ (.A(net189),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][62] ),
    .S(_02332_),
    .Z(_01860_));
 MUX2_X1 _15317_ (.A(net190),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][63] ),
    .S(_02332_),
    .Z(_01861_));
 MUX2_X1 _15318_ (.A(net191),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][6] ),
    .S(_02326_),
    .Z(_01862_));
 MUX2_X1 _15319_ (.A(net192),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][7] ),
    .S(_02326_),
    .Z(_01863_));
 MUX2_X1 _15320_ (.A(net193),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][8] ),
    .S(_02326_),
    .Z(_01864_));
 MUX2_X1 _15321_ (.A(net194),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[1][9] ),
    .S(_02326_),
    .Z(_01865_));
 NAND2_X1 _15322_ (.A1(_10603_),
    .A2(_02316_),
    .ZN(_02333_));
 BUF_X4 _15323_ (.A(_02333_),
    .Z(_02334_));
 CLKBUF_X3 _15324_ (.A(_02334_),
    .Z(_02335_));
 MUX2_X1 _15325_ (.A(net131),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][0] ),
    .S(_02335_),
    .Z(_01866_));
 MUX2_X1 _15326_ (.A(net132),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][10] ),
    .S(_02335_),
    .Z(_01867_));
 MUX2_X1 _15327_ (.A(net133),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][11] ),
    .S(_02335_),
    .Z(_01868_));
 MUX2_X1 _15328_ (.A(net134),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][12] ),
    .S(_02335_),
    .Z(_01869_));
 MUX2_X1 _15329_ (.A(net135),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][13] ),
    .S(_02335_),
    .Z(_01870_));
 MUX2_X1 _15330_ (.A(net136),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][14] ),
    .S(_02335_),
    .Z(_01871_));
 MUX2_X1 _15331_ (.A(net137),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][15] ),
    .S(_02335_),
    .Z(_01872_));
 MUX2_X1 _15332_ (.A(net138),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][16] ),
    .S(_02335_),
    .Z(_01873_));
 MUX2_X1 _15333_ (.A(net139),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][17] ),
    .S(_02335_),
    .Z(_01874_));
 MUX2_X1 _15334_ (.A(net140),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][18] ),
    .S(_02335_),
    .Z(_01875_));
 BUF_X4 _15335_ (.A(_02334_),
    .Z(_02336_));
 MUX2_X1 _15336_ (.A(net141),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][19] ),
    .S(_02336_),
    .Z(_01876_));
 MUX2_X1 _15337_ (.A(net142),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][1] ),
    .S(_02336_),
    .Z(_01877_));
 MUX2_X1 _15338_ (.A(net143),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][20] ),
    .S(_02336_),
    .Z(_01878_));
 MUX2_X1 _15339_ (.A(net144),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][21] ),
    .S(_02336_),
    .Z(_01879_));
 MUX2_X1 _15340_ (.A(net145),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][22] ),
    .S(_02336_),
    .Z(_01880_));
 MUX2_X1 _15341_ (.A(net146),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][23] ),
    .S(_02336_),
    .Z(_01881_));
 MUX2_X1 _15342_ (.A(net147),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][24] ),
    .S(_02336_),
    .Z(_01882_));
 MUX2_X1 _15343_ (.A(net148),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][25] ),
    .S(_02336_),
    .Z(_01883_));
 MUX2_X1 _15344_ (.A(net149),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][26] ),
    .S(_02336_),
    .Z(_01884_));
 MUX2_X1 _15345_ (.A(net150),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][27] ),
    .S(_02336_),
    .Z(_01885_));
 BUF_X4 _15346_ (.A(_02334_),
    .Z(_02337_));
 MUX2_X1 _15347_ (.A(net151),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][28] ),
    .S(_02337_),
    .Z(_01886_));
 MUX2_X1 _15348_ (.A(net152),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][29] ),
    .S(_02337_),
    .Z(_01887_));
 MUX2_X1 _15349_ (.A(net153),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][2] ),
    .S(_02337_),
    .Z(_01888_));
 MUX2_X1 _15350_ (.A(net154),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][30] ),
    .S(_02337_),
    .Z(_01889_));
 MUX2_X1 _15351_ (.A(net155),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][31] ),
    .S(_02337_),
    .Z(_01890_));
 MUX2_X1 _15352_ (.A(net156),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][32] ),
    .S(_02337_),
    .Z(_01891_));
 MUX2_X1 _15353_ (.A(net157),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][33] ),
    .S(_02337_),
    .Z(_01892_));
 MUX2_X1 _15354_ (.A(net158),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][34] ),
    .S(_02337_),
    .Z(_01893_));
 MUX2_X1 _15355_ (.A(net159),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][35] ),
    .S(_02337_),
    .Z(_01894_));
 MUX2_X1 _15356_ (.A(net160),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][36] ),
    .S(_02337_),
    .Z(_01895_));
 BUF_X4 _15357_ (.A(_02334_),
    .Z(_02338_));
 MUX2_X1 _15358_ (.A(net161),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][37] ),
    .S(_02338_),
    .Z(_01896_));
 MUX2_X1 _15359_ (.A(net162),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][38] ),
    .S(_02338_),
    .Z(_01897_));
 MUX2_X1 _15360_ (.A(net163),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][39] ),
    .S(_02338_),
    .Z(_01898_));
 MUX2_X1 _15361_ (.A(net164),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][3] ),
    .S(_02338_),
    .Z(_01899_));
 MUX2_X1 _15362_ (.A(net165),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][40] ),
    .S(_02338_),
    .Z(_01900_));
 MUX2_X1 _15363_ (.A(net166),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][41] ),
    .S(_02338_),
    .Z(_01901_));
 MUX2_X1 _15364_ (.A(net167),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][42] ),
    .S(_02338_),
    .Z(_01902_));
 MUX2_X1 _15365_ (.A(net168),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][43] ),
    .S(_02338_),
    .Z(_01903_));
 MUX2_X1 _15366_ (.A(net169),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][44] ),
    .S(_02338_),
    .Z(_01904_));
 MUX2_X1 _15367_ (.A(net170),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][45] ),
    .S(_02338_),
    .Z(_01905_));
 BUF_X4 _15368_ (.A(_02334_),
    .Z(_02339_));
 MUX2_X1 _15369_ (.A(net171),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][46] ),
    .S(_02339_),
    .Z(_01906_));
 MUX2_X1 _15370_ (.A(net172),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][47] ),
    .S(_02339_),
    .Z(_01907_));
 MUX2_X1 _15371_ (.A(net173),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][48] ),
    .S(_02339_),
    .Z(_01908_));
 MUX2_X1 _15372_ (.A(net174),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][49] ),
    .S(_02339_),
    .Z(_01909_));
 MUX2_X1 _15373_ (.A(net175),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][4] ),
    .S(_02339_),
    .Z(_01910_));
 MUX2_X1 _15374_ (.A(net176),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][50] ),
    .S(_02339_),
    .Z(_01911_));
 MUX2_X1 _15375_ (.A(net177),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][51] ),
    .S(_02339_),
    .Z(_01912_));
 MUX2_X1 _15376_ (.A(net178),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][52] ),
    .S(_02339_),
    .Z(_01913_));
 MUX2_X1 _15377_ (.A(net179),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][53] ),
    .S(_02339_),
    .Z(_01914_));
 MUX2_X1 _15378_ (.A(net180),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][54] ),
    .S(_02339_),
    .Z(_01915_));
 BUF_X4 _15379_ (.A(_02334_),
    .Z(_02340_));
 MUX2_X1 _15380_ (.A(net181),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][55] ),
    .S(_02340_),
    .Z(_01916_));
 MUX2_X1 _15381_ (.A(net182),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][56] ),
    .S(_02340_),
    .Z(_01917_));
 MUX2_X1 _15382_ (.A(net183),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][57] ),
    .S(_02340_),
    .Z(_01918_));
 MUX2_X1 _15383_ (.A(net184),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][58] ),
    .S(_02340_),
    .Z(_01919_));
 MUX2_X1 _15384_ (.A(net185),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][59] ),
    .S(_02340_),
    .Z(_01920_));
 MUX2_X1 _15385_ (.A(net186),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][5] ),
    .S(_02340_),
    .Z(_01921_));
 MUX2_X1 _15386_ (.A(net187),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][60] ),
    .S(_02340_),
    .Z(_01922_));
 MUX2_X1 _15387_ (.A(net188),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][61] ),
    .S(_02340_),
    .Z(_01923_));
 MUX2_X1 _15388_ (.A(net189),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][62] ),
    .S(_02340_),
    .Z(_01924_));
 MUX2_X1 _15389_ (.A(net190),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][63] ),
    .S(_02340_),
    .Z(_01925_));
 MUX2_X1 _15390_ (.A(net191),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][6] ),
    .S(_02334_),
    .Z(_01926_));
 MUX2_X1 _15391_ (.A(net192),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][7] ),
    .S(_02334_),
    .Z(_01927_));
 MUX2_X1 _15392_ (.A(net193),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][8] ),
    .S(_02334_),
    .Z(_01928_));
 MUX2_X1 _15393_ (.A(net194),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][9] ),
    .S(_02334_),
    .Z(_01929_));
 NAND2_X1 _15394_ (.A1(_10607_),
    .A2(_02316_),
    .ZN(_02341_));
 BUF_X4 _15395_ (.A(_02341_),
    .Z(_02342_));
 CLKBUF_X3 _15396_ (.A(_02342_),
    .Z(_02343_));
 MUX2_X1 _15397_ (.A(net131),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][0] ),
    .S(_02343_),
    .Z(_01930_));
 MUX2_X1 _15398_ (.A(net132),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][10] ),
    .S(_02343_),
    .Z(_01931_));
 MUX2_X1 _15399_ (.A(net133),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][11] ),
    .S(_02343_),
    .Z(_01932_));
 MUX2_X1 _15400_ (.A(net134),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][12] ),
    .S(_02343_),
    .Z(_01933_));
 MUX2_X1 _15401_ (.A(net135),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][13] ),
    .S(_02343_),
    .Z(_01934_));
 MUX2_X1 _15402_ (.A(net136),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][14] ),
    .S(_02343_),
    .Z(_01935_));
 MUX2_X1 _15403_ (.A(net137),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][15] ),
    .S(_02343_),
    .Z(_01936_));
 MUX2_X1 _15404_ (.A(net138),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][16] ),
    .S(_02343_),
    .Z(_01937_));
 MUX2_X1 _15405_ (.A(net139),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][17] ),
    .S(_02343_),
    .Z(_01938_));
 MUX2_X1 _15406_ (.A(net140),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][18] ),
    .S(_02343_),
    .Z(_01939_));
 CLKBUF_X3 _15407_ (.A(_02342_),
    .Z(_02344_));
 MUX2_X1 _15408_ (.A(net141),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][19] ),
    .S(_02344_),
    .Z(_01940_));
 MUX2_X1 _15409_ (.A(net142),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][1] ),
    .S(_02344_),
    .Z(_01941_));
 MUX2_X1 _15410_ (.A(net143),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][20] ),
    .S(_02344_),
    .Z(_01942_));
 MUX2_X1 _15411_ (.A(net144),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][21] ),
    .S(_02344_),
    .Z(_01943_));
 MUX2_X1 _15412_ (.A(net145),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][22] ),
    .S(_02344_),
    .Z(_01944_));
 MUX2_X1 _15413_ (.A(net146),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][23] ),
    .S(_02344_),
    .Z(_01945_));
 MUX2_X1 _15414_ (.A(net147),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][24] ),
    .S(_02344_),
    .Z(_01946_));
 MUX2_X1 _15415_ (.A(net148),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][25] ),
    .S(_02344_),
    .Z(_01947_));
 MUX2_X1 _15416_ (.A(net149),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][26] ),
    .S(_02344_),
    .Z(_01948_));
 MUX2_X1 _15417_ (.A(net150),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][27] ),
    .S(_02344_),
    .Z(_01949_));
 BUF_X4 _15418_ (.A(_02342_),
    .Z(_02345_));
 MUX2_X1 _15419_ (.A(net151),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][28] ),
    .S(_02345_),
    .Z(_01950_));
 MUX2_X1 _15420_ (.A(net152),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][29] ),
    .S(_02345_),
    .Z(_01951_));
 MUX2_X1 _15421_ (.A(net153),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][2] ),
    .S(_02345_),
    .Z(_01952_));
 MUX2_X1 _15422_ (.A(net154),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][30] ),
    .S(_02345_),
    .Z(_01953_));
 MUX2_X1 _15423_ (.A(net155),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][31] ),
    .S(_02345_),
    .Z(_01954_));
 MUX2_X1 _15424_ (.A(net156),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][32] ),
    .S(_02345_),
    .Z(_01955_));
 MUX2_X1 _15425_ (.A(net157),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][33] ),
    .S(_02345_),
    .Z(_01956_));
 MUX2_X1 _15426_ (.A(net158),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][34] ),
    .S(_02345_),
    .Z(_01957_));
 MUX2_X1 _15427_ (.A(net159),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][35] ),
    .S(_02345_),
    .Z(_01958_));
 MUX2_X1 _15428_ (.A(net160),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][36] ),
    .S(_02345_),
    .Z(_01959_));
 BUF_X4 _15429_ (.A(_02342_),
    .Z(_02346_));
 MUX2_X1 _15430_ (.A(net161),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][37] ),
    .S(_02346_),
    .Z(_01960_));
 MUX2_X1 _15431_ (.A(net162),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][38] ),
    .S(_02346_),
    .Z(_01961_));
 MUX2_X1 _15432_ (.A(net163),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][39] ),
    .S(_02346_),
    .Z(_01962_));
 MUX2_X1 _15433_ (.A(net164),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][3] ),
    .S(_02346_),
    .Z(_01963_));
 MUX2_X1 _15434_ (.A(net165),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][40] ),
    .S(_02346_),
    .Z(_01964_));
 MUX2_X1 _15435_ (.A(net166),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][41] ),
    .S(_02346_),
    .Z(_01965_));
 MUX2_X1 _15436_ (.A(net167),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][42] ),
    .S(_02346_),
    .Z(_01966_));
 MUX2_X1 _15437_ (.A(net168),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][43] ),
    .S(_02346_),
    .Z(_01967_));
 MUX2_X1 _15438_ (.A(net169),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][44] ),
    .S(_02346_),
    .Z(_01968_));
 MUX2_X1 _15439_ (.A(net170),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][45] ),
    .S(_02346_),
    .Z(_01969_));
 BUF_X4 _15440_ (.A(_02342_),
    .Z(_02347_));
 MUX2_X1 _15441_ (.A(net171),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][46] ),
    .S(_02347_),
    .Z(_01970_));
 MUX2_X1 _15442_ (.A(net172),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][47] ),
    .S(_02347_),
    .Z(_01971_));
 MUX2_X1 _15443_ (.A(net173),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][48] ),
    .S(_02347_),
    .Z(_01972_));
 MUX2_X1 _15444_ (.A(net174),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][49] ),
    .S(_02347_),
    .Z(_01973_));
 MUX2_X1 _15445_ (.A(net175),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][4] ),
    .S(_02347_),
    .Z(_01974_));
 MUX2_X1 _15446_ (.A(net176),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][50] ),
    .S(_02347_),
    .Z(_01975_));
 MUX2_X1 _15447_ (.A(net177),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][51] ),
    .S(_02347_),
    .Z(_01976_));
 MUX2_X1 _15448_ (.A(net178),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][52] ),
    .S(_02347_),
    .Z(_01977_));
 MUX2_X1 _15449_ (.A(net179),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][53] ),
    .S(_02347_),
    .Z(_01978_));
 MUX2_X1 _15450_ (.A(net180),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][54] ),
    .S(_02347_),
    .Z(_01979_));
 BUF_X4 _15451_ (.A(_02342_),
    .Z(_02348_));
 MUX2_X1 _15452_ (.A(net181),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][55] ),
    .S(_02348_),
    .Z(_01980_));
 MUX2_X1 _15453_ (.A(net182),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][56] ),
    .S(_02348_),
    .Z(_01981_));
 MUX2_X1 _15454_ (.A(net183),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][57] ),
    .S(_02348_),
    .Z(_01982_));
 MUX2_X1 _15455_ (.A(net184),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][58] ),
    .S(_02348_),
    .Z(_01983_));
 MUX2_X1 _15456_ (.A(net185),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][59] ),
    .S(_02348_),
    .Z(_01984_));
 MUX2_X1 _15457_ (.A(net186),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][5] ),
    .S(_02348_),
    .Z(_01985_));
 MUX2_X1 _15458_ (.A(net187),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][60] ),
    .S(_02348_),
    .Z(_01986_));
 MUX2_X1 _15459_ (.A(net188),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][61] ),
    .S(_02348_),
    .Z(_01987_));
 MUX2_X1 _15460_ (.A(net189),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][62] ),
    .S(_02348_),
    .Z(_01988_));
 MUX2_X1 _15461_ (.A(net190),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][63] ),
    .S(_02348_),
    .Z(_01989_));
 MUX2_X1 _15462_ (.A(net191),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][6] ),
    .S(_02342_),
    .Z(_01990_));
 MUX2_X1 _15463_ (.A(net192),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][7] ),
    .S(_02342_),
    .Z(_01991_));
 MUX2_X1 _15464_ (.A(net193),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][8] ),
    .S(_02342_),
    .Z(_01992_));
 MUX2_X1 _15465_ (.A(net194),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][9] ),
    .S(_02342_),
    .Z(_01993_));
 NOR2_X2 _15466_ (.A1(_06540_),
    .A2(_10497_),
    .ZN(_02349_));
 NAND2_X1 _15467_ (.A1(_10610_),
    .A2(_02349_),
    .ZN(_02350_));
 BUF_X4 _15468_ (.A(_02350_),
    .Z(_02351_));
 BUF_X4 _15469_ (.A(_02351_),
    .Z(_02352_));
 MUX2_X1 _15470_ (.A(net195),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][0] ),
    .S(_02352_),
    .Z(_02019_));
 MUX2_X1 _15471_ (.A(net196),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][10] ),
    .S(_02352_),
    .Z(_02020_));
 MUX2_X1 _15472_ (.A(net197),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][11] ),
    .S(_02352_),
    .Z(_02021_));
 MUX2_X1 _15473_ (.A(net198),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][12] ),
    .S(_02352_),
    .Z(_02022_));
 MUX2_X1 _15474_ (.A(net199),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][13] ),
    .S(_02352_),
    .Z(_02023_));
 MUX2_X1 _15475_ (.A(net200),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][14] ),
    .S(_02352_),
    .Z(_02024_));
 MUX2_X1 _15476_ (.A(net201),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][15] ),
    .S(_02352_),
    .Z(_02025_));
 MUX2_X1 _15477_ (.A(net202),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][16] ),
    .S(_02352_),
    .Z(_02026_));
 MUX2_X1 _15478_ (.A(net203),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][17] ),
    .S(_02352_),
    .Z(_02027_));
 MUX2_X1 _15479_ (.A(net204),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][18] ),
    .S(_02352_),
    .Z(_02028_));
 BUF_X4 _15480_ (.A(_02351_),
    .Z(_02353_));
 MUX2_X1 _15481_ (.A(net205),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][19] ),
    .S(_02353_),
    .Z(_02029_));
 MUX2_X1 _15482_ (.A(net206),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][1] ),
    .S(_02353_),
    .Z(_02030_));
 MUX2_X1 _15483_ (.A(net207),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][20] ),
    .S(_02353_),
    .Z(_02031_));
 MUX2_X1 _15484_ (.A(net208),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][21] ),
    .S(_02353_),
    .Z(_02032_));
 MUX2_X1 _15485_ (.A(net209),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][22] ),
    .S(_02353_),
    .Z(_02033_));
 MUX2_X1 _15486_ (.A(net210),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][23] ),
    .S(_02353_),
    .Z(_02034_));
 MUX2_X1 _15487_ (.A(net211),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][24] ),
    .S(_02353_),
    .Z(_02035_));
 MUX2_X1 _15488_ (.A(net212),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][25] ),
    .S(_02353_),
    .Z(_02036_));
 MUX2_X1 _15489_ (.A(net213),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][26] ),
    .S(_02353_),
    .Z(_02037_));
 MUX2_X1 _15490_ (.A(net214),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][27] ),
    .S(_02353_),
    .Z(_02038_));
 BUF_X4 _15491_ (.A(_02351_),
    .Z(_02354_));
 MUX2_X1 _15492_ (.A(net215),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][28] ),
    .S(_02354_),
    .Z(_02039_));
 MUX2_X1 _15493_ (.A(net216),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][29] ),
    .S(_02354_),
    .Z(_02040_));
 MUX2_X1 _15494_ (.A(net217),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][2] ),
    .S(_02354_),
    .Z(_02041_));
 MUX2_X1 _15495_ (.A(net218),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][30] ),
    .S(_02354_),
    .Z(_02042_));
 MUX2_X1 _15496_ (.A(net219),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][31] ),
    .S(_02354_),
    .Z(_02043_));
 MUX2_X1 _15497_ (.A(net220),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][32] ),
    .S(_02354_),
    .Z(_02044_));
 MUX2_X1 _15498_ (.A(net221),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][33] ),
    .S(_02354_),
    .Z(_02045_));
 MUX2_X1 _15499_ (.A(net222),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][34] ),
    .S(_02354_),
    .Z(_02046_));
 MUX2_X1 _15500_ (.A(net223),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][35] ),
    .S(_02354_),
    .Z(_02047_));
 MUX2_X1 _15501_ (.A(net224),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][36] ),
    .S(_02354_),
    .Z(_02048_));
 BUF_X4 _15502_ (.A(_02351_),
    .Z(_02355_));
 MUX2_X1 _15503_ (.A(net225),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][37] ),
    .S(_02355_),
    .Z(_02049_));
 MUX2_X1 _15504_ (.A(net226),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][38] ),
    .S(_02355_),
    .Z(_02050_));
 MUX2_X1 _15505_ (.A(net227),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][39] ),
    .S(_02355_),
    .Z(_02051_));
 MUX2_X1 _15506_ (.A(net228),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][3] ),
    .S(_02355_),
    .Z(_02052_));
 MUX2_X1 _15507_ (.A(net229),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][40] ),
    .S(_02355_),
    .Z(_02053_));
 MUX2_X1 _15508_ (.A(net230),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][41] ),
    .S(_02355_),
    .Z(_02054_));
 MUX2_X1 _15509_ (.A(net231),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][42] ),
    .S(_02355_),
    .Z(_02055_));
 MUX2_X1 _15510_ (.A(net232),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][43] ),
    .S(_02355_),
    .Z(_02056_));
 MUX2_X1 _15511_ (.A(net233),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][44] ),
    .S(_02355_),
    .Z(_02057_));
 MUX2_X1 _15512_ (.A(net234),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][45] ),
    .S(_02355_),
    .Z(_02058_));
 BUF_X4 _15513_ (.A(_02351_),
    .Z(_02356_));
 MUX2_X1 _15514_ (.A(net235),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][46] ),
    .S(_02356_),
    .Z(_02059_));
 MUX2_X1 _15515_ (.A(net236),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][47] ),
    .S(_02356_),
    .Z(_02060_));
 MUX2_X1 _15516_ (.A(net237),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][48] ),
    .S(_02356_),
    .Z(_02061_));
 MUX2_X1 _15517_ (.A(net238),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][49] ),
    .S(_02356_),
    .Z(_02062_));
 MUX2_X1 _15518_ (.A(net239),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][4] ),
    .S(_02356_),
    .Z(_02063_));
 MUX2_X1 _15519_ (.A(net240),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][50] ),
    .S(_02356_),
    .Z(_02064_));
 MUX2_X1 _15520_ (.A(net241),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][51] ),
    .S(_02356_),
    .Z(_02065_));
 MUX2_X1 _15521_ (.A(net242),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][52] ),
    .S(_02356_),
    .Z(_02066_));
 MUX2_X1 _15522_ (.A(net243),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][53] ),
    .S(_02356_),
    .Z(_02067_));
 MUX2_X1 _15523_ (.A(net244),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][54] ),
    .S(_02356_),
    .Z(_02068_));
 BUF_X4 _15524_ (.A(_02351_),
    .Z(_02357_));
 MUX2_X1 _15525_ (.A(net245),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][55] ),
    .S(_02357_),
    .Z(_02069_));
 MUX2_X1 _15526_ (.A(net246),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][56] ),
    .S(_02357_),
    .Z(_02070_));
 MUX2_X1 _15527_ (.A(net247),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][57] ),
    .S(_02357_),
    .Z(_02071_));
 MUX2_X1 _15528_ (.A(net248),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][58] ),
    .S(_02357_),
    .Z(_02072_));
 MUX2_X1 _15529_ (.A(net249),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][59] ),
    .S(_02357_),
    .Z(_02073_));
 MUX2_X1 _15530_ (.A(net250),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][5] ),
    .S(_02357_),
    .Z(_02074_));
 MUX2_X1 _15531_ (.A(net251),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][60] ),
    .S(_02357_),
    .Z(_02075_));
 MUX2_X1 _15532_ (.A(net252),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][61] ),
    .S(_02357_),
    .Z(_02076_));
 MUX2_X1 _15533_ (.A(net253),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][62] ),
    .S(_02357_),
    .Z(_02077_));
 MUX2_X1 _15534_ (.A(net254),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][63] ),
    .S(_02357_),
    .Z(_02078_));
 MUX2_X1 _15535_ (.A(net255),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][6] ),
    .S(_02351_),
    .Z(_02079_));
 MUX2_X1 _15536_ (.A(net256),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][7] ),
    .S(_02351_),
    .Z(_02080_));
 MUX2_X1 _15537_ (.A(net257),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][8] ),
    .S(_02351_),
    .Z(_02081_));
 MUX2_X1 _15538_ (.A(net258),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[0][9] ),
    .S(_02351_),
    .Z(_02082_));
 NAND2_X1 _15539_ (.A1(_10613_),
    .A2(_02349_),
    .ZN(_02358_));
 BUF_X4 _15540_ (.A(_02358_),
    .Z(_02359_));
 BUF_X4 _15541_ (.A(_02359_),
    .Z(_02360_));
 MUX2_X1 _15542_ (.A(net195),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][0] ),
    .S(_02360_),
    .Z(_02083_));
 MUX2_X1 _15543_ (.A(net196),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][10] ),
    .S(_02360_),
    .Z(_02084_));
 MUX2_X1 _15544_ (.A(net197),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][11] ),
    .S(_02360_),
    .Z(_02085_));
 MUX2_X1 _15545_ (.A(net198),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][12] ),
    .S(_02360_),
    .Z(_02086_));
 MUX2_X1 _15546_ (.A(net199),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][13] ),
    .S(_02360_),
    .Z(_02087_));
 MUX2_X1 _15547_ (.A(net200),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][14] ),
    .S(_02360_),
    .Z(_02088_));
 MUX2_X1 _15548_ (.A(net201),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][15] ),
    .S(_02360_),
    .Z(_02089_));
 MUX2_X1 _15549_ (.A(net202),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][16] ),
    .S(_02360_),
    .Z(_02090_));
 MUX2_X1 _15550_ (.A(net203),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][17] ),
    .S(_02360_),
    .Z(_02091_));
 MUX2_X1 _15551_ (.A(net204),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][18] ),
    .S(_02360_),
    .Z(_02092_));
 BUF_X4 _15552_ (.A(_02359_),
    .Z(_02361_));
 MUX2_X1 _15553_ (.A(net205),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][19] ),
    .S(_02361_),
    .Z(_02093_));
 MUX2_X1 _15554_ (.A(net206),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][1] ),
    .S(_02361_),
    .Z(_02094_));
 MUX2_X1 _15555_ (.A(net207),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][20] ),
    .S(_02361_),
    .Z(_02095_));
 MUX2_X1 _15556_ (.A(net208),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][21] ),
    .S(_02361_),
    .Z(_02096_));
 MUX2_X1 _15557_ (.A(net209),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][22] ),
    .S(_02361_),
    .Z(_02097_));
 MUX2_X1 _15558_ (.A(net210),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][23] ),
    .S(_02361_),
    .Z(_02098_));
 MUX2_X1 _15559_ (.A(net211),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][24] ),
    .S(_02361_),
    .Z(_02099_));
 MUX2_X1 _15560_ (.A(net212),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][25] ),
    .S(_02361_),
    .Z(_02100_));
 MUX2_X1 _15561_ (.A(net213),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][26] ),
    .S(_02361_),
    .Z(_02101_));
 MUX2_X1 _15562_ (.A(net214),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][27] ),
    .S(_02361_),
    .Z(_02102_));
 BUF_X4 _15563_ (.A(_02359_),
    .Z(_02362_));
 MUX2_X1 _15564_ (.A(net215),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][28] ),
    .S(_02362_),
    .Z(_02103_));
 MUX2_X1 _15565_ (.A(net216),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][29] ),
    .S(_02362_),
    .Z(_02104_));
 MUX2_X1 _15566_ (.A(net217),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][2] ),
    .S(_02362_),
    .Z(_02105_));
 MUX2_X1 _15567_ (.A(net218),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][30] ),
    .S(_02362_),
    .Z(_02106_));
 MUX2_X1 _15568_ (.A(net219),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][31] ),
    .S(_02362_),
    .Z(_02107_));
 MUX2_X1 _15569_ (.A(net220),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][32] ),
    .S(_02362_),
    .Z(_02108_));
 MUX2_X1 _15570_ (.A(net221),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][33] ),
    .S(_02362_),
    .Z(_02109_));
 MUX2_X1 _15571_ (.A(net222),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][34] ),
    .S(_02362_),
    .Z(_02110_));
 MUX2_X1 _15572_ (.A(net223),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][35] ),
    .S(_02362_),
    .Z(_02111_));
 MUX2_X1 _15573_ (.A(net224),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][36] ),
    .S(_02362_),
    .Z(_02112_));
 BUF_X4 _15574_ (.A(_02359_),
    .Z(_02363_));
 MUX2_X1 _15575_ (.A(net225),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][37] ),
    .S(_02363_),
    .Z(_02113_));
 MUX2_X1 _15576_ (.A(net226),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][38] ),
    .S(_02363_),
    .Z(_02114_));
 MUX2_X1 _15577_ (.A(net227),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][39] ),
    .S(_02363_),
    .Z(_02115_));
 MUX2_X1 _15578_ (.A(net228),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][3] ),
    .S(_02363_),
    .Z(_02116_));
 MUX2_X1 _15579_ (.A(net229),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][40] ),
    .S(_02363_),
    .Z(_02117_));
 MUX2_X1 _15580_ (.A(net230),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][41] ),
    .S(_02363_),
    .Z(_02118_));
 MUX2_X1 _15581_ (.A(net231),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][42] ),
    .S(_02363_),
    .Z(_02119_));
 MUX2_X1 _15582_ (.A(net232),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][43] ),
    .S(_02363_),
    .Z(_02120_));
 MUX2_X1 _15583_ (.A(net233),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][44] ),
    .S(_02363_),
    .Z(_02121_));
 MUX2_X1 _15584_ (.A(net234),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][45] ),
    .S(_02363_),
    .Z(_02122_));
 BUF_X4 _15585_ (.A(_02359_),
    .Z(_02364_));
 MUX2_X1 _15586_ (.A(net235),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][46] ),
    .S(_02364_),
    .Z(_02123_));
 MUX2_X1 _15587_ (.A(net236),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][47] ),
    .S(_02364_),
    .Z(_02124_));
 MUX2_X1 _15588_ (.A(net237),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][48] ),
    .S(_02364_),
    .Z(_02125_));
 MUX2_X1 _15589_ (.A(net238),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][49] ),
    .S(_02364_),
    .Z(_02126_));
 MUX2_X1 _15590_ (.A(net239),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][4] ),
    .S(_02364_),
    .Z(_02127_));
 MUX2_X1 _15591_ (.A(net240),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][50] ),
    .S(_02364_),
    .Z(_02128_));
 MUX2_X1 _15592_ (.A(net241),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][51] ),
    .S(_02364_),
    .Z(_02129_));
 MUX2_X1 _15593_ (.A(net242),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][52] ),
    .S(_02364_),
    .Z(_02130_));
 MUX2_X1 _15594_ (.A(net243),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][53] ),
    .S(_02364_),
    .Z(_02131_));
 MUX2_X1 _15595_ (.A(net244),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][54] ),
    .S(_02364_),
    .Z(_02132_));
 BUF_X4 _15596_ (.A(_02359_),
    .Z(_02365_));
 MUX2_X1 _15597_ (.A(net245),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][55] ),
    .S(_02365_),
    .Z(_02133_));
 MUX2_X1 _15598_ (.A(net246),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][56] ),
    .S(_02365_),
    .Z(_02134_));
 MUX2_X1 _15599_ (.A(net247),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][57] ),
    .S(_02365_),
    .Z(_02135_));
 MUX2_X1 _15600_ (.A(net248),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][58] ),
    .S(_02365_),
    .Z(_02136_));
 MUX2_X1 _15601_ (.A(net249),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][59] ),
    .S(_02365_),
    .Z(_02137_));
 MUX2_X1 _15602_ (.A(net250),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][5] ),
    .S(_02365_),
    .Z(_02138_));
 MUX2_X1 _15603_ (.A(net251),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][60] ),
    .S(_02365_),
    .Z(_02139_));
 MUX2_X1 _15604_ (.A(net252),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][61] ),
    .S(_02365_),
    .Z(_02140_));
 MUX2_X1 _15605_ (.A(net253),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][62] ),
    .S(_02365_),
    .Z(_02141_));
 MUX2_X1 _15606_ (.A(net254),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][63] ),
    .S(_02365_),
    .Z(_02142_));
 MUX2_X1 _15607_ (.A(net255),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][6] ),
    .S(_02359_),
    .Z(_02143_));
 MUX2_X1 _15608_ (.A(net256),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][7] ),
    .S(_02359_),
    .Z(_02144_));
 MUX2_X1 _15609_ (.A(net257),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][8] ),
    .S(_02359_),
    .Z(_02145_));
 MUX2_X1 _15610_ (.A(net258),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[1][9] ),
    .S(_02359_),
    .Z(_02146_));
 NAND2_X1 _15611_ (.A1(_10611_),
    .A2(_02349_),
    .ZN(_02366_));
 BUF_X4 _15612_ (.A(_02366_),
    .Z(_02367_));
 BUF_X4 _15613_ (.A(_02367_),
    .Z(_02368_));
 MUX2_X1 _15614_ (.A(net195),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][0] ),
    .S(_02368_),
    .Z(_02147_));
 MUX2_X1 _15615_ (.A(net196),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][10] ),
    .S(_02368_),
    .Z(_02148_));
 MUX2_X1 _15616_ (.A(net197),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][11] ),
    .S(_02368_),
    .Z(_02149_));
 MUX2_X1 _15617_ (.A(net198),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][12] ),
    .S(_02368_),
    .Z(_02150_));
 MUX2_X1 _15618_ (.A(net199),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][13] ),
    .S(_02368_),
    .Z(_02151_));
 MUX2_X1 _15619_ (.A(net200),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][14] ),
    .S(_02368_),
    .Z(_02152_));
 MUX2_X1 _15620_ (.A(net201),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][15] ),
    .S(_02368_),
    .Z(_02153_));
 MUX2_X1 _15621_ (.A(net202),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][16] ),
    .S(_02368_),
    .Z(_02154_));
 MUX2_X1 _15622_ (.A(net203),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][17] ),
    .S(_02368_),
    .Z(_02155_));
 MUX2_X1 _15623_ (.A(net204),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][18] ),
    .S(_02368_),
    .Z(_02156_));
 BUF_X4 _15624_ (.A(_02367_),
    .Z(_02369_));
 MUX2_X1 _15625_ (.A(net205),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][19] ),
    .S(_02369_),
    .Z(_02157_));
 MUX2_X1 _15626_ (.A(net206),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][1] ),
    .S(_02369_),
    .Z(_02158_));
 MUX2_X1 _15627_ (.A(net207),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][20] ),
    .S(_02369_),
    .Z(_02159_));
 MUX2_X1 _15628_ (.A(net208),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][21] ),
    .S(_02369_),
    .Z(_02160_));
 MUX2_X1 _15629_ (.A(net209),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][22] ),
    .S(_02369_),
    .Z(_02161_));
 MUX2_X1 _15630_ (.A(net210),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][23] ),
    .S(_02369_),
    .Z(_02162_));
 MUX2_X1 _15631_ (.A(net211),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][24] ),
    .S(_02369_),
    .Z(_02163_));
 MUX2_X1 _15632_ (.A(net212),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][25] ),
    .S(_02369_),
    .Z(_02164_));
 MUX2_X1 _15633_ (.A(net213),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][26] ),
    .S(_02369_),
    .Z(_02165_));
 MUX2_X1 _15634_ (.A(net214),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][27] ),
    .S(_02369_),
    .Z(_02166_));
 BUF_X4 _15635_ (.A(_02367_),
    .Z(_02370_));
 MUX2_X1 _15636_ (.A(net215),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][28] ),
    .S(_02370_),
    .Z(_02167_));
 MUX2_X1 _15637_ (.A(net216),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][29] ),
    .S(_02370_),
    .Z(_02168_));
 MUX2_X1 _15638_ (.A(net217),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][2] ),
    .S(_02370_),
    .Z(_02169_));
 MUX2_X1 _15639_ (.A(net218),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][30] ),
    .S(_02370_),
    .Z(_02170_));
 MUX2_X1 _15640_ (.A(net219),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][31] ),
    .S(_02370_),
    .Z(_02171_));
 MUX2_X1 _15641_ (.A(net220),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][32] ),
    .S(_02370_),
    .Z(_02172_));
 MUX2_X1 _15642_ (.A(net221),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][33] ),
    .S(_02370_),
    .Z(_02173_));
 MUX2_X1 _15643_ (.A(net222),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][34] ),
    .S(_02370_),
    .Z(_02174_));
 MUX2_X1 _15644_ (.A(net223),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][35] ),
    .S(_02370_),
    .Z(_02175_));
 MUX2_X1 _15645_ (.A(net224),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][36] ),
    .S(_02370_),
    .Z(_02176_));
 BUF_X4 _15646_ (.A(_02367_),
    .Z(_02371_));
 MUX2_X1 _15647_ (.A(net225),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][37] ),
    .S(_02371_),
    .Z(_02177_));
 MUX2_X1 _15648_ (.A(net226),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][38] ),
    .S(_02371_),
    .Z(_02178_));
 MUX2_X1 _15649_ (.A(net227),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][39] ),
    .S(_02371_),
    .Z(_02179_));
 MUX2_X1 _15650_ (.A(net228),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][3] ),
    .S(_02371_),
    .Z(_02180_));
 MUX2_X1 _15651_ (.A(net229),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][40] ),
    .S(_02371_),
    .Z(_02181_));
 MUX2_X1 _15652_ (.A(net230),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][41] ),
    .S(_02371_),
    .Z(_02182_));
 MUX2_X1 _15653_ (.A(net231),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][42] ),
    .S(_02371_),
    .Z(_02183_));
 MUX2_X1 _15654_ (.A(net232),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][43] ),
    .S(_02371_),
    .Z(_02184_));
 MUX2_X1 _15655_ (.A(net233),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][44] ),
    .S(_02371_),
    .Z(_02185_));
 MUX2_X1 _15656_ (.A(net234),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][45] ),
    .S(_02371_),
    .Z(_02186_));
 BUF_X4 _15657_ (.A(_02367_),
    .Z(_02372_));
 MUX2_X1 _15658_ (.A(net235),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][46] ),
    .S(_02372_),
    .Z(_02187_));
 MUX2_X1 _15659_ (.A(net236),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][47] ),
    .S(_02372_),
    .Z(_02188_));
 MUX2_X1 _15660_ (.A(net237),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][48] ),
    .S(_02372_),
    .Z(_02189_));
 MUX2_X1 _15661_ (.A(net238),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][49] ),
    .S(_02372_),
    .Z(_02190_));
 MUX2_X1 _15662_ (.A(net239),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][4] ),
    .S(_02372_),
    .Z(_02191_));
 MUX2_X1 _15663_ (.A(net240),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][50] ),
    .S(_02372_),
    .Z(_02192_));
 MUX2_X1 _15664_ (.A(net241),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][51] ),
    .S(_02372_),
    .Z(_02193_));
 MUX2_X1 _15665_ (.A(net242),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][52] ),
    .S(_02372_),
    .Z(_02194_));
 MUX2_X1 _15666_ (.A(net243),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][53] ),
    .S(_02372_),
    .Z(_02195_));
 MUX2_X1 _15667_ (.A(net244),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][54] ),
    .S(_02372_),
    .Z(_02196_));
 BUF_X4 _15668_ (.A(_02367_),
    .Z(_02373_));
 MUX2_X1 _15669_ (.A(net245),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][55] ),
    .S(_02373_),
    .Z(_02197_));
 MUX2_X1 _15670_ (.A(net246),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][56] ),
    .S(_02373_),
    .Z(_02198_));
 MUX2_X1 _15671_ (.A(net247),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][57] ),
    .S(_02373_),
    .Z(_02199_));
 MUX2_X1 _15672_ (.A(net248),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][58] ),
    .S(_02373_),
    .Z(_02200_));
 MUX2_X1 _15673_ (.A(net249),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][59] ),
    .S(_02373_),
    .Z(_02201_));
 MUX2_X1 _15674_ (.A(net250),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][5] ),
    .S(_02373_),
    .Z(_02202_));
 MUX2_X1 _15675_ (.A(net251),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][60] ),
    .S(_02373_),
    .Z(_02203_));
 MUX2_X1 _15676_ (.A(net252),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][61] ),
    .S(_02373_),
    .Z(_02204_));
 MUX2_X1 _15677_ (.A(net253),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][62] ),
    .S(_02373_),
    .Z(_02205_));
 MUX2_X1 _15678_ (.A(net254),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][63] ),
    .S(_02373_),
    .Z(_02206_));
 MUX2_X1 _15679_ (.A(net255),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][6] ),
    .S(_02367_),
    .Z(_02207_));
 MUX2_X1 _15680_ (.A(net256),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][7] ),
    .S(_02367_),
    .Z(_02208_));
 MUX2_X1 _15681_ (.A(net257),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][8] ),
    .S(_02367_),
    .Z(_02209_));
 MUX2_X1 _15682_ (.A(net258),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][9] ),
    .S(_02367_),
    .Z(_02210_));
 NAND2_X1 _15683_ (.A1(_10615_),
    .A2(_02349_),
    .ZN(_02374_));
 BUF_X4 _15684_ (.A(_02374_),
    .Z(_02375_));
 BUF_X4 _15685_ (.A(_02375_),
    .Z(_02376_));
 MUX2_X1 _15686_ (.A(net195),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][0] ),
    .S(_02376_),
    .Z(_02211_));
 MUX2_X1 _15687_ (.A(net196),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][10] ),
    .S(_02376_),
    .Z(_02212_));
 MUX2_X1 _15688_ (.A(net197),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][11] ),
    .S(_02376_),
    .Z(_02213_));
 MUX2_X1 _15689_ (.A(net198),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][12] ),
    .S(_02376_),
    .Z(_02214_));
 MUX2_X1 _15690_ (.A(net199),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][13] ),
    .S(_02376_),
    .Z(_02215_));
 MUX2_X1 _15691_ (.A(net200),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][14] ),
    .S(_02376_),
    .Z(_02216_));
 MUX2_X1 _15692_ (.A(net201),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][15] ),
    .S(_02376_),
    .Z(_02217_));
 MUX2_X1 _15693_ (.A(net202),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][16] ),
    .S(_02376_),
    .Z(_02218_));
 MUX2_X1 _15694_ (.A(net203),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][17] ),
    .S(_02376_),
    .Z(_02219_));
 MUX2_X1 _15695_ (.A(net204),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][18] ),
    .S(_02376_),
    .Z(_02220_));
 BUF_X4 _15696_ (.A(_02375_),
    .Z(_02377_));
 MUX2_X1 _15697_ (.A(net205),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][19] ),
    .S(_02377_),
    .Z(_02221_));
 MUX2_X1 _15698_ (.A(net206),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][1] ),
    .S(_02377_),
    .Z(_02222_));
 MUX2_X1 _15699_ (.A(net207),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][20] ),
    .S(_02377_),
    .Z(_02223_));
 MUX2_X1 _15700_ (.A(net208),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][21] ),
    .S(_02377_),
    .Z(_02224_));
 MUX2_X1 _15701_ (.A(net209),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][22] ),
    .S(_02377_),
    .Z(_02225_));
 MUX2_X1 _15702_ (.A(net210),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][23] ),
    .S(_02377_),
    .Z(_02226_));
 MUX2_X1 _15703_ (.A(net211),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][24] ),
    .S(_02377_),
    .Z(_02227_));
 MUX2_X1 _15704_ (.A(net212),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][25] ),
    .S(_02377_),
    .Z(_02228_));
 MUX2_X1 _15705_ (.A(net213),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][26] ),
    .S(_02377_),
    .Z(_02229_));
 MUX2_X1 _15706_ (.A(net214),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][27] ),
    .S(_02377_),
    .Z(_02230_));
 BUF_X4 _15707_ (.A(_02375_),
    .Z(_02378_));
 MUX2_X1 _15708_ (.A(net215),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][28] ),
    .S(_02378_),
    .Z(_02231_));
 MUX2_X1 _15709_ (.A(net216),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][29] ),
    .S(_02378_),
    .Z(_02232_));
 MUX2_X1 _15710_ (.A(net217),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][2] ),
    .S(_02378_),
    .Z(_02233_));
 MUX2_X1 _15711_ (.A(net218),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][30] ),
    .S(_02378_),
    .Z(_02234_));
 MUX2_X1 _15712_ (.A(net219),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][31] ),
    .S(_02378_),
    .Z(_02235_));
 MUX2_X1 _15713_ (.A(net220),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][32] ),
    .S(_02378_),
    .Z(_02236_));
 MUX2_X1 _15714_ (.A(net221),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][33] ),
    .S(_02378_),
    .Z(_02237_));
 MUX2_X1 _15715_ (.A(net222),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][34] ),
    .S(_02378_),
    .Z(_02238_));
 MUX2_X1 _15716_ (.A(net223),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][35] ),
    .S(_02378_),
    .Z(_02239_));
 MUX2_X1 _15717_ (.A(net224),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][36] ),
    .S(_02378_),
    .Z(_02240_));
 CLKBUF_X3 _15718_ (.A(_02375_),
    .Z(_02379_));
 MUX2_X1 _15719_ (.A(net225),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][37] ),
    .S(_02379_),
    .Z(_02241_));
 MUX2_X1 _15720_ (.A(net226),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][38] ),
    .S(_02379_),
    .Z(_02242_));
 MUX2_X1 _15721_ (.A(net227),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][39] ),
    .S(_02379_),
    .Z(_02243_));
 MUX2_X1 _15722_ (.A(net228),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][3] ),
    .S(_02379_),
    .Z(_02244_));
 MUX2_X1 _15723_ (.A(net229),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][40] ),
    .S(_02379_),
    .Z(_02245_));
 MUX2_X1 _15724_ (.A(net230),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][41] ),
    .S(_02379_),
    .Z(_02246_));
 MUX2_X1 _15725_ (.A(net231),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][42] ),
    .S(_02379_),
    .Z(_02247_));
 MUX2_X1 _15726_ (.A(net232),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][43] ),
    .S(_02379_),
    .Z(_02248_));
 MUX2_X1 _15727_ (.A(net233),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][44] ),
    .S(_02379_),
    .Z(_02249_));
 MUX2_X1 _15728_ (.A(net234),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][45] ),
    .S(_02379_),
    .Z(_02250_));
 BUF_X4 _15729_ (.A(_02375_),
    .Z(_02380_));
 MUX2_X1 _15730_ (.A(net235),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][46] ),
    .S(_02380_),
    .Z(_02251_));
 MUX2_X1 _15731_ (.A(net236),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][47] ),
    .S(_02380_),
    .Z(_02252_));
 MUX2_X1 _15732_ (.A(net237),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][48] ),
    .S(_02380_),
    .Z(_02253_));
 MUX2_X1 _15733_ (.A(net238),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][49] ),
    .S(_02380_),
    .Z(_02254_));
 MUX2_X1 _15734_ (.A(net239),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][4] ),
    .S(_02380_),
    .Z(_02255_));
 MUX2_X1 _15735_ (.A(net240),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][50] ),
    .S(_02380_),
    .Z(_02256_));
 MUX2_X1 _15736_ (.A(net241),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][51] ),
    .S(_02380_),
    .Z(_02257_));
 MUX2_X1 _15737_ (.A(net242),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][52] ),
    .S(_02380_),
    .Z(_02258_));
 MUX2_X1 _15738_ (.A(net243),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][53] ),
    .S(_02380_),
    .Z(_02259_));
 MUX2_X1 _15739_ (.A(net244),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][54] ),
    .S(_02380_),
    .Z(_02260_));
 BUF_X4 _15740_ (.A(_02375_),
    .Z(_02381_));
 MUX2_X1 _15741_ (.A(net245),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][55] ),
    .S(_02381_),
    .Z(_02261_));
 MUX2_X1 _15742_ (.A(net246),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][56] ),
    .S(_02381_),
    .Z(_02262_));
 MUX2_X1 _15743_ (.A(net247),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][57] ),
    .S(_02381_),
    .Z(_02263_));
 MUX2_X1 _15744_ (.A(net248),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][58] ),
    .S(_02381_),
    .Z(_02264_));
 MUX2_X1 _15745_ (.A(net249),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][59] ),
    .S(_02381_),
    .Z(_02265_));
 MUX2_X1 _15746_ (.A(net250),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][5] ),
    .S(_02381_),
    .Z(_02266_));
 MUX2_X1 _15747_ (.A(net251),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][60] ),
    .S(_02381_),
    .Z(_02267_));
 MUX2_X1 _15748_ (.A(net252),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][61] ),
    .S(_02381_),
    .Z(_02268_));
 MUX2_X1 _15749_ (.A(net253),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][62] ),
    .S(_02381_),
    .Z(_02269_));
 MUX2_X1 _15750_ (.A(net254),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][63] ),
    .S(_02381_),
    .Z(_02270_));
 MUX2_X1 _15751_ (.A(net255),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][6] ),
    .S(_02375_),
    .Z(_02271_));
 MUX2_X1 _15752_ (.A(net256),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][7] ),
    .S(_02375_),
    .Z(_02272_));
 MUX2_X1 _15753_ (.A(net257),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][8] ),
    .S(_02375_),
    .Z(_02273_));
 MUX2_X1 _15754_ (.A(net258),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][9] ),
    .S(_02375_),
    .Z(_02274_));
 BUF_X4 _15755_ (.A(_06589_),
    .Z(_02382_));
 NOR2_X1 _15756_ (.A1(_10499_),
    .A2(_10503_),
    .ZN(_02383_));
 XOR2_X1 _15757_ (.A(\dynamic_node_top.west_input.NIB.head_ptr_next[0] ),
    .B(_02383_),
    .Z(_02384_));
 NOR2_X1 _15758_ (.A1(_02382_),
    .A2(_02384_),
    .ZN(_00077_));
 NAND2_X1 _15759_ (.A1(\dynamic_node_top.west_input.NIB.head_ptr_f[0] ),
    .A2(_02383_),
    .ZN(_02385_));
 XOR2_X2 _15760_ (.A(\dynamic_node_top.west_input.NIB.head_ptr_f[1] ),
    .B(_02385_),
    .Z(_02386_));
 NOR2_X2 _15761_ (.A1(_02382_),
    .A2(_02386_),
    .ZN(_00078_));
 NOR2_X4 _15762_ (.A1(_10469_),
    .A2(_10465_),
    .ZN(_02387_));
 XOR2_X1 _15763_ (.A(\dynamic_node_top.south_input.NIB.head_ptr_next[0] ),
    .B(_02387_),
    .Z(_02388_));
 NOR2_X1 _15764_ (.A1(_02382_),
    .A2(_02388_),
    .ZN(_00079_));
 NAND2_X1 _15765_ (.A1(\dynamic_node_top.south_input.NIB.head_ptr_f[0] ),
    .A2(_02387_),
    .ZN(_02389_));
 XOR2_X1 _15766_ (.A(\dynamic_node_top.south_input.NIB.head_ptr_f[1] ),
    .B(_02389_),
    .Z(_02390_));
 NOR2_X1 _15767_ (.A1(_02382_),
    .A2(_02390_),
    .ZN(_00080_));
 NOR2_X4 _15768_ (.A1(_10507_),
    .A2(_10511_),
    .ZN(_02391_));
 XOR2_X1 _15769_ (.A(\dynamic_node_top.east_input.NIB.head_ptr_next[0] ),
    .B(_02391_),
    .Z(_02392_));
 NOR2_X1 _15770_ (.A1(_02382_),
    .A2(_02392_),
    .ZN(_00081_));
 NAND2_X1 _15771_ (.A1(\dynamic_node_top.east_input.NIB.head_ptr_f[0] ),
    .A2(_02391_),
    .ZN(_02393_));
 XOR2_X1 _15772_ (.A(\dynamic_node_top.east_input.NIB.head_ptr_f[1] ),
    .B(_02393_),
    .Z(_02394_));
 NOR2_X1 _15773_ (.A1(_02382_),
    .A2(_02394_),
    .ZN(_00082_));
 NOR2_X4 _15774_ (.A1(_10458_),
    .A2(_10169_),
    .ZN(_02395_));
 XOR2_X1 _15775_ (.A(\dynamic_node_top.proc_input.NIB.head_ptr_next[0] ),
    .B(_02395_),
    .Z(_02396_));
 NOR2_X1 _15776_ (.A1(_02382_),
    .A2(_02396_),
    .ZN(_00083_));
 MUX2_X1 _15777_ (.A(\dynamic_node_top.proc_input.NIB.head_ptr_f[1] ),
    .B(\dynamic_node_top.proc_input.NIB.head_ptr_next[1] ),
    .S(_02395_),
    .Z(_02397_));
 AND2_X1 _15778_ (.A1(_06892_),
    .A2(_02397_),
    .ZN(_00084_));
 NAND2_X1 _15779_ (.A1(_10592_),
    .A2(_02395_),
    .ZN(_02398_));
 XOR2_X1 _15780_ (.A(\dynamic_node_top.proc_input.NIB.head_ptr_f[2] ),
    .B(_02398_),
    .Z(_02399_));
 NOR2_X1 _15781_ (.A1(_02382_),
    .A2(_02399_),
    .ZN(_00085_));
 NAND4_X1 _15782_ (.A1(\dynamic_node_top.proc_input.NIB.head_ptr_f[2] ),
    .A2(\dynamic_node_top.proc_input.NIB.head_ptr_f[1] ),
    .A3(\dynamic_node_top.proc_input.NIB.head_ptr_f[0] ),
    .A4(_02395_),
    .ZN(_02400_));
 XOR2_X1 _15783_ (.A(\dynamic_node_top.proc_input.NIB.head_ptr_f[3] ),
    .B(_02400_),
    .Z(_02401_));
 NOR2_X1 _15784_ (.A1(_02382_),
    .A2(_02401_),
    .ZN(_00086_));
 NOR2_X2 _15785_ (.A1(_10477_),
    .A2(_10473_),
    .ZN(_02402_));
 XOR2_X1 _15786_ (.A(\dynamic_node_top.north_input.NIB.head_ptr_next[0] ),
    .B(_02402_),
    .Z(_02403_));
 NOR2_X1 _15787_ (.A1(_02382_),
    .A2(_02403_),
    .ZN(_00087_));
 BUF_X4 _15788_ (.A(_06589_),
    .Z(_02404_));
 NAND2_X1 _15789_ (.A1(\dynamic_node_top.north_input.NIB.head_ptr_f[0] ),
    .A2(_02402_),
    .ZN(_02405_));
 XOR2_X2 _15790_ (.A(\dynamic_node_top.north_input.NIB.head_ptr_f[1] ),
    .B(_02405_),
    .Z(_02406_));
 NOR2_X2 _15791_ (.A1(_02404_),
    .A2(_02406_),
    .ZN(_00088_));
 MUX2_X1 _15792_ (.A(\dynamic_node_top.east_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.east_input.NIB.elements_in_array_next[0] ),
    .S(_10508_),
    .Z(_02407_));
 AND2_X1 _15793_ (.A1(_06892_),
    .A2(_02407_),
    .ZN(_00089_));
 NAND2_X1 _15794_ (.A1(_10164_),
    .A2(_10508_),
    .ZN(_02408_));
 OAI21_X1 _15795_ (.A(_02408_),
    .B1(_10508_),
    .B2(\dynamic_node_top.east_input.NIB.elements_in_array_f[1] ),
    .ZN(_02409_));
 NOR2_X1 _15796_ (.A1(_02404_),
    .A2(_02409_),
    .ZN(_00090_));
 XNOR2_X1 _15797_ (.A(_10511_),
    .B(_10163_),
    .ZN(_02410_));
 NAND2_X1 _15798_ (.A1(_10508_),
    .A2(_02410_),
    .ZN(_02411_));
 XOR2_X1 _15799_ (.A(\dynamic_node_top.east_input.NIB.elements_in_array_f[2] ),
    .B(_02411_),
    .Z(_02412_));
 NOR2_X1 _15800_ (.A1(_02404_),
    .A2(_02412_),
    .ZN(_00091_));
 MUX2_X1 _15801_ (.A(\dynamic_node_top.east_input.NIB.head_ptr_f[0] ),
    .B(\dynamic_node_top.east_input.NIB.head_ptr_next[0] ),
    .S(_02391_),
    .Z(_02413_));
 AND2_X1 _15802_ (.A1(_06892_),
    .A2(_02413_),
    .ZN(_00092_));
 NOR2_X4 _15803_ (.A1(_10509_),
    .A2(_10507_),
    .ZN(_02414_));
 MUX2_X1 _15804_ (.A(\dynamic_node_top.east_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.east_input.NIB.tail_ptr_next[0] ),
    .S(_02414_),
    .Z(_02415_));
 AND2_X1 _15805_ (.A1(_06892_),
    .A2(_02415_),
    .ZN(_00349_));
 MUX2_X1 _15806_ (.A(\dynamic_node_top.east_input.NIB.tail_ptr_f[1] ),
    .B(\dynamic_node_top.east_input.NIB.tail_ptr_next[1] ),
    .S(_02414_),
    .Z(_02416_));
 AND2_X1 _15807_ (.A1(_06892_),
    .A2(_02416_),
    .ZN(_00350_));
 AND2_X1 _15808_ (.A1(_06754_),
    .A2(_07211_),
    .ZN(_00351_));
 NOR2_X1 _15809_ (.A1(_05787_),
    .A2(\dynamic_node_top.east_input.control.count_f[1] ),
    .ZN(_02417_));
 AOI221_X2 _15810_ (.A(_02417_),
    .B1(_10441_),
    .B2(_05787_),
    .C1(_05488_),
    .C2(_05177_),
    .ZN(_02418_));
 AOI21_X1 _15811_ (.A(_02418_),
    .B1(_05765_),
    .B2(_06787_),
    .ZN(_02419_));
 NOR2_X1 _15812_ (.A1(_02404_),
    .A2(_02419_),
    .ZN(_00352_));
 BUF_X4 _15813_ (.A(_06589_),
    .Z(_02420_));
 NOR2_X1 _15814_ (.A1(_06793_),
    .A2(_05771_),
    .ZN(_02421_));
 XNOR2_X1 _15815_ (.A(_07212_),
    .B(_07213_),
    .ZN(_02422_));
 NOR2_X1 _15816_ (.A1(_06787_),
    .A2(_02422_),
    .ZN(_02423_));
 NOR3_X1 _15817_ (.A1(_02420_),
    .A2(_02421_),
    .A3(_02423_),
    .ZN(_00353_));
 NOR2_X1 _15818_ (.A1(_06793_),
    .A2(_05768_),
    .ZN(_02424_));
 NOR2_X1 _15819_ (.A1(_06787_),
    .A2(_07219_),
    .ZN(_02425_));
 NOR3_X1 _15820_ (.A1(_02420_),
    .A2(_02424_),
    .A3(_02425_),
    .ZN(_00354_));
 NOR3_X1 _15821_ (.A1(_02420_),
    .A2(_05761_),
    .A3(_07216_),
    .ZN(_00355_));
 NOR2_X1 _15822_ (.A1(_02404_),
    .A2(_07235_),
    .ZN(_00356_));
 NOR2_X1 _15823_ (.A1(_02404_),
    .A2(_07232_),
    .ZN(_00357_));
 AND2_X1 _15824_ (.A1(_06892_),
    .A2(_07228_),
    .ZN(_00358_));
 INV_X1 _15825_ (.A(_00351_),
    .ZN(_02426_));
 NOR4_X1 _15826_ (.A1(_07224_),
    .A2(_07228_),
    .A3(_07236_),
    .A4(_02426_),
    .ZN(_00359_));
 NOR2_X1 _15827_ (.A1(_02404_),
    .A2(_06599_),
    .ZN(_00360_));
 NOR2_X1 _15828_ (.A1(_02404_),
    .A2(_10506_),
    .ZN(_00361_));
 NAND2_X1 _15829_ (.A1(_00046_),
    .A2(_06721_),
    .ZN(_02427_));
 NAND2_X1 _15830_ (.A1(_05307_),
    .A2(_06757_),
    .ZN(_02428_));
 MUX2_X1 _15831_ (.A(_02427_),
    .B(_02428_),
    .S(_06720_),
    .Z(_02429_));
 NAND2_X1 _15832_ (.A1(_00046_),
    .A2(_06756_),
    .ZN(_02430_));
 NAND3_X1 _15833_ (.A1(_06545_),
    .A2(_06789_),
    .A3(_05500_),
    .ZN(_02431_));
 NOR4_X1 _15834_ (.A1(_05304_),
    .A2(_06793_),
    .A3(_06567_),
    .A4(_02431_),
    .ZN(_02432_));
 NOR2_X1 _15835_ (.A1(_06793_),
    .A2(_06839_),
    .ZN(_02433_));
 AOI21_X1 _15836_ (.A(_02432_),
    .B1(_02433_),
    .B2(_06567_),
    .ZN(_02434_));
 AND4_X1 _15837_ (.A1(_05306_),
    .A2(_06752_),
    .A3(_06765_),
    .A4(_02434_),
    .ZN(_02435_));
 NAND3_X1 _15838_ (.A1(_05184_),
    .A2(_06833_),
    .A3(_02435_),
    .ZN(_02436_));
 OAI211_X2 _15839_ (.A(_06755_),
    .B(_02429_),
    .C1(_02430_),
    .C2(_02436_),
    .ZN(_02437_));
 OAI21_X1 _15840_ (.A(_06721_),
    .B1(_06833_),
    .B2(_05158_),
    .ZN(_02438_));
 OAI21_X1 _15841_ (.A(_02438_),
    .B1(_06745_),
    .B2(_05306_),
    .ZN(_02439_));
 NOR2_X1 _15842_ (.A1(_00046_),
    .A2(_05184_),
    .ZN(_02440_));
 AND3_X1 _15843_ (.A1(_06714_),
    .A2(_06719_),
    .A3(_02440_),
    .ZN(_02441_));
 OAI222_X2 _15844_ (.A1(_05173_),
    .A2(_06736_),
    .B1(_06841_),
    .B2(_06724_),
    .C1(_06752_),
    .C2(_05167_),
    .ZN(_02442_));
 NOR2_X1 _15845_ (.A1(_06757_),
    .A2(_06719_),
    .ZN(_02443_));
 OAI21_X1 _15846_ (.A(_06714_),
    .B1(_06765_),
    .B2(_05171_),
    .ZN(_02444_));
 MUX2_X1 _15847_ (.A(_06954_),
    .B(_02444_),
    .S(_06721_),
    .Z(_02445_));
 NOR4_X1 _15848_ (.A1(_02441_),
    .A2(_02442_),
    .A3(_02443_),
    .A4(_02445_),
    .ZN(_02446_));
 AOI21_X1 _15849_ (.A(_02437_),
    .B1(_02439_),
    .B2(_02446_),
    .ZN(_00362_));
 BUF_X2 _15850_ (.A(_10432_),
    .Z(_02447_));
 NAND2_X1 _15851_ (.A1(\dynamic_node_top.east_output.space.count_f[2] ),
    .A2(_02447_),
    .ZN(_02448_));
 BUF_X2 _15852_ (.A(_00057_),
    .Z(_02449_));
 NAND2_X1 _15853_ (.A1(_02449_),
    .A2(_02447_),
    .ZN(_02450_));
 OAI22_X1 _15854_ (.A1(_10566_),
    .A2(_02448_),
    .B1(_02450_),
    .B2(_10568_),
    .ZN(_02451_));
 BUF_X1 _15855_ (.A(_10426_),
    .Z(_02452_));
 NOR3_X1 _15856_ (.A1(_02452_),
    .A2(_10567_),
    .A3(_10565_),
    .ZN(_02453_));
 AOI21_X1 _15857_ (.A(_02453_),
    .B1(_10430_),
    .B2(_02452_),
    .ZN(_02454_));
 OAI21_X2 _15858_ (.A(_02447_),
    .B1(_02449_),
    .B2(\dynamic_node_top.east_output.space.count_f[2] ),
    .ZN(_02455_));
 AOI21_X1 _15859_ (.A(_02451_),
    .B1(_02454_),
    .B2(_02455_),
    .ZN(_02456_));
 NOR2_X1 _15860_ (.A1(_02404_),
    .A2(_02456_),
    .ZN(_00363_));
 CLKBUF_X2 _15861_ (.A(_10428_),
    .Z(_02457_));
 NAND4_X1 _15862_ (.A1(_10433_),
    .A2(_02457_),
    .A3(_02449_),
    .A4(_02447_),
    .ZN(_02458_));
 INV_X1 _15863_ (.A(_10433_),
    .ZN(_02459_));
 NAND2_X1 _15864_ (.A1(_10425_),
    .A2(_02459_),
    .ZN(_02460_));
 OAI21_X1 _15865_ (.A(_02458_),
    .B1(_02460_),
    .B2(_02448_),
    .ZN(_02461_));
 INV_X1 _15866_ (.A(_02457_),
    .ZN(_02462_));
 OAI21_X1 _15867_ (.A(_02460_),
    .B1(_02462_),
    .B2(_02459_),
    .ZN(_02463_));
 MUX2_X1 _15868_ (.A(_02463_),
    .B(\dynamic_node_top.east_output.space.count_f[1] ),
    .S(_02452_),
    .Z(_02464_));
 INV_X1 _15869_ (.A(_10431_),
    .ZN(_02465_));
 OAI22_X2 _15870_ (.A1(_10425_),
    .A2(_02448_),
    .B1(_02450_),
    .B2(_02457_),
    .ZN(_02466_));
 AOI221_X2 _15871_ (.A(_02461_),
    .B1(_02464_),
    .B2(_02455_),
    .C1(_02465_),
    .C2(_02466_),
    .ZN(_02467_));
 NOR2_X1 _15872_ (.A1(_02404_),
    .A2(_02467_),
    .ZN(_00364_));
 NAND2_X1 _15873_ (.A1(_10425_),
    .A2(_10434_),
    .ZN(_02468_));
 XOR2_X1 _15874_ (.A(_02449_),
    .B(_02468_),
    .Z(_02469_));
 MUX2_X1 _15875_ (.A(_02452_),
    .B(_02469_),
    .S(_02447_),
    .Z(_02470_));
 NAND2_X1 _15876_ (.A1(\dynamic_node_top.east_output.space.count_f[2] ),
    .A2(_02470_),
    .ZN(_02471_));
 INV_X1 _15877_ (.A(_02455_),
    .ZN(_02472_));
 XNOR2_X1 _15878_ (.A(_02449_),
    .B(_10436_),
    .ZN(_02473_));
 XNOR2_X1 _15879_ (.A(_02449_),
    .B(_10434_),
    .ZN(_02474_));
 AOI22_X1 _15880_ (.A1(_02457_),
    .A2(_02473_),
    .B1(_02474_),
    .B2(_10425_),
    .ZN(_02475_));
 OR3_X1 _15881_ (.A1(_02452_),
    .A2(_02472_),
    .A3(_02475_),
    .ZN(_02476_));
 NAND4_X1 _15882_ (.A1(_02457_),
    .A2(_02449_),
    .A3(_10436_),
    .A4(_02447_),
    .ZN(_02477_));
 AND2_X1 _15883_ (.A1(_06754_),
    .A2(_02477_),
    .ZN(_02478_));
 NAND3_X1 _15884_ (.A1(_02471_),
    .A2(_02476_),
    .A3(_02478_),
    .ZN(_00365_));
 NAND4_X1 _15885_ (.A1(_02467_),
    .A2(_02471_),
    .A3(_02476_),
    .A4(_02478_),
    .ZN(_00367_));
 NOR2_X1 _15886_ (.A1(_02456_),
    .A2(_00367_),
    .ZN(_00366_));
 CLKBUF_X3 _15887_ (.A(_06589_),
    .Z(_02479_));
 NOR2_X1 _15888_ (.A1(_02479_),
    .A2(_05308_),
    .ZN(_00368_));
 AND2_X1 _15889_ (.A1(_06892_),
    .A2(net295),
    .ZN(_00369_));
 CLKBUF_X3 _15890_ (.A(_06755_),
    .Z(_02480_));
 AND2_X1 _15891_ (.A1(_02480_),
    .A2(net259),
    .ZN(_00370_));
 AND2_X1 _15892_ (.A1(_02480_),
    .A2(net260),
    .ZN(_00371_));
 AND2_X1 _15893_ (.A1(_02480_),
    .A2(net261),
    .ZN(_00372_));
 AND2_X1 _15894_ (.A1(_02480_),
    .A2(net262),
    .ZN(_00373_));
 AND2_X1 _15895_ (.A1(_02480_),
    .A2(net263),
    .ZN(_00374_));
 AND2_X1 _15896_ (.A1(_02480_),
    .A2(net264),
    .ZN(_00375_));
 AND2_X1 _15897_ (.A1(_02480_),
    .A2(net265),
    .ZN(_00376_));
 AND2_X1 _15898_ (.A1(_02480_),
    .A2(net266),
    .ZN(_00377_));
 AND2_X1 _15899_ (.A1(_02480_),
    .A2(net267),
    .ZN(_00378_));
 AND2_X1 _15900_ (.A1(_02480_),
    .A2(net268),
    .ZN(_00379_));
 CLKBUF_X3 _15901_ (.A(_06880_),
    .Z(_02481_));
 AND2_X1 _15902_ (.A1(_02481_),
    .A2(net269),
    .ZN(_00380_));
 AND2_X1 _15903_ (.A1(_02481_),
    .A2(net270),
    .ZN(_00381_));
 AND2_X1 _15904_ (.A1(_02481_),
    .A2(net271),
    .ZN(_00382_));
 AND2_X1 _15905_ (.A1(_02481_),
    .A2(net272),
    .ZN(_00383_));
 AND2_X1 _15906_ (.A1(_02481_),
    .A2(net273),
    .ZN(_00384_));
 AND2_X1 _15907_ (.A1(_02481_),
    .A2(net274),
    .ZN(_00385_));
 AND2_X1 _15908_ (.A1(_02481_),
    .A2(net275),
    .ZN(_00386_));
 AND2_X1 _15909_ (.A1(_02481_),
    .A2(net276),
    .ZN(_00387_));
 AND2_X1 _15910_ (.A1(_02481_),
    .A2(net277),
    .ZN(_00388_));
 AND2_X1 _15911_ (.A1(_02481_),
    .A2(net278),
    .ZN(_00389_));
 CLKBUF_X2 _15912_ (.A(_06880_),
    .Z(_02482_));
 AND2_X1 _15913_ (.A1(_02482_),
    .A2(net279),
    .ZN(_00390_));
 AND2_X1 _15914_ (.A1(_02482_),
    .A2(net280),
    .ZN(_00391_));
 AND2_X1 _15915_ (.A1(_02482_),
    .A2(net281),
    .ZN(_00392_));
 AND2_X1 _15916_ (.A1(_02482_),
    .A2(net282),
    .ZN(_00393_));
 AND2_X1 _15917_ (.A1(_02482_),
    .A2(net283),
    .ZN(_00394_));
 AND2_X1 _15918_ (.A1(_02482_),
    .A2(net284),
    .ZN(_00395_));
 AND2_X1 _15919_ (.A1(_02482_),
    .A2(net285),
    .ZN(_00396_));
 AND2_X1 _15920_ (.A1(_02482_),
    .A2(net286),
    .ZN(_00397_));
 AND2_X1 _15921_ (.A1(_02482_),
    .A2(net287),
    .ZN(_00398_));
 AND2_X1 _15922_ (.A1(_02482_),
    .A2(net288),
    .ZN(_00399_));
 CLKBUF_X3 _15923_ (.A(_06880_),
    .Z(_02483_));
 MUX2_X1 _15924_ (.A(\dynamic_node_top.north_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.north_input.NIB.elements_in_array_next[0] ),
    .S(_10474_),
    .Z(_02484_));
 AND2_X1 _15925_ (.A1(_02483_),
    .A2(_02484_),
    .ZN(_00400_));
 NAND2_X1 _15926_ (.A1(_10167_),
    .A2(_10474_),
    .ZN(_02485_));
 OAI21_X1 _15927_ (.A(_02485_),
    .B1(_10474_),
    .B2(\dynamic_node_top.north_input.NIB.elements_in_array_f[1] ),
    .ZN(_02486_));
 NOR2_X1 _15928_ (.A1(_02479_),
    .A2(_02486_),
    .ZN(_00401_));
 XNOR2_X1 _15929_ (.A(_10477_),
    .B(_10166_),
    .ZN(_02487_));
 NAND2_X1 _15930_ (.A1(_10474_),
    .A2(_02487_),
    .ZN(_02488_));
 XOR2_X1 _15931_ (.A(\dynamic_node_top.north_input.NIB.elements_in_array_f[2] ),
    .B(_02488_),
    .Z(_02489_));
 NOR2_X1 _15932_ (.A1(_02479_),
    .A2(_02489_),
    .ZN(_00402_));
 MUX2_X1 _15933_ (.A(\dynamic_node_top.north_input.NIB.head_ptr_f[0] ),
    .B(\dynamic_node_top.north_input.NIB.head_ptr_next[0] ),
    .S(_02402_),
    .Z(_02490_));
 AND2_X1 _15934_ (.A1(_02483_),
    .A2(_02490_),
    .ZN(_00403_));
 NOR2_X2 _15935_ (.A1(_10473_),
    .A2(_10475_),
    .ZN(_02491_));
 MUX2_X1 _15936_ (.A(\dynamic_node_top.north_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.north_input.NIB.tail_ptr_next[0] ),
    .S(_02491_),
    .Z(_02492_));
 AND2_X1 _15937_ (.A1(_02483_),
    .A2(_02492_),
    .ZN(_00660_));
 MUX2_X1 _15938_ (.A(\dynamic_node_top.north_input.NIB.tail_ptr_f[1] ),
    .B(\dynamic_node_top.north_input.NIB.tail_ptr_next[1] ),
    .S(_02491_),
    .Z(_02493_));
 AND2_X1 _15939_ (.A1(_02483_),
    .A2(_02493_),
    .ZN(_00661_));
 NOR2_X1 _15940_ (.A1(_02479_),
    .A2(_10472_),
    .ZN(_00662_));
 INV_X2 _15941_ (.A(_05846_),
    .ZN(_02494_));
 NOR2_X1 _15942_ (.A1(_06909_),
    .A2(_02494_),
    .ZN(_02495_));
 AOI21_X1 _15943_ (.A(_02495_),
    .B1(_07087_),
    .B2(_06909_),
    .ZN(_02496_));
 NOR2_X1 _15944_ (.A1(_02479_),
    .A2(_02496_),
    .ZN(_00663_));
 AND2_X1 _15945_ (.A1(_02483_),
    .A2(_07091_),
    .ZN(_00664_));
 AND2_X1 _15946_ (.A1(_02483_),
    .A2(_07094_),
    .ZN(_00665_));
 OAI21_X1 _15947_ (.A(_06755_),
    .B1(_06909_),
    .B2(_05829_),
    .ZN(_02497_));
 AOI21_X1 _15948_ (.A(_02497_),
    .B1(_07098_),
    .B2(_06909_),
    .ZN(_00666_));
 NOR2_X1 _15949_ (.A1(_06909_),
    .A2(_05832_),
    .ZN(_02498_));
 NOR3_X1 _15950_ (.A1(_02420_),
    .A2(_02498_),
    .A3(_07102_),
    .ZN(_00667_));
 NOR2_X1 _15951_ (.A1(_02479_),
    .A2(_07118_),
    .ZN(_00668_));
 NOR2_X1 _15952_ (.A1(_02479_),
    .A2(_07115_),
    .ZN(_00669_));
 NOR2_X1 _15953_ (.A1(_02479_),
    .A2(_07111_),
    .ZN(_00670_));
 NOR3_X1 _15954_ (.A1(_02420_),
    .A2(_02496_),
    .A3(_07119_),
    .ZN(_00671_));
 NOR2_X1 _15955_ (.A1(_02479_),
    .A2(_06601_),
    .ZN(_00672_));
 OR3_X1 _15956_ (.A1(_05821_),
    .A2(_06510_),
    .A3(_06518_),
    .ZN(_02499_));
 AOI22_X2 _15957_ (.A1(_07021_),
    .A2(_06568_),
    .B1(_02499_),
    .B2(_06124_),
    .ZN(_02500_));
 INV_X1 _15958_ (.A(_06124_),
    .ZN(_02501_));
 AND2_X1 _15959_ (.A1(_06051_),
    .A2(_06084_),
    .ZN(_02502_));
 AOI22_X2 _15960_ (.A1(_06122_),
    .A2(_02501_),
    .B1(_02502_),
    .B2(net622),
    .ZN(_02503_));
 NOR2_X1 _15961_ (.A1(_05757_),
    .A2(_06568_),
    .ZN(_02504_));
 NOR2_X1 _15962_ (.A1(_06090_),
    .A2(_06120_),
    .ZN(_02505_));
 NOR3_X2 _15963_ (.A1(_06580_),
    .A2(_02504_),
    .A3(_02505_),
    .ZN(_02506_));
 OAI211_X2 _15964_ (.A(_06124_),
    .B(_02506_),
    .C1(_07038_),
    .C2(_05823_),
    .ZN(_02507_));
 NAND3_X1 _15965_ (.A1(_07038_),
    .A2(_06578_),
    .A3(_02506_),
    .ZN(_02508_));
 AOI211_X2 _15966_ (.A(_02500_),
    .B(_02503_),
    .C1(_02507_),
    .C2(_02508_),
    .ZN(_02509_));
 NAND2_X1 _15967_ (.A1(_06122_),
    .A2(_02502_),
    .ZN(_02510_));
 NOR2_X1 _15968_ (.A1(_06095_),
    .A2(net667),
    .ZN(_02511_));
 NAND4_X1 _15969_ (.A1(_07038_),
    .A2(_07021_),
    .A3(_06585_),
    .A4(_02511_),
    .ZN(_02512_));
 AOI21_X1 _15970_ (.A(_02510_),
    .B1(_02512_),
    .B2(_02501_),
    .ZN(_02513_));
 NOR3_X1 _15971_ (.A1(_06122_),
    .A2(_06124_),
    .A3(_02502_),
    .ZN(_02514_));
 NOR4_X1 _15972_ (.A1(_06573_),
    .A2(_02509_),
    .A3(_02513_),
    .A4(_02514_),
    .ZN(_00673_));
 BUF_X2 _15973_ (.A(_10543_),
    .Z(_02515_));
 NAND2_X1 _15974_ (.A1(\dynamic_node_top.north_output.space.count_f[2] ),
    .A2(_02515_),
    .ZN(_02516_));
 BUF_X2 _15975_ (.A(_00061_),
    .Z(_02517_));
 NAND2_X1 _15976_ (.A1(_02517_),
    .A2(_02515_),
    .ZN(_02518_));
 OAI22_X1 _15977_ (.A1(_10562_),
    .A2(_02516_),
    .B1(_02518_),
    .B2(_10564_),
    .ZN(_02519_));
 BUF_X1 _15978_ (.A(_10537_),
    .Z(_02520_));
 NOR3_X1 _15979_ (.A1(_02520_),
    .A2(_10563_),
    .A3(_10561_),
    .ZN(_02521_));
 AOI21_X1 _15980_ (.A(_02521_),
    .B1(_10541_),
    .B2(_02520_),
    .ZN(_02522_));
 OAI21_X2 _15981_ (.A(_02515_),
    .B1(_02517_),
    .B2(\dynamic_node_top.north_output.space.count_f[2] ),
    .ZN(_02523_));
 AOI21_X1 _15982_ (.A(_02519_),
    .B1(_02522_),
    .B2(_02523_),
    .ZN(_02524_));
 NOR2_X1 _15983_ (.A1(_02479_),
    .A2(_02524_),
    .ZN(_00674_));
 BUF_X4 _15984_ (.A(_06589_),
    .Z(_02525_));
 CLKBUF_X2 _15985_ (.A(_10539_),
    .Z(_02526_));
 NAND4_X1 _15986_ (.A1(_10544_),
    .A2(_02526_),
    .A3(_02517_),
    .A4(_02515_),
    .ZN(_02527_));
 INV_X1 _15987_ (.A(_10544_),
    .ZN(_02528_));
 NAND2_X1 _15988_ (.A1(_10536_),
    .A2(_02528_),
    .ZN(_02529_));
 OAI21_X1 _15989_ (.A(_02527_),
    .B1(_02529_),
    .B2(_02516_),
    .ZN(_02530_));
 INV_X1 _15990_ (.A(_02526_),
    .ZN(_02531_));
 OAI21_X1 _15991_ (.A(_02529_),
    .B1(_02531_),
    .B2(_02528_),
    .ZN(_02532_));
 MUX2_X1 _15992_ (.A(_02532_),
    .B(\dynamic_node_top.north_output.space.count_f[1] ),
    .S(_02520_),
    .Z(_02533_));
 INV_X1 _15993_ (.A(_10542_),
    .ZN(_02534_));
 OAI22_X2 _15994_ (.A1(_10536_),
    .A2(_02516_),
    .B1(_02518_),
    .B2(_02526_),
    .ZN(_02535_));
 AOI221_X2 _15995_ (.A(_02530_),
    .B1(_02533_),
    .B2(_02523_),
    .C1(_02534_),
    .C2(_02535_),
    .ZN(_02536_));
 NOR2_X1 _15996_ (.A1(_02525_),
    .A2(_02536_),
    .ZN(_00675_));
 NAND2_X1 _15997_ (.A1(_10536_),
    .A2(_10545_),
    .ZN(_02537_));
 XOR2_X1 _15998_ (.A(_02517_),
    .B(_02537_),
    .Z(_02538_));
 MUX2_X1 _15999_ (.A(_02520_),
    .B(_02538_),
    .S(_02515_),
    .Z(_02539_));
 NAND2_X1 _16000_ (.A1(\dynamic_node_top.north_output.space.count_f[2] ),
    .A2(_02539_),
    .ZN(_02540_));
 INV_X1 _16001_ (.A(_02523_),
    .ZN(_02541_));
 XNOR2_X1 _16002_ (.A(_02517_),
    .B(_10547_),
    .ZN(_02542_));
 XNOR2_X1 _16003_ (.A(_02517_),
    .B(_10545_),
    .ZN(_02543_));
 AOI22_X1 _16004_ (.A1(_02526_),
    .A2(_02542_),
    .B1(_02543_),
    .B2(_10536_),
    .ZN(_02544_));
 OR3_X1 _16005_ (.A1(_02520_),
    .A2(_02541_),
    .A3(_02544_),
    .ZN(_02545_));
 NAND4_X1 _16006_ (.A1(_02526_),
    .A2(_02517_),
    .A3(_10547_),
    .A4(_02515_),
    .ZN(_02546_));
 AND2_X1 _16007_ (.A1(_06754_),
    .A2(_02546_),
    .ZN(_02547_));
 NAND3_X1 _16008_ (.A1(_02540_),
    .A2(_02545_),
    .A3(_02547_),
    .ZN(_00676_));
 NAND4_X1 _16009_ (.A1(_02536_),
    .A2(_02540_),
    .A3(_02545_),
    .A4(_02547_),
    .ZN(_00678_));
 NOR2_X1 _16010_ (.A1(_02524_),
    .A2(_00678_),
    .ZN(_00677_));
 AND2_X1 _16011_ (.A1(_06892_),
    .A2(net622),
    .ZN(_00679_));
 AND2_X1 _16012_ (.A1(_02483_),
    .A2(net296),
    .ZN(_00680_));
 BUF_X2 _16013_ (.A(_10459_),
    .Z(_02548_));
 MUX2_X1 _16014_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.proc_input.NIB.elements_in_array_next[0] ),
    .S(_02548_),
    .Z(_02549_));
 AND2_X1 _16015_ (.A1(_02483_),
    .A2(_02549_),
    .ZN(_00681_));
 NAND2_X1 _16016_ (.A1(_10171_),
    .A2(_02548_),
    .ZN(_02550_));
 OAI21_X1 _16017_ (.A(_02550_),
    .B1(_02548_),
    .B2(\dynamic_node_top.proc_input.NIB.elements_in_array_f[1] ),
    .ZN(_02551_));
 NOR2_X1 _16018_ (.A1(_02525_),
    .A2(_02551_),
    .ZN(_00682_));
 XNOR2_X1 _16019_ (.A(_10170_),
    .B(_10573_),
    .ZN(_02552_));
 MUX2_X1 _16020_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[2] ),
    .B(_02552_),
    .S(_02548_),
    .Z(_02553_));
 AND2_X1 _16021_ (.A1(_02483_),
    .A2(_02553_),
    .ZN(_00683_));
 INV_X1 _16022_ (.A(_10572_),
    .ZN(_02554_));
 AOI21_X1 _16023_ (.A(_10570_),
    .B1(_10571_),
    .B2(\dynamic_node_top.proc_input.NIB.elements_in_array_f[0] ),
    .ZN(_02555_));
 INV_X1 _16024_ (.A(_10573_),
    .ZN(_02556_));
 OAI21_X1 _16025_ (.A(_02554_),
    .B1(_02555_),
    .B2(_02556_),
    .ZN(_02557_));
 XOR2_X1 _16026_ (.A(_10575_),
    .B(_02557_),
    .Z(_02558_));
 MUX2_X1 _16027_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[3] ),
    .B(_02558_),
    .S(_02548_),
    .Z(_02559_));
 AND2_X1 _16028_ (.A1(_02483_),
    .A2(_02559_),
    .ZN(_00684_));
 OAI21_X1 _16029_ (.A(_02554_),
    .B1(_02556_),
    .B2(_10170_),
    .ZN(_02560_));
 AOI21_X1 _16030_ (.A(_10574_),
    .B1(_10575_),
    .B2(_02560_),
    .ZN(_02561_));
 XNOR2_X1 _16031_ (.A(_10569_),
    .B(_02561_),
    .ZN(_02562_));
 NAND2_X1 _16032_ (.A1(_02548_),
    .A2(_02562_),
    .ZN(_02563_));
 XOR2_X1 _16033_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[4] ),
    .B(_02563_),
    .Z(_02564_));
 NOR2_X1 _16034_ (.A1(_02525_),
    .A2(_02564_),
    .ZN(_00685_));
 BUF_X4 _16035_ (.A(_06880_),
    .Z(_02565_));
 MUX2_X1 _16036_ (.A(\dynamic_node_top.proc_input.NIB.head_ptr_f[0] ),
    .B(\dynamic_node_top.proc_input.NIB.head_ptr_next[0] ),
    .S(_02395_),
    .Z(_02566_));
 AND2_X1 _16037_ (.A1(_02565_),
    .A2(_02566_),
    .ZN(_00686_));
 NOR2_X4 _16038_ (.A1(_10461_),
    .A2(_10458_),
    .ZN(_02567_));
 MUX2_X1 _16039_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.proc_input.NIB.tail_ptr_next[0] ),
    .S(_02567_),
    .Z(_02568_));
 AND2_X1 _16040_ (.A1(_02565_),
    .A2(_02568_),
    .ZN(_01711_));
 MUX2_X1 _16041_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_f[1] ),
    .B(\dynamic_node_top.proc_input.NIB.tail_ptr_next[1] ),
    .S(_02567_),
    .Z(_02569_));
 AND2_X1 _16042_ (.A1(_02565_),
    .A2(_02569_),
    .ZN(_01712_));
 NAND2_X1 _16043_ (.A1(_07895_),
    .A2(_02567_),
    .ZN(_02570_));
 XNOR2_X1 _16044_ (.A(_07883_),
    .B(_02570_),
    .ZN(_02571_));
 NOR2_X1 _16045_ (.A1(_02525_),
    .A2(_02571_),
    .ZN(_01713_));
 NAND4_X1 _16046_ (.A1(_07747_),
    .A2(\dynamic_node_top.proc_input.NIB.tail_ptr_f[1] ),
    .A3(\dynamic_node_top.proc_input.NIB.tail_ptr_f[0] ),
    .A4(_02567_),
    .ZN(_02572_));
 XOR2_X1 _16047_ (.A(_07746_),
    .B(_02572_),
    .Z(_02573_));
 NOR2_X1 _16048_ (.A1(_02525_),
    .A2(_02573_),
    .ZN(_01714_));
 NOR2_X1 _16049_ (.A1(_02525_),
    .A2(_10456_),
    .ZN(_01715_));
 NOR2_X1 _16050_ (.A1(_02525_),
    .A2(_07133_),
    .ZN(_01716_));
 NOR2_X1 _16051_ (.A1(_02525_),
    .A2(_07157_),
    .ZN(_01717_));
 NOR2_X1 _16052_ (.A1(_02525_),
    .A2(_07138_),
    .ZN(_01718_));
 AND2_X1 _16053_ (.A1(_02565_),
    .A2(_07151_),
    .ZN(_01719_));
 NOR2_X1 _16054_ (.A1(_02525_),
    .A2(_07159_),
    .ZN(_01720_));
 AND2_X1 _16055_ (.A1(_02565_),
    .A2(_07149_),
    .ZN(_01721_));
 BUF_X4 _16056_ (.A(_06589_),
    .Z(_02574_));
 NOR2_X1 _16057_ (.A1(_02574_),
    .A2(_07142_),
    .ZN(_01722_));
 NOR2_X1 _16058_ (.A1(_02574_),
    .A2(_07163_),
    .ZN(_01723_));
 NOR3_X1 _16059_ (.A1(_02420_),
    .A2(_07133_),
    .A3(_07164_),
    .ZN(_01724_));
 NOR2_X1 _16060_ (.A1(_02574_),
    .A2(_06050_),
    .ZN(_01725_));
 OR3_X1 _16061_ (.A1(_05697_),
    .A2(_06931_),
    .A3(_06938_),
    .ZN(_02575_));
 NAND4_X1 _16062_ (.A1(_06987_),
    .A2(_06975_),
    .A3(_06920_),
    .A4(_06948_),
    .ZN(_02576_));
 NOR4_X2 _16063_ (.A1(_05610_),
    .A2(_06936_),
    .A3(_06937_),
    .A4(_02576_),
    .ZN(_02577_));
 OAI211_X2 _16064_ (.A(_05697_),
    .B(_02577_),
    .C1(_06945_),
    .C2(_06944_),
    .ZN(_02578_));
 NAND3_X1 _16065_ (.A1(_05697_),
    .A2(_06931_),
    .A3(_06938_),
    .ZN(_02579_));
 NAND4_X1 _16066_ (.A1(_06755_),
    .A2(_02575_),
    .A3(_02578_),
    .A4(_02579_),
    .ZN(_02580_));
 INV_X1 _16067_ (.A(_06931_),
    .ZN(_02581_));
 AOI21_X1 _16068_ (.A(_02581_),
    .B1(net744),
    .B2(_06938_),
    .ZN(_02582_));
 NAND2_X1 _16069_ (.A1(_05595_),
    .A2(_06931_),
    .ZN(_02583_));
 AOI22_X1 _16070_ (.A1(_06934_),
    .A2(_06914_),
    .B1(_06926_),
    .B2(_02583_),
    .ZN(_02584_));
 OAI21_X1 _16071_ (.A(_06931_),
    .B1(_05696_),
    .B2(_05603_),
    .ZN(_02585_));
 OAI21_X1 _16072_ (.A(_02585_),
    .B1(_06914_),
    .B2(_06987_),
    .ZN(_02586_));
 NAND2_X1 _16073_ (.A1(_02584_),
    .A2(_02586_),
    .ZN(_02587_));
 NAND2_X1 _16074_ (.A1(_06787_),
    .A2(_06789_),
    .ZN(_02588_));
 INV_X1 _16075_ (.A(_06907_),
    .ZN(_02589_));
 OAI33_X1 _16076_ (.A1(_06163_),
    .A2(_06740_),
    .A3(_06944_),
    .B1(_02588_),
    .B2(_02589_),
    .B3(_06905_),
    .ZN(_02590_));
 AOI211_X2 _16077_ (.A(_02582_),
    .B(_02587_),
    .C1(_02581_),
    .C2(_02590_),
    .ZN(_02591_));
 OR2_X1 _16078_ (.A1(_05605_),
    .A2(_06908_),
    .ZN(_02592_));
 NAND3_X1 _16079_ (.A1(net744),
    .A2(_06938_),
    .A3(_02592_),
    .ZN(_02593_));
 NOR3_X1 _16080_ (.A1(_06916_),
    .A2(_06944_),
    .A3(_06945_),
    .ZN(_02594_));
 OAI21_X1 _16081_ (.A(_07124_),
    .B1(_02593_),
    .B2(_02594_),
    .ZN(_02595_));
 AOI21_X1 _16082_ (.A(_02580_),
    .B1(_02591_),
    .B2(_02595_),
    .ZN(_01726_));
 BUF_X2 _16083_ (.A(_10525_),
    .Z(_02596_));
 NAND2_X1 _16084_ (.A1(\dynamic_node_top.proc_output.space.count_f[2] ),
    .A2(_02596_),
    .ZN(_02597_));
 BUF_X2 _16085_ (.A(_00060_),
    .Z(_02598_));
 NAND2_X1 _16086_ (.A1(_02598_),
    .A2(_02596_),
    .ZN(_02599_));
 OAI22_X1 _16087_ (.A1(_10554_),
    .A2(_02597_),
    .B1(_02599_),
    .B2(_10556_),
    .ZN(_02600_));
 BUF_X1 _16088_ (.A(_10519_),
    .Z(_02601_));
 NOR3_X1 _16089_ (.A1(_02601_),
    .A2(_10555_),
    .A3(_10553_),
    .ZN(_02602_));
 AOI21_X1 _16090_ (.A(_02602_),
    .B1(_10523_),
    .B2(_02601_),
    .ZN(_02603_));
 OAI21_X2 _16091_ (.A(_02596_),
    .B1(_02598_),
    .B2(\dynamic_node_top.proc_output.space.count_f[2] ),
    .ZN(_02604_));
 AOI21_X1 _16092_ (.A(_02600_),
    .B1(_02603_),
    .B2(_02604_),
    .ZN(_02605_));
 NOR2_X1 _16093_ (.A1(_02574_),
    .A2(_02605_),
    .ZN(_01727_));
 CLKBUF_X2 _16094_ (.A(_10521_),
    .Z(_02606_));
 NAND4_X1 _16095_ (.A1(_10526_),
    .A2(_02606_),
    .A3(_02598_),
    .A4(_02596_),
    .ZN(_02607_));
 INV_X1 _16096_ (.A(_10526_),
    .ZN(_02608_));
 NAND2_X1 _16097_ (.A1(_10518_),
    .A2(_02608_),
    .ZN(_02609_));
 OAI21_X1 _16098_ (.A(_02607_),
    .B1(_02609_),
    .B2(_02597_),
    .ZN(_02610_));
 INV_X1 _16099_ (.A(_02606_),
    .ZN(_02611_));
 OAI21_X1 _16100_ (.A(_02609_),
    .B1(_02611_),
    .B2(_02608_),
    .ZN(_02612_));
 MUX2_X1 _16101_ (.A(_02612_),
    .B(\dynamic_node_top.proc_output.space.count_f[1] ),
    .S(_02601_),
    .Z(_02613_));
 INV_X1 _16102_ (.A(_10524_),
    .ZN(_02614_));
 OAI22_X2 _16103_ (.A1(_10518_),
    .A2(_02597_),
    .B1(_02599_),
    .B2(_02606_),
    .ZN(_02615_));
 AOI221_X2 _16104_ (.A(_02610_),
    .B1(_02613_),
    .B2(_02604_),
    .C1(_02614_),
    .C2(_02615_),
    .ZN(_02616_));
 NOR2_X1 _16105_ (.A1(_02574_),
    .A2(_02616_),
    .ZN(_01728_));
 NAND2_X1 _16106_ (.A1(_10518_),
    .A2(_10527_),
    .ZN(_02617_));
 XOR2_X1 _16107_ (.A(_02598_),
    .B(_02617_),
    .Z(_02618_));
 MUX2_X1 _16108_ (.A(_02601_),
    .B(_02618_),
    .S(_02596_),
    .Z(_02619_));
 NAND2_X1 _16109_ (.A1(\dynamic_node_top.proc_output.space.count_f[2] ),
    .A2(_02619_),
    .ZN(_02620_));
 INV_X1 _16110_ (.A(_02604_),
    .ZN(_02621_));
 XNOR2_X1 _16111_ (.A(_02598_),
    .B(_10529_),
    .ZN(_02622_));
 XNOR2_X1 _16112_ (.A(_02598_),
    .B(_10527_),
    .ZN(_02623_));
 AOI22_X1 _16113_ (.A1(_02606_),
    .A2(_02622_),
    .B1(_02623_),
    .B2(_10518_),
    .ZN(_02624_));
 OR3_X1 _16114_ (.A1(_02601_),
    .A2(_02621_),
    .A3(_02624_),
    .ZN(_02625_));
 NAND4_X1 _16115_ (.A1(_02606_),
    .A2(_02598_),
    .A3(_10529_),
    .A4(_02596_),
    .ZN(_02626_));
 AND2_X1 _16116_ (.A1(_06754_),
    .A2(_02626_),
    .ZN(_02627_));
 NAND3_X1 _16117_ (.A1(_02620_),
    .A2(_02625_),
    .A3(_02627_),
    .ZN(_01729_));
 NAND4_X1 _16118_ (.A1(_02616_),
    .A2(_02620_),
    .A3(_02625_),
    .A4(_02627_),
    .ZN(_01731_));
 NOR2_X1 _16119_ (.A1(_02605_),
    .A2(_01731_),
    .ZN(_01730_));
 AND2_X1 _16120_ (.A1(_02565_),
    .A2(net744),
    .ZN(_01732_));
 AND2_X1 _16121_ (.A1(_02565_),
    .A2(net297),
    .ZN(_01733_));
 MUX2_X1 _16122_ (.A(\dynamic_node_top.south_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.south_input.NIB.elements_in_array_next[0] ),
    .S(_10466_),
    .Z(_02628_));
 AND2_X1 _16123_ (.A1(_02565_),
    .A2(_02628_),
    .ZN(_01734_));
 NAND2_X1 _16124_ (.A1(_10174_),
    .A2(_10466_),
    .ZN(_02629_));
 OAI21_X1 _16125_ (.A(_02629_),
    .B1(_10466_),
    .B2(\dynamic_node_top.south_input.NIB.elements_in_array_f[1] ),
    .ZN(_02630_));
 NOR2_X1 _16126_ (.A1(_02574_),
    .A2(_02630_),
    .ZN(_01735_));
 XNOR2_X1 _16127_ (.A(_10469_),
    .B(_10173_),
    .ZN(_02631_));
 NAND2_X1 _16128_ (.A1(_10466_),
    .A2(_02631_),
    .ZN(_02632_));
 XOR2_X1 _16129_ (.A(\dynamic_node_top.south_input.NIB.elements_in_array_f[2] ),
    .B(_02632_),
    .Z(_02633_));
 NOR2_X1 _16130_ (.A1(_02574_),
    .A2(_02633_),
    .ZN(_01736_));
 MUX2_X1 _16131_ (.A(\dynamic_node_top.south_input.NIB.head_ptr_f[0] ),
    .B(\dynamic_node_top.south_input.NIB.head_ptr_next[0] ),
    .S(_02387_),
    .Z(_02634_));
 AND2_X1 _16132_ (.A1(_02565_),
    .A2(_02634_),
    .ZN(_01737_));
 NOR2_X4 _16133_ (.A1(_10465_),
    .A2(_10467_),
    .ZN(_02635_));
 MUX2_X1 _16134_ (.A(\dynamic_node_top.south_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.south_input.NIB.tail_ptr_next[0] ),
    .S(_02635_),
    .Z(_02636_));
 AND2_X1 _16135_ (.A1(_02565_),
    .A2(_02636_),
    .ZN(_01994_));
 BUF_X4 _16136_ (.A(_06880_),
    .Z(_02637_));
 MUX2_X1 _16137_ (.A(\dynamic_node_top.south_input.NIB.tail_ptr_f[1] ),
    .B(\dynamic_node_top.south_input.NIB.tail_ptr_next[1] ),
    .S(_02635_),
    .Z(_02638_));
 AND2_X1 _16138_ (.A1(_02637_),
    .A2(_02638_),
    .ZN(_01995_));
 NOR2_X1 _16139_ (.A1(_02574_),
    .A2(_10464_),
    .ZN(_01996_));
 AND2_X1 _16140_ (.A1(_06754_),
    .A2(_07173_),
    .ZN(_01997_));
 NOR2_X1 _16141_ (.A1(_06052_),
    .A2(\dynamic_node_top.south_input.control.count_f[1] ),
    .ZN(_02639_));
 AOI221_X1 _16142_ (.A(_02639_),
    .B1(_10516_),
    .B2(_06052_),
    .C1(\dynamic_node_top.south_input.control.header_last_temp ),
    .C2(_05170_),
    .ZN(_02640_));
 AOI21_X1 _16143_ (.A(_02640_),
    .B1(_06060_),
    .B2(_06103_),
    .ZN(_02641_));
 NOR2_X1 _16144_ (.A1(_02574_),
    .A2(_02641_),
    .ZN(_01998_));
 NAND2_X1 _16145_ (.A1(_06103_),
    .A2(_06064_),
    .ZN(_02642_));
 XNOR2_X1 _16146_ (.A(_07175_),
    .B(_07176_),
    .ZN(_02643_));
 NAND2_X1 _16147_ (.A1(_06096_),
    .A2(_02643_),
    .ZN(_02644_));
 AOI21_X1 _16148_ (.A(_06573_),
    .B1(_02642_),
    .B2(_02644_),
    .ZN(_01999_));
 NOR2_X1 _16149_ (.A1(_06096_),
    .A2(_06067_),
    .ZN(_02645_));
 NOR2_X1 _16150_ (.A1(_06103_),
    .A2(_07182_),
    .ZN(_02646_));
 NOR3_X1 _16151_ (.A1(_02420_),
    .A2(_02645_),
    .A3(_02646_),
    .ZN(_02000_));
 INV_X1 _16152_ (.A(_06057_),
    .ZN(_02647_));
 NOR3_X1 _16153_ (.A1(_06573_),
    .A2(_02647_),
    .A3(_07179_),
    .ZN(_02001_));
 NOR2_X1 _16154_ (.A1(_02574_),
    .A2(_07198_),
    .ZN(_02002_));
 BUF_X4 _16155_ (.A(_06589_),
    .Z(_02648_));
 NOR2_X1 _16156_ (.A1(_02648_),
    .A2(_07195_),
    .ZN(_02003_));
 AND2_X1 _16157_ (.A1(_02637_),
    .A2(_07191_),
    .ZN(_02004_));
 INV_X1 _16158_ (.A(_01997_),
    .ZN(_02649_));
 NOR4_X1 _16159_ (.A1(_07187_),
    .A2(_07191_),
    .A3(_07199_),
    .A4(_02649_),
    .ZN(_02005_));
 NOR2_X1 _16160_ (.A1(_02648_),
    .A2(_06083_),
    .ZN(_02006_));
 AND2_X1 _16161_ (.A1(_05454_),
    .A2(_06812_),
    .ZN(_02650_));
 NAND2_X1 _16162_ (.A1(_06818_),
    .A2(_02650_),
    .ZN(_02651_));
 OR3_X1 _16163_ (.A1(_05454_),
    .A2(_06812_),
    .A3(_06818_),
    .ZN(_02652_));
 NAND3_X1 _16164_ (.A1(_06880_),
    .A2(_02651_),
    .A3(_02652_),
    .ZN(_02653_));
 OR4_X1 _16165_ (.A1(_06865_),
    .A2(_06802_),
    .A3(_06828_),
    .A4(_06881_),
    .ZN(_02654_));
 NAND4_X1 _16166_ (.A1(_05454_),
    .A2(_05344_),
    .A3(_06856_),
    .A4(_06818_),
    .ZN(_02655_));
 NOR2_X1 _16167_ (.A1(_02654_),
    .A2(_02655_),
    .ZN(_02656_));
 AOI22_X1 _16168_ (.A1(_05454_),
    .A2(_06813_),
    .B1(_05344_),
    .B2(_06818_),
    .ZN(_02657_));
 NAND2_X1 _16169_ (.A1(_05452_),
    .A2(_02650_),
    .ZN(_02658_));
 OAI221_X1 _16170_ (.A(_02658_),
    .B1(_06851_),
    .B2(_06806_),
    .C1(_05338_),
    .C2(net680),
    .ZN(_02659_));
 NOR3_X1 _16171_ (.A1(_05330_),
    .A2(_06613_),
    .A3(_06801_),
    .ZN(_02660_));
 NOR3_X1 _16172_ (.A1(_02657_),
    .A2(_02659_),
    .A3(_02660_),
    .ZN(_02661_));
 OAI221_X1 _16173_ (.A(_06812_),
    .B1(_06798_),
    .B2(_05331_),
    .C1(_06876_),
    .C2(_05329_),
    .ZN(_02662_));
 OAI21_X1 _16174_ (.A(_02662_),
    .B1(_02654_),
    .B2(_06856_),
    .ZN(_02663_));
 AOI211_X2 _16175_ (.A(_02653_),
    .B(_02656_),
    .C1(_02661_),
    .C2(_02663_),
    .ZN(_02007_));
 BUF_X2 _16176_ (.A(_10491_),
    .Z(_02664_));
 NAND2_X1 _16177_ (.A1(\dynamic_node_top.south_output.space.count_f[2] ),
    .A2(_02664_),
    .ZN(_02665_));
 BUF_X2 _16178_ (.A(_00059_),
    .Z(_02666_));
 NAND2_X1 _16179_ (.A1(_02666_),
    .A2(_02664_),
    .ZN(_02667_));
 OAI22_X1 _16180_ (.A1(_10558_),
    .A2(_02665_),
    .B1(_02667_),
    .B2(_10560_),
    .ZN(_02668_));
 BUF_X1 _16181_ (.A(_10485_),
    .Z(_02669_));
 NOR3_X1 _16182_ (.A1(_02669_),
    .A2(_10559_),
    .A3(_10557_),
    .ZN(_02670_));
 AOI21_X1 _16183_ (.A(_02670_),
    .B1(_10489_),
    .B2(_02669_),
    .ZN(_02671_));
 OAI21_X2 _16184_ (.A(_02664_),
    .B1(_02666_),
    .B2(\dynamic_node_top.south_output.space.count_f[2] ),
    .ZN(_02672_));
 AOI21_X1 _16185_ (.A(_02668_),
    .B1(_02671_),
    .B2(_02672_),
    .ZN(_02673_));
 NOR2_X1 _16186_ (.A1(_02648_),
    .A2(_02673_),
    .ZN(_02008_));
 CLKBUF_X2 _16187_ (.A(_10487_),
    .Z(_02674_));
 NAND4_X1 _16188_ (.A1(_10492_),
    .A2(_02674_),
    .A3(_02666_),
    .A4(_02664_),
    .ZN(_02675_));
 INV_X1 _16189_ (.A(_10492_),
    .ZN(_02676_));
 NAND2_X1 _16190_ (.A1(_10484_),
    .A2(_02676_),
    .ZN(_02677_));
 OAI21_X1 _16191_ (.A(_02675_),
    .B1(_02677_),
    .B2(_02665_),
    .ZN(_02678_));
 INV_X1 _16192_ (.A(_02674_),
    .ZN(_02679_));
 OAI21_X1 _16193_ (.A(_02677_),
    .B1(_02679_),
    .B2(_02676_),
    .ZN(_02680_));
 MUX2_X1 _16194_ (.A(_02680_),
    .B(\dynamic_node_top.south_output.space.count_f[1] ),
    .S(_02669_),
    .Z(_02681_));
 INV_X1 _16195_ (.A(_10490_),
    .ZN(_02682_));
 OAI22_X2 _16196_ (.A1(_10484_),
    .A2(_02665_),
    .B1(_02667_),
    .B2(_02674_),
    .ZN(_02683_));
 AOI221_X2 _16197_ (.A(_02678_),
    .B1(_02681_),
    .B2(_02672_),
    .C1(_02682_),
    .C2(_02683_),
    .ZN(_02684_));
 NOR2_X1 _16198_ (.A1(_02648_),
    .A2(_02684_),
    .ZN(_02009_));
 NAND2_X1 _16199_ (.A1(_10484_),
    .A2(_10493_),
    .ZN(_02685_));
 XOR2_X1 _16200_ (.A(_02666_),
    .B(_02685_),
    .Z(_02686_));
 MUX2_X1 _16201_ (.A(_02669_),
    .B(_02686_),
    .S(_02664_),
    .Z(_02687_));
 NAND2_X1 _16202_ (.A1(\dynamic_node_top.south_output.space.count_f[2] ),
    .A2(_02687_),
    .ZN(_02688_));
 INV_X1 _16203_ (.A(_02672_),
    .ZN(_02689_));
 XNOR2_X1 _16204_ (.A(_02666_),
    .B(_10495_),
    .ZN(_02690_));
 XNOR2_X1 _16205_ (.A(_02666_),
    .B(_10493_),
    .ZN(_02691_));
 AOI22_X1 _16206_ (.A1(_02674_),
    .A2(_02690_),
    .B1(_02691_),
    .B2(_10484_),
    .ZN(_02692_));
 OR3_X1 _16207_ (.A1(_02669_),
    .A2(_02689_),
    .A3(_02692_),
    .ZN(_02693_));
 NAND4_X1 _16208_ (.A1(_02674_),
    .A2(_02666_),
    .A3(_10495_),
    .A4(_02664_),
    .ZN(_02694_));
 AND2_X1 _16209_ (.A1(_06754_),
    .A2(_02694_),
    .ZN(_02695_));
 NAND3_X1 _16210_ (.A1(_02688_),
    .A2(_02693_),
    .A3(_02695_),
    .ZN(_02010_));
 NAND4_X1 _16211_ (.A1(_02684_),
    .A2(_02688_),
    .A3(_02693_),
    .A4(_02695_),
    .ZN(_02012_));
 NOR2_X1 _16212_ (.A1(_02673_),
    .A2(_02012_),
    .ZN(_02011_));
 AND2_X1 _16213_ (.A1(_02637_),
    .A2(net1),
    .ZN(_02013_));
 AND2_X1 _16214_ (.A1(_02637_),
    .A2(net298),
    .ZN(_02014_));
 MUX2_X1 _16215_ (.A(\dynamic_node_top.west_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.west_input.NIB.elements_in_array_next[0] ),
    .S(_10500_),
    .Z(_02696_));
 AND2_X1 _16216_ (.A1(_02637_),
    .A2(_02696_),
    .ZN(_02015_));
 NAND2_X1 _16217_ (.A1(_10177_),
    .A2(_10500_),
    .ZN(_02697_));
 OAI21_X1 _16218_ (.A(_02697_),
    .B1(_10500_),
    .B2(\dynamic_node_top.west_input.NIB.elements_in_array_f[1] ),
    .ZN(_02698_));
 NOR2_X1 _16219_ (.A1(_02648_),
    .A2(_02698_),
    .ZN(_02016_));
 XNOR2_X1 _16220_ (.A(_10503_),
    .B(_10176_),
    .ZN(_02699_));
 NAND2_X1 _16221_ (.A1(_10500_),
    .A2(_02699_),
    .ZN(_02700_));
 XOR2_X1 _16222_ (.A(\dynamic_node_top.west_input.NIB.elements_in_array_f[2] ),
    .B(_02700_),
    .Z(_02701_));
 NOR2_X1 _16223_ (.A1(_02648_),
    .A2(_02701_),
    .ZN(_02017_));
 MUX2_X1 _16224_ (.A(\dynamic_node_top.west_input.NIB.head_ptr_f[0] ),
    .B(\dynamic_node_top.west_input.NIB.head_ptr_next[0] ),
    .S(_02383_),
    .Z(_02702_));
 AND2_X1 _16225_ (.A1(_02637_),
    .A2(_02702_),
    .ZN(_02018_));
 NOR2_X2 _16226_ (.A1(_10501_),
    .A2(_10499_),
    .ZN(_02703_));
 MUX2_X1 _16227_ (.A(\dynamic_node_top.west_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.west_input.NIB.tail_ptr_next[0] ),
    .S(_02703_),
    .Z(_02704_));
 AND2_X1 _16228_ (.A1(_02637_),
    .A2(_02704_),
    .ZN(_02275_));
 MUX2_X1 _16229_ (.A(\dynamic_node_top.west_input.NIB.tail_ptr_f[1] ),
    .B(\dynamic_node_top.west_input.NIB.tail_ptr_next[1] ),
    .S(_02703_),
    .Z(_02705_));
 AND2_X1 _16230_ (.A1(_02637_),
    .A2(_02705_),
    .ZN(_02276_));
 NOR2_X1 _16231_ (.A1(_02648_),
    .A2(_10498_),
    .ZN(_02277_));
 AND2_X1 _16232_ (.A1(_06754_),
    .A2(_07048_),
    .ZN(_02278_));
 NOR2_X1 _16233_ (.A1(_05818_),
    .A2(\dynamic_node_top.west_input.control.count_f[1] ),
    .ZN(_02706_));
 AOI221_X1 _16234_ (.A(_02706_),
    .B1(_10482_),
    .B2(_05818_),
    .C1(\dynamic_node_top.west_input.control.header_last_temp ),
    .C2(_05175_),
    .ZN(_02707_));
 AOI21_X1 _16235_ (.A(_02707_),
    .B1(_05796_),
    .B2(_06701_),
    .ZN(_02708_));
 NOR2_X1 _16236_ (.A1(_02648_),
    .A2(_02708_),
    .ZN(_02279_));
 NOR2_X1 _16237_ (.A1(_06613_),
    .A2(_05799_),
    .ZN(_02709_));
 XNOR2_X1 _16238_ (.A(_07049_),
    .B(_07050_),
    .ZN(_02710_));
 NOR2_X1 _16239_ (.A1(_06701_),
    .A2(_02710_),
    .ZN(_02711_));
 NOR3_X1 _16240_ (.A1(_06573_),
    .A2(_02709_),
    .A3(_02711_),
    .ZN(_02280_));
 NOR2_X1 _16241_ (.A1(_06613_),
    .A2(_05802_),
    .ZN(_02712_));
 NOR2_X1 _16242_ (.A1(_06701_),
    .A2(_07056_),
    .ZN(_02713_));
 NOR3_X1 _16243_ (.A1(_06573_),
    .A2(_02712_),
    .A3(_02713_),
    .ZN(_02281_));
 NOR3_X1 _16244_ (.A1(_06573_),
    .A2(_05793_),
    .A3(_07053_),
    .ZN(_02282_));
 NOR2_X1 _16245_ (.A1(_02648_),
    .A2(_07072_),
    .ZN(_02283_));
 NOR2_X1 _16246_ (.A1(_02648_),
    .A2(_07069_),
    .ZN(_02284_));
 AND2_X1 _16247_ (.A1(_02637_),
    .A2(_07065_),
    .ZN(_02285_));
 INV_X1 _16248_ (.A(_02278_),
    .ZN(_02714_));
 NOR4_X1 _16249_ (.A1(_07061_),
    .A2(_07065_),
    .A3(_07073_),
    .A4(_02714_),
    .ZN(_02286_));
 NOR2_X1 _16250_ (.A1(_02420_),
    .A2(_06713_),
    .ZN(_02287_));
 NAND3_X1 _16251_ (.A1(_06755_),
    .A2(\dynamic_node_top.west_output.control.planned_f ),
    .A3(_06605_),
    .ZN(_02715_));
 OR3_X1 _16252_ (.A1(_05487_),
    .A2(_05590_),
    .A3(_06605_),
    .ZN(_02716_));
 NOR4_X1 _16253_ (.A1(_06618_),
    .A2(_06697_),
    .A3(_06778_),
    .A4(_02716_),
    .ZN(_02717_));
 NAND2_X1 _16254_ (.A1(_00052_),
    .A2(_06581_),
    .ZN(_02718_));
 OR3_X1 _16255_ (.A1(\dynamic_node_top.west_output.control.planned_f ),
    .A2(_02717_),
    .A3(_02718_),
    .ZN(_02719_));
 AOI211_X2 _16256_ (.A(_06609_),
    .B(_05185_),
    .C1(_06615_),
    .C2(_06617_),
    .ZN(_02720_));
 OAI222_X2 _16257_ (.A1(_05478_),
    .A2(_06636_),
    .B1(_06659_),
    .B2(_05470_),
    .C1(_05481_),
    .C2(_05590_),
    .ZN(_02721_));
 OR2_X1 _16258_ (.A1(_02720_),
    .A2(_02721_),
    .ZN(_02722_));
 OAI21_X1 _16259_ (.A(\dynamic_node_top.west_output.control.planned_f ),
    .B1(_06687_),
    .B2(_05484_),
    .ZN(_02723_));
 NAND4_X2 _16260_ (.A1(_06707_),
    .A2(_06636_),
    .A3(_06687_),
    .A4(_06690_),
    .ZN(_02724_));
 AOI21_X1 _16261_ (.A(_02722_),
    .B1(_02723_),
    .B2(_02724_),
    .ZN(_02725_));
 OR3_X1 _16262_ (.A1(_00052_),
    .A2(_06572_),
    .A3(_06605_),
    .ZN(_02726_));
 AOI211_X2 _16263_ (.A(_05487_),
    .B(_02722_),
    .C1(_02723_),
    .C2(_02724_),
    .ZN(_02727_));
 OAI221_X1 _16264_ (.A(_02715_),
    .B1(_02719_),
    .B2(_02725_),
    .C1(_02726_),
    .C2(_02727_),
    .ZN(_02288_));
 BUF_X2 _16265_ (.A(_10450_),
    .Z(_02728_));
 NAND2_X1 _16266_ (.A1(\dynamic_node_top.west_output.space.count_f[2] ),
    .A2(_02728_),
    .ZN(_02729_));
 BUF_X2 _16267_ (.A(_00058_),
    .Z(_02730_));
 NAND2_X1 _16268_ (.A1(_02730_),
    .A2(_02728_),
    .ZN(_02731_));
 OAI22_X1 _16269_ (.A1(_10550_),
    .A2(_02729_),
    .B1(_02731_),
    .B2(_10552_),
    .ZN(_02732_));
 BUF_X1 _16270_ (.A(_10444_),
    .Z(_02733_));
 NOR3_X1 _16271_ (.A1(_02733_),
    .A2(_10551_),
    .A3(_10549_),
    .ZN(_02734_));
 AOI21_X1 _16272_ (.A(_02734_),
    .B1(_10448_),
    .B2(_02733_),
    .ZN(_02735_));
 OAI21_X2 _16273_ (.A(_02728_),
    .B1(_02730_),
    .B2(\dynamic_node_top.west_output.space.count_f[2] ),
    .ZN(_02736_));
 AOI21_X1 _16274_ (.A(_02732_),
    .B1(_02735_),
    .B2(_02736_),
    .ZN(_02737_));
 NOR2_X1 _16275_ (.A1(_02420_),
    .A2(_02737_),
    .ZN(_02289_));
 CLKBUF_X2 _16276_ (.A(_10446_),
    .Z(_02738_));
 NAND4_X1 _16277_ (.A1(_10451_),
    .A2(_02738_),
    .A3(_02730_),
    .A4(_02728_),
    .ZN(_02739_));
 INV_X1 _16278_ (.A(_10451_),
    .ZN(_02740_));
 NAND2_X1 _16279_ (.A1(_10443_),
    .A2(_02740_),
    .ZN(_02741_));
 OAI21_X1 _16280_ (.A(_02739_),
    .B1(_02741_),
    .B2(_02729_),
    .ZN(_02742_));
 INV_X1 _16281_ (.A(_02738_),
    .ZN(_02743_));
 OAI21_X1 _16282_ (.A(_02741_),
    .B1(_02743_),
    .B2(_02740_),
    .ZN(_02744_));
 MUX2_X1 _16283_ (.A(_02744_),
    .B(\dynamic_node_top.west_output.space.count_f[1] ),
    .S(_02733_),
    .Z(_02745_));
 INV_X1 _16284_ (.A(_10449_),
    .ZN(_02746_));
 OAI22_X2 _16285_ (.A1(_10443_),
    .A2(_02729_),
    .B1(_02731_),
    .B2(_02738_),
    .ZN(_02747_));
 AOI221_X2 _16286_ (.A(_02742_),
    .B1(_02745_),
    .B2(_02736_),
    .C1(_02746_),
    .C2(_02747_),
    .ZN(_02748_));
 NOR2_X1 _16287_ (.A1(_02420_),
    .A2(_02748_),
    .ZN(_02290_));
 NAND2_X1 _16288_ (.A1(_10443_),
    .A2(_10452_),
    .ZN(_02749_));
 XOR2_X1 _16289_ (.A(_02730_),
    .B(_02749_),
    .Z(_02750_));
 MUX2_X1 _16290_ (.A(_02733_),
    .B(_02750_),
    .S(_02728_),
    .Z(_02751_));
 NAND2_X1 _16291_ (.A1(\dynamic_node_top.west_output.space.count_f[2] ),
    .A2(_02751_),
    .ZN(_02752_));
 INV_X1 _16292_ (.A(_02736_),
    .ZN(_02753_));
 XNOR2_X1 _16293_ (.A(_02730_),
    .B(_10454_),
    .ZN(_02754_));
 XNOR2_X1 _16294_ (.A(_02730_),
    .B(_10452_),
    .ZN(_02755_));
 AOI22_X1 _16295_ (.A1(_02738_),
    .A2(_02754_),
    .B1(_02755_),
    .B2(_10443_),
    .ZN(_02756_));
 OR3_X1 _16296_ (.A1(_02733_),
    .A2(_02753_),
    .A3(_02756_),
    .ZN(_02757_));
 NAND4_X1 _16297_ (.A1(_02738_),
    .A2(_02730_),
    .A3(_10454_),
    .A4(_02728_),
    .ZN(_02758_));
 AND2_X1 _16298_ (.A1(_06754_),
    .A2(_02758_),
    .ZN(_02759_));
 NAND3_X1 _16299_ (.A1(_02752_),
    .A2(_02757_),
    .A3(_02759_),
    .ZN(_02291_));
 NAND4_X1 _16300_ (.A1(_02748_),
    .A2(_02752_),
    .A3(_02757_),
    .A4(_02759_),
    .ZN(_02293_));
 NOR2_X1 _16301_ (.A1(_02737_),
    .A2(_02293_),
    .ZN(_02292_));
 AND2_X1 _16302_ (.A1(_02637_),
    .A2(net756),
    .ZN(_02294_));
 AND2_X1 _16303_ (.A1(_06755_),
    .A2(net299),
    .ZN(_02295_));
 BUF_X4 _16304_ (.A(_05163_),
    .Z(_02760_));
 BUF_X4 _16305_ (.A(_06960_),
    .Z(_02761_));
 BUF_X2 _16306_ (.A(_05468_),
    .Z(_02762_));
 BUF_X4 _16307_ (.A(_07286_),
    .Z(_02763_));
 MUX2_X1 _16308_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][0] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][0] ),
    .S(_02763_),
    .Z(_02764_));
 OR2_X1 _16309_ (.A1(_02762_),
    .A2(_02764_),
    .ZN(_02765_));
 MUX2_X1 _16310_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][0] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][0] ),
    .S(_07523_),
    .Z(_02766_));
 BUF_X8 _16311_ (.A(_07525_),
    .Z(_02767_));
 OAI21_X4 _16312_ (.A(_02765_),
    .B1(_02766_),
    .B2(_02767_),
    .ZN(_02768_));
 BUF_X8 _16313_ (.A(_07244_),
    .Z(_02769_));
 BUF_X4 _16314_ (.A(net743),
    .Z(_02770_));
 MUX2_X1 _16315_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][0] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][0] ),
    .S(_02770_),
    .Z(_02771_));
 INV_X1 _16316_ (.A(_02771_),
    .ZN(_02772_));
 NAND2_X1 _16317_ (.A1(_02769_),
    .A2(_02772_),
    .ZN(_02773_));
 BUF_X4 _16318_ (.A(net745),
    .Z(_02774_));
 MUX2_X1 _16319_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][0] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][0] ),
    .S(_02774_),
    .Z(_02775_));
 BUF_X4 _16320_ (.A(_07244_),
    .Z(_02776_));
 OAI21_X4 _16321_ (.A(_02773_),
    .B1(_02775_),
    .B2(_02776_),
    .ZN(_02777_));
 BUF_X4 _16322_ (.A(_00074_),
    .Z(_02778_));
 BUF_X4 _16323_ (.A(_02778_),
    .Z(_02779_));
 BUF_X4 _16324_ (.A(_02779_),
    .Z(_02780_));
 OAI22_X1 _16325_ (.A1(_02761_),
    .A2(_02768_),
    .B1(_02777_),
    .B2(_02780_),
    .ZN(_02781_));
 BUF_X4 _16326_ (.A(_05156_),
    .Z(_02782_));
 BUF_X4 _16327_ (.A(_02782_),
    .Z(_02783_));
 BUF_X2 _16328_ (.A(_07268_),
    .Z(_02784_));
 BUF_X4 _16329_ (.A(_07273_),
    .Z(_02785_));
 MUX2_X1 _16330_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][0] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][0] ),
    .S(_02785_),
    .Z(_02786_));
 OR2_X1 _16331_ (.A1(_02784_),
    .A2(_02786_),
    .ZN(_02787_));
 MUX2_X1 _16332_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][0] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][0] ),
    .S(_07440_),
    .Z(_02788_));
 BUF_X8 _16333_ (.A(_07445_),
    .Z(_02789_));
 OAI21_X4 _16334_ (.A(_02787_),
    .B1(_02788_),
    .B2(_02789_),
    .ZN(_02790_));
 CLKBUF_X3 _16335_ (.A(_05321_),
    .Z(_02791_));
 BUF_X4 _16336_ (.A(_05314_),
    .Z(_02792_));
 MUX2_X1 _16337_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][0] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][0] ),
    .S(_02792_),
    .Z(_02793_));
 OR2_X1 _16338_ (.A1(_02791_),
    .A2(_02793_),
    .ZN(_02794_));
 BUF_X4 _16339_ (.A(_05315_),
    .Z(_02795_));
 MUX2_X1 _16340_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][0] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][0] ),
    .S(_02795_),
    .Z(_02796_));
 BUF_X8 _16341_ (.A(_05326_),
    .Z(_02797_));
 OAI21_X4 _16342_ (.A(_02794_),
    .B1(_02796_),
    .B2(_02797_),
    .ZN(_02798_));
 BUF_X4 _16343_ (.A(_00075_),
    .Z(_02799_));
 BUF_X4 _16344_ (.A(_02799_),
    .Z(_02800_));
 BUF_X4 _16345_ (.A(_02800_),
    .Z(_02801_));
 OAI22_X1 _16346_ (.A1(_02783_),
    .A2(_02790_),
    .B1(_02798_),
    .B2(_02801_),
    .ZN(_02802_));
 BUF_X4 _16347_ (.A(_00076_),
    .Z(_02803_));
 CLKBUF_X3 _16348_ (.A(_02803_),
    .Z(_02804_));
 BUF_X8 _16349_ (.A(_05977_),
    .Z(_02805_));
 BUF_X4 _16350_ (.A(_07130_),
    .Z(_02806_));
 BUF_X8 _16351_ (.A(_05702_),
    .Z(_02807_));
 BUF_X4 _16352_ (.A(_02807_),
    .Z(_02808_));
 MUX2_X1 _16353_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][0] ),
    .S(_02808_),
    .Z(_02809_));
 BUF_X4 _16354_ (.A(_02807_),
    .Z(_02810_));
 MUX2_X1 _16355_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][0] ),
    .S(_02810_),
    .Z(_02811_));
 BUF_X4 _16356_ (.A(_05710_),
    .Z(_02812_));
 MUX2_X1 _16357_ (.A(_02809_),
    .B(_02811_),
    .S(_02812_),
    .Z(_02813_));
 NAND2_X1 _16358_ (.A1(_02806_),
    .A2(_02813_),
    .ZN(_02814_));
 BUF_X4 _16359_ (.A(_05720_),
    .Z(_02815_));
 BUF_X4 _16360_ (.A(_02807_),
    .Z(_02816_));
 MUX2_X1 _16361_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][0] ),
    .S(_02816_),
    .Z(_02817_));
 BUF_X4 _16362_ (.A(_02807_),
    .Z(_02818_));
 MUX2_X1 _16363_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][0] ),
    .S(_02818_),
    .Z(_02819_));
 BUF_X4 _16364_ (.A(_05710_),
    .Z(_02820_));
 MUX2_X1 _16365_ (.A(_02817_),
    .B(_02819_),
    .S(_02820_),
    .Z(_02821_));
 NAND2_X1 _16366_ (.A1(_02815_),
    .A2(_02821_),
    .ZN(_02822_));
 NAND3_X2 _16367_ (.A1(_02805_),
    .A2(_02814_),
    .A3(_02822_),
    .ZN(_02823_));
 BUF_X4 _16368_ (.A(_05702_),
    .Z(_02824_));
 MUX2_X1 _16369_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][0] ),
    .S(_02824_),
    .Z(_02825_));
 BUF_X4 _16370_ (.A(_05702_),
    .Z(_02826_));
 MUX2_X1 _16371_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][0] ),
    .S(_02826_),
    .Z(_02827_));
 BUF_X4 _16372_ (.A(_05709_),
    .Z(_02828_));
 MUX2_X1 _16373_ (.A(_02825_),
    .B(_02827_),
    .S(_02828_),
    .Z(_02829_));
 BUF_X4 _16374_ (.A(_05702_),
    .Z(_02830_));
 MUX2_X1 _16375_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][0] ),
    .S(_02830_),
    .Z(_02831_));
 BUF_X8 _16376_ (.A(_02807_),
    .Z(_02832_));
 MUX2_X1 _16377_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][0] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][0] ),
    .S(_02832_),
    .Z(_02833_));
 BUF_X4 _16378_ (.A(_05709_),
    .Z(_02834_));
 MUX2_X1 _16379_ (.A(_02831_),
    .B(_02833_),
    .S(_02834_),
    .Z(_02835_));
 BUF_X4 _16380_ (.A(_05720_),
    .Z(_02836_));
 MUX2_X1 _16381_ (.A(_02829_),
    .B(_02835_),
    .S(_02836_),
    .Z(_02837_));
 BUF_X4 _16382_ (.A(_05977_),
    .Z(_02838_));
 BUF_X8 _16383_ (.A(_02838_),
    .Z(_02839_));
 OAI21_X4 _16384_ (.A(_02823_),
    .B1(_02837_),
    .B2(_02839_),
    .ZN(_02840_));
 NOR2_X1 _16385_ (.A1(_02804_),
    .A2(_02840_),
    .ZN(_02841_));
 NOR3_X1 _16386_ (.A1(_02781_),
    .A2(_02802_),
    .A3(_02841_),
    .ZN(_02842_));
 NOR2_X2 _16387_ (.A1(_02760_),
    .A2(_02842_),
    .ZN(net300));
 BUF_X8 _16388_ (.A(_05163_),
    .Z(_02843_));
 BUF_X4 _16389_ (.A(_02779_),
    .Z(_02844_));
 BUF_X4 _16390_ (.A(_07244_),
    .Z(_02845_));
 MUX2_X1 _16391_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][10] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][10] ),
    .S(_07246_),
    .Z(_02846_));
 INV_X1 _16392_ (.A(_02846_),
    .ZN(_02847_));
 NAND2_X1 _16393_ (.A1(_02845_),
    .A2(_02847_),
    .ZN(_02848_));
 MUX2_X1 _16394_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][10] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][10] ),
    .S(_07250_),
    .Z(_02849_));
 OAI21_X4 _16395_ (.A(_02848_),
    .B1(_02849_),
    .B2(_07244_),
    .ZN(_02850_));
 MUX2_X1 _16396_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][10] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][10] ),
    .S(_07520_),
    .Z(_02851_));
 OR2_X1 _16397_ (.A1(_07519_),
    .A2(_02851_),
    .ZN(_02852_));
 MUX2_X1 _16398_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][10] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][10] ),
    .S(_07523_),
    .Z(_02853_));
 OAI21_X4 _16399_ (.A(_02852_),
    .B1(_02853_),
    .B2(_07526_),
    .ZN(_02854_));
 BUF_X4 _16400_ (.A(_06960_),
    .Z(_02855_));
 OAI22_X1 _16401_ (.A1(_02844_),
    .A2(_02850_),
    .B1(_02854_),
    .B2(_02855_),
    .ZN(_02856_));
 BUF_X4 _16402_ (.A(_02782_),
    .Z(_02857_));
 BUF_X2 _16403_ (.A(_07268_),
    .Z(_02858_));
 BUF_X4 _16404_ (.A(_07273_),
    .Z(_02859_));
 MUX2_X1 _16405_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][10] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][10] ),
    .S(_02859_),
    .Z(_02860_));
 OR2_X1 _16406_ (.A1(_02858_),
    .A2(_02860_),
    .ZN(_02861_));
 MUX2_X1 _16407_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][10] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][10] ),
    .S(_07443_),
    .Z(_02862_));
 BUF_X8 _16408_ (.A(_07445_),
    .Z(_02863_));
 OAI21_X4 _16409_ (.A(_02861_),
    .B1(_02862_),
    .B2(_02863_),
    .ZN(_02864_));
 MUX2_X1 _16410_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][10] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][10] ),
    .S(_07494_),
    .Z(_02865_));
 OR2_X1 _16411_ (.A1(_07493_),
    .A2(_02865_),
    .ZN(_02866_));
 MUX2_X1 _16412_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][10] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][10] ),
    .S(_07497_),
    .Z(_02867_));
 OAI21_X2 _16413_ (.A(_02866_),
    .B1(_02867_),
    .B2(_07499_),
    .ZN(_02868_));
 BUF_X4 _16414_ (.A(_02800_),
    .Z(_02869_));
 OAI22_X1 _16415_ (.A1(_02857_),
    .A2(_02864_),
    .B1(_02868_),
    .B2(_02869_),
    .ZN(_02870_));
 NOR2_X1 _16416_ (.A1(_02856_),
    .A2(_02870_),
    .ZN(_02871_));
 INV_X1 _16417_ (.A(_02803_),
    .ZN(_02872_));
 CLKBUF_X3 _16418_ (.A(_02872_),
    .Z(_02873_));
 BUF_X4 _16419_ (.A(_02873_),
    .Z(_02874_));
 BUF_X4 _16420_ (.A(_02807_),
    .Z(_02875_));
 MUX2_X1 _16421_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][10] ),
    .S(_02875_),
    .Z(_02876_));
 BUF_X4 _16422_ (.A(_02807_),
    .Z(_02877_));
 MUX2_X1 _16423_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][10] ),
    .S(_02877_),
    .Z(_02878_));
 BUF_X4 _16424_ (.A(_05710_),
    .Z(_02879_));
 MUX2_X1 _16425_ (.A(_02876_),
    .B(_02878_),
    .S(_02879_),
    .Z(_02880_));
 MUX2_X1 _16426_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][10] ),
    .S(_02877_),
    .Z(_02881_));
 BUF_X4 _16427_ (.A(_05703_),
    .Z(_02882_));
 MUX2_X1 _16428_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][10] ),
    .S(_02882_),
    .Z(_02883_));
 MUX2_X1 _16429_ (.A(_02881_),
    .B(_02883_),
    .S(_02879_),
    .Z(_02884_));
 BUF_X4 _16430_ (.A(_05720_),
    .Z(_02885_));
 MUX2_X1 _16431_ (.A(_02880_),
    .B(_02884_),
    .S(_02885_),
    .Z(_02886_));
 MUX2_X1 _16432_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][10] ),
    .S(_02882_),
    .Z(_02887_));
 BUF_X4 _16433_ (.A(_05703_),
    .Z(_02888_));
 MUX2_X1 _16434_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][10] ),
    .S(_02888_),
    .Z(_02889_));
 BUF_X4 _16435_ (.A(_05710_),
    .Z(_02890_));
 MUX2_X1 _16436_ (.A(_02887_),
    .B(_02889_),
    .S(_02890_),
    .Z(_02891_));
 MUX2_X1 _16437_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][10] ),
    .S(_02888_),
    .Z(_02892_));
 MUX2_X1 _16438_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][10] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][10] ),
    .S(_02888_),
    .Z(_02893_));
 MUX2_X1 _16439_ (.A(_02892_),
    .B(_02893_),
    .S(_05711_),
    .Z(_02894_));
 MUX2_X1 _16440_ (.A(_02891_),
    .B(_02894_),
    .S(_05721_),
    .Z(_02895_));
 MUX2_X2 _16441_ (.A(_02886_),
    .B(_02895_),
    .S(_07393_),
    .Z(_02896_));
 NAND2_X1 _16442_ (.A1(_02874_),
    .A2(_02896_),
    .ZN(_02897_));
 AOI21_X2 _16443_ (.A(_02843_),
    .B1(_02871_),
    .B2(_02897_),
    .ZN(net301));
 MUX2_X1 _16444_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][11] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][11] ),
    .S(_02763_),
    .Z(_02898_));
 OR2_X1 _16445_ (.A1(_07519_),
    .A2(_02898_),
    .ZN(_02899_));
 MUX2_X1 _16446_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][11] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][11] ),
    .S(_07523_),
    .Z(_02900_));
 OAI21_X4 _16447_ (.A(_02899_),
    .B1(_02900_),
    .B2(_07526_),
    .ZN(_02901_));
 MUX2_X1 _16448_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][11] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][11] ),
    .S(_02859_),
    .Z(_02902_));
 OR2_X1 _16449_ (.A1(_02858_),
    .A2(_02902_),
    .ZN(_02903_));
 MUX2_X1 _16450_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][11] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][11] ),
    .S(_07443_),
    .Z(_02904_));
 OAI21_X4 _16451_ (.A(_02903_),
    .B1(_02904_),
    .B2(_07446_),
    .ZN(_02905_));
 BUF_X4 _16452_ (.A(_02782_),
    .Z(_02906_));
 OAI22_X2 _16453_ (.A1(_02761_),
    .A2(_02901_),
    .B1(_02905_),
    .B2(_02906_),
    .ZN(_02907_));
 MUX2_X1 _16454_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][11] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][11] ),
    .S(_07246_),
    .Z(_02908_));
 INV_X1 _16455_ (.A(_02908_),
    .ZN(_02909_));
 NAND2_X1 _16456_ (.A1(_02845_),
    .A2(_02909_),
    .ZN(_02910_));
 MUX2_X1 _16457_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][11] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][11] ),
    .S(_07250_),
    .Z(_02911_));
 OAI21_X4 _16458_ (.A(_02910_),
    .B1(_02911_),
    .B2(_07244_),
    .ZN(_02912_));
 MUX2_X1 _16459_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][11] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][11] ),
    .S(_02792_),
    .Z(_02913_));
 OR2_X1 _16460_ (.A1(_07493_),
    .A2(_02913_),
    .ZN(_02914_));
 MUX2_X1 _16461_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][11] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][11] ),
    .S(_07497_),
    .Z(_02915_));
 OAI21_X4 _16462_ (.A(_02914_),
    .B1(_02915_),
    .B2(_07499_),
    .ZN(_02916_));
 OAI22_X2 _16463_ (.A1(_02844_),
    .A2(_02912_),
    .B1(_02916_),
    .B2(_02869_),
    .ZN(_02917_));
 NOR2_X2 _16464_ (.A1(_02907_),
    .A2(_02917_),
    .ZN(_02918_));
 MUX2_X1 _16465_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][11] ),
    .S(_02810_),
    .Z(_02919_));
 MUX2_X1 _16466_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][11] ),
    .S(_02877_),
    .Z(_02920_));
 MUX2_X1 _16467_ (.A(_02919_),
    .B(_02920_),
    .S(_02879_),
    .Z(_02921_));
 MUX2_X1 _16468_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][11] ),
    .S(_02877_),
    .Z(_02922_));
 MUX2_X1 _16469_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][11] ),
    .S(_02882_),
    .Z(_02923_));
 MUX2_X1 _16470_ (.A(_02922_),
    .B(_02923_),
    .S(_02879_),
    .Z(_02924_));
 MUX2_X1 _16471_ (.A(_02921_),
    .B(_02924_),
    .S(_02885_),
    .Z(_02925_));
 MUX2_X1 _16472_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][11] ),
    .S(_02882_),
    .Z(_02926_));
 MUX2_X1 _16473_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][11] ),
    .S(_02888_),
    .Z(_02927_));
 MUX2_X1 _16474_ (.A(_02926_),
    .B(_02927_),
    .S(_02890_),
    .Z(_02928_));
 BUF_X4 _16475_ (.A(_05703_),
    .Z(_02929_));
 MUX2_X1 _16476_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][11] ),
    .S(_02929_),
    .Z(_02930_));
 MUX2_X1 _16477_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][11] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][11] ),
    .S(_02888_),
    .Z(_02931_));
 MUX2_X1 _16478_ (.A(_02930_),
    .B(_02931_),
    .S(_05711_),
    .Z(_02932_));
 MUX2_X1 _16479_ (.A(_02928_),
    .B(_02932_),
    .S(_02885_),
    .Z(_02933_));
 MUX2_X2 _16480_ (.A(_02925_),
    .B(_02933_),
    .S(_07393_),
    .Z(_02934_));
 NAND2_X1 _16481_ (.A1(_02874_),
    .A2(_02934_),
    .ZN(_02935_));
 AOI21_X4 _16482_ (.A(_02843_),
    .B1(_02918_),
    .B2(_02935_),
    .ZN(net302));
 MUX2_X1 _16483_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][12] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][12] ),
    .S(_02763_),
    .Z(_02936_));
 OR2_X1 _16484_ (.A1(_02762_),
    .A2(_02936_),
    .ZN(_02937_));
 BUF_X4 _16485_ (.A(net721),
    .Z(_02938_));
 MUX2_X1 _16486_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][12] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][12] ),
    .S(_02938_),
    .Z(_02939_));
 OAI21_X4 _16487_ (.A(_02937_),
    .B1(_02939_),
    .B2(_02767_),
    .ZN(_02940_));
 BUF_X4 _16488_ (.A(_07244_),
    .Z(_02941_));
 MUX2_X1 _16489_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][12] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][12] ),
    .S(_02770_),
    .Z(_02942_));
 INV_X1 _16490_ (.A(_02942_),
    .ZN(_02943_));
 NAND2_X1 _16491_ (.A1(_02941_),
    .A2(_02943_),
    .ZN(_02944_));
 MUX2_X1 _16492_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][12] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][12] ),
    .S(_02774_),
    .Z(_02945_));
 OAI21_X4 _16493_ (.A(_02944_),
    .B1(_02945_),
    .B2(_02769_),
    .ZN(_02946_));
 OAI22_X1 _16494_ (.A1(_02761_),
    .A2(_02940_),
    .B1(_02946_),
    .B2(_02780_),
    .ZN(_02947_));
 MUX2_X1 _16495_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][12] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][12] ),
    .S(_02785_),
    .Z(_02948_));
 OR2_X1 _16496_ (.A1(_02784_),
    .A2(_02948_),
    .ZN(_02949_));
 BUF_X4 _16497_ (.A(_05147_),
    .Z(_02950_));
 MUX2_X1 _16498_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][12] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][12] ),
    .S(_02950_),
    .Z(_02951_));
 OAI21_X4 _16499_ (.A(_02949_),
    .B1(_02951_),
    .B2(_02789_),
    .ZN(_02952_));
 MUX2_X1 _16500_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][12] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][12] ),
    .S(_02792_),
    .Z(_02953_));
 OR2_X1 _16501_ (.A1(_02791_),
    .A2(_02953_),
    .ZN(_02954_));
 MUX2_X1 _16502_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][12] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][12] ),
    .S(_02795_),
    .Z(_02955_));
 OAI21_X4 _16503_ (.A(_02954_),
    .B1(_02955_),
    .B2(_02797_),
    .ZN(_02956_));
 OAI22_X1 _16504_ (.A1(_02783_),
    .A2(_02952_),
    .B1(_02956_),
    .B2(_02801_),
    .ZN(_02957_));
 MUX2_X1 _16505_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][12] ),
    .S(_02808_),
    .Z(_02958_));
 MUX2_X1 _16506_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][12] ),
    .S(_02810_),
    .Z(_02959_));
 MUX2_X1 _16507_ (.A(_02958_),
    .B(_02959_),
    .S(_02812_),
    .Z(_02960_));
 NAND2_X1 _16508_ (.A1(_02806_),
    .A2(_02960_),
    .ZN(_02961_));
 MUX2_X1 _16509_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][12] ),
    .S(_02816_),
    .Z(_02962_));
 MUX2_X1 _16510_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][12] ),
    .S(_02818_),
    .Z(_02963_));
 MUX2_X1 _16511_ (.A(_02962_),
    .B(_02963_),
    .S(_02820_),
    .Z(_02964_));
 NAND2_X1 _16512_ (.A1(_02815_),
    .A2(_02964_),
    .ZN(_02965_));
 NAND3_X2 _16513_ (.A1(_02805_),
    .A2(_02961_),
    .A3(_02965_),
    .ZN(_02966_));
 MUX2_X1 _16514_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][12] ),
    .S(_02824_),
    .Z(_02967_));
 MUX2_X1 _16515_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][12] ),
    .S(_02826_),
    .Z(_02968_));
 MUX2_X1 _16516_ (.A(_02967_),
    .B(_02968_),
    .S(_02828_),
    .Z(_02969_));
 MUX2_X1 _16517_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][12] ),
    .S(_02830_),
    .Z(_02970_));
 MUX2_X1 _16518_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][12] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][12] ),
    .S(_02832_),
    .Z(_02971_));
 MUX2_X1 _16519_ (.A(_02970_),
    .B(_02971_),
    .S(_02834_),
    .Z(_02972_));
 MUX2_X1 _16520_ (.A(_02969_),
    .B(_02972_),
    .S(_02836_),
    .Z(_02973_));
 OAI21_X4 _16521_ (.A(_02966_),
    .B1(_02973_),
    .B2(_02839_),
    .ZN(_02974_));
 NOR2_X1 _16522_ (.A1(_02804_),
    .A2(_02974_),
    .ZN(_02975_));
 NOR3_X1 _16523_ (.A1(_02947_),
    .A2(_02957_),
    .A3(_02975_),
    .ZN(_02976_));
 NOR2_X2 _16524_ (.A1(_02760_),
    .A2(_02976_),
    .ZN(net303));
 MUX2_X1 _16525_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][13] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][13] ),
    .S(_02770_),
    .Z(_02977_));
 INV_X1 _16526_ (.A(_02977_),
    .ZN(_02978_));
 NAND2_X1 _16527_ (.A1(_02845_),
    .A2(_02978_),
    .ZN(_02979_));
 MUX2_X1 _16528_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][13] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][13] ),
    .S(_07250_),
    .Z(_02980_));
 OAI21_X4 _16529_ (.A(_02979_),
    .B1(_02980_),
    .B2(_07244_),
    .ZN(_02981_));
 MUX2_X1 _16530_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][13] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][13] ),
    .S(_07520_),
    .Z(_02982_));
 OR2_X1 _16531_ (.A1(_07519_),
    .A2(_02982_),
    .ZN(_02983_));
 MUX2_X1 _16532_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][13] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][13] ),
    .S(_07523_),
    .Z(_02984_));
 OAI21_X4 _16533_ (.A(_02983_),
    .B1(_02984_),
    .B2(_07526_),
    .ZN(_02985_));
 OAI22_X1 _16534_ (.A1(_02844_),
    .A2(_02981_),
    .B1(_02985_),
    .B2(_02855_),
    .ZN(_02986_));
 MUX2_X1 _16535_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][13] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][13] ),
    .S(_02859_),
    .Z(_02987_));
 OR2_X1 _16536_ (.A1(_02858_),
    .A2(_02987_),
    .ZN(_02988_));
 MUX2_X1 _16537_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][13] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][13] ),
    .S(_07443_),
    .Z(_02989_));
 OAI21_X4 _16538_ (.A(_02988_),
    .B1(_02989_),
    .B2(_02863_),
    .ZN(_02990_));
 CLKBUF_X3 _16539_ (.A(_05321_),
    .Z(_02991_));
 MUX2_X1 _16540_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][13] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][13] ),
    .S(_02792_),
    .Z(_02992_));
 OR2_X1 _16541_ (.A1(_02991_),
    .A2(_02992_),
    .ZN(_02993_));
 MUX2_X1 _16542_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][13] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][13] ),
    .S(_07497_),
    .Z(_02994_));
 BUF_X8 _16543_ (.A(_07499_),
    .Z(_02995_));
 OAI21_X2 _16544_ (.A(_02993_),
    .B1(_02994_),
    .B2(_02995_),
    .ZN(_02996_));
 OAI22_X1 _16545_ (.A1(_02857_),
    .A2(_02990_),
    .B1(_02996_),
    .B2(_02869_),
    .ZN(_02997_));
 NOR2_X1 _16546_ (.A1(_02986_),
    .A2(_02997_),
    .ZN(_02998_));
 MUX2_X1 _16547_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][13] ),
    .S(_02810_),
    .Z(_02999_));
 MUX2_X1 _16548_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][13] ),
    .S(_02877_),
    .Z(_03000_));
 MUX2_X1 _16549_ (.A(_02999_),
    .B(_03000_),
    .S(_02879_),
    .Z(_03001_));
 MUX2_X1 _16550_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][13] ),
    .S(_02875_),
    .Z(_03002_));
 MUX2_X1 _16551_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][13] ),
    .S(_02882_),
    .Z(_03003_));
 MUX2_X1 _16552_ (.A(_03002_),
    .B(_03003_),
    .S(_02879_),
    .Z(_03004_));
 MUX2_X1 _16553_ (.A(_03001_),
    .B(_03004_),
    .S(_02885_),
    .Z(_03005_));
 MUX2_X1 _16554_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][13] ),
    .S(_02877_),
    .Z(_03006_));
 MUX2_X1 _16555_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][13] ),
    .S(_02929_),
    .Z(_03007_));
 MUX2_X1 _16556_ (.A(_03006_),
    .B(_03007_),
    .S(_02890_),
    .Z(_03008_));
 MUX2_X1 _16557_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][13] ),
    .S(_02929_),
    .Z(_03009_));
 MUX2_X1 _16558_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][13] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][13] ),
    .S(_02888_),
    .Z(_03010_));
 MUX2_X1 _16559_ (.A(_03009_),
    .B(_03010_),
    .S(_05711_),
    .Z(_03011_));
 MUX2_X1 _16560_ (.A(_03008_),
    .B(_03011_),
    .S(_02885_),
    .Z(_03012_));
 MUX2_X2 _16561_ (.A(_03005_),
    .B(_03012_),
    .S(_07393_),
    .Z(_03013_));
 NAND2_X1 _16562_ (.A1(_02874_),
    .A2(_03013_),
    .ZN(_03014_));
 AOI21_X2 _16563_ (.A(_02843_),
    .B1(_02998_),
    .B2(_03014_),
    .ZN(net304));
 CLKBUF_X3 _16564_ (.A(_06960_),
    .Z(_03015_));
 MUX2_X1 _16565_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][14] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][14] ),
    .S(_02763_),
    .Z(_03016_));
 OR2_X1 _16566_ (.A1(_02762_),
    .A2(_03016_),
    .ZN(_03017_));
 MUX2_X1 _16567_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][14] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][14] ),
    .S(_02938_),
    .Z(_03018_));
 OAI21_X4 _16568_ (.A(_03017_),
    .B1(_03018_),
    .B2(_02767_),
    .ZN(_03019_));
 MUX2_X1 _16569_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][14] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][14] ),
    .S(_02770_),
    .Z(_03020_));
 INV_X1 _16570_ (.A(_03020_),
    .ZN(_03021_));
 NAND2_X1 _16571_ (.A1(_02769_),
    .A2(_03021_),
    .ZN(_03022_));
 MUX2_X1 _16572_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][14] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][14] ),
    .S(_02774_),
    .Z(_03023_));
 OAI21_X4 _16573_ (.A(_03022_),
    .B1(_03023_),
    .B2(_02776_),
    .ZN(_03024_));
 BUF_X4 _16574_ (.A(_02778_),
    .Z(_03025_));
 OAI22_X1 _16575_ (.A1(_03015_),
    .A2(_03019_),
    .B1(_03024_),
    .B2(_03025_),
    .ZN(_03026_));
 MUX2_X1 _16576_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][14] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][14] ),
    .S(_02785_),
    .Z(_03027_));
 OR2_X1 _16577_ (.A1(_02784_),
    .A2(_03027_),
    .ZN(_03028_));
 MUX2_X1 _16578_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][14] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][14] ),
    .S(_07440_),
    .Z(_03029_));
 OAI21_X4 _16579_ (.A(_03028_),
    .B1(_03029_),
    .B2(_02789_),
    .ZN(_03030_));
 MUX2_X1 _16580_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][14] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][14] ),
    .S(_02792_),
    .Z(_03031_));
 OR2_X1 _16581_ (.A1(_02791_),
    .A2(_03031_),
    .ZN(_03032_));
 MUX2_X1 _16582_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][14] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][14] ),
    .S(_02795_),
    .Z(_03033_));
 OAI21_X4 _16583_ (.A(_03032_),
    .B1(_03033_),
    .B2(_02797_),
    .ZN(_03034_));
 OAI22_X1 _16584_ (.A1(_02783_),
    .A2(_03030_),
    .B1(_03034_),
    .B2(_02801_),
    .ZN(_03035_));
 BUF_X4 _16585_ (.A(_05977_),
    .Z(_03036_));
 MUX2_X1 _16586_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][14] ),
    .S(_02808_),
    .Z(_03037_));
 MUX2_X1 _16587_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][14] ),
    .S(_02810_),
    .Z(_03038_));
 MUX2_X1 _16588_ (.A(_03037_),
    .B(_03038_),
    .S(_02812_),
    .Z(_03039_));
 NAND2_X1 _16589_ (.A1(_02806_),
    .A2(_03039_),
    .ZN(_03040_));
 MUX2_X1 _16590_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][14] ),
    .S(_02816_),
    .Z(_03041_));
 BUF_X4 _16591_ (.A(_02807_),
    .Z(_03042_));
 MUX2_X1 _16592_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][14] ),
    .S(_03042_),
    .Z(_03043_));
 MUX2_X1 _16593_ (.A(_03041_),
    .B(_03043_),
    .S(_02820_),
    .Z(_03044_));
 NAND2_X1 _16594_ (.A1(_02815_),
    .A2(_03044_),
    .ZN(_03045_));
 NAND3_X2 _16595_ (.A1(_03036_),
    .A2(_03040_),
    .A3(_03045_),
    .ZN(_03046_));
 BUF_X4 _16596_ (.A(_05702_),
    .Z(_03047_));
 MUX2_X1 _16597_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][14] ),
    .S(_03047_),
    .Z(_03048_));
 MUX2_X1 _16598_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][14] ),
    .S(_02826_),
    .Z(_03049_));
 MUX2_X1 _16599_ (.A(_03048_),
    .B(_03049_),
    .S(_02828_),
    .Z(_03050_));
 MUX2_X1 _16600_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][14] ),
    .S(_02830_),
    .Z(_03051_));
 MUX2_X1 _16601_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][14] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][14] ),
    .S(_02832_),
    .Z(_03052_));
 MUX2_X1 _16602_ (.A(_03051_),
    .B(_03052_),
    .S(_02834_),
    .Z(_03053_));
 MUX2_X1 _16603_ (.A(_03050_),
    .B(_03053_),
    .S(_02836_),
    .Z(_03054_));
 OAI21_X4 _16604_ (.A(_03046_),
    .B1(_03054_),
    .B2(_02839_),
    .ZN(_03055_));
 NOR2_X1 _16605_ (.A1(_02804_),
    .A2(_03055_),
    .ZN(_03056_));
 NOR3_X1 _16606_ (.A1(_03026_),
    .A2(_03035_),
    .A3(_03056_),
    .ZN(_03057_));
 NOR2_X2 _16607_ (.A1(_02760_),
    .A2(_03057_),
    .ZN(net305));
 MUX2_X1 _16608_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][15] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][15] ),
    .S(_02763_),
    .Z(_03058_));
 OR2_X1 _16609_ (.A1(_02762_),
    .A2(_03058_),
    .ZN(_03059_));
 MUX2_X1 _16610_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][15] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][15] ),
    .S(_02938_),
    .Z(_03060_));
 OAI21_X4 _16611_ (.A(_03059_),
    .B1(_03060_),
    .B2(_02767_),
    .ZN(_03061_));
 MUX2_X1 _16612_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][15] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][15] ),
    .S(_02859_),
    .Z(_03062_));
 OR2_X1 _16613_ (.A1(_02858_),
    .A2(_03062_),
    .ZN(_03063_));
 MUX2_X1 _16614_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][15] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][15] ),
    .S(_02950_),
    .Z(_03064_));
 OAI21_X4 _16615_ (.A(_03063_),
    .B1(_03064_),
    .B2(_02863_),
    .ZN(_03065_));
 BUF_X4 _16616_ (.A(_02782_),
    .Z(_03066_));
 OAI22_X1 _16617_ (.A1(_03015_),
    .A2(_03061_),
    .B1(_03065_),
    .B2(_03066_),
    .ZN(_03067_));
 BUF_X4 _16618_ (.A(net743),
    .Z(_03068_));
 MUX2_X1 _16619_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][15] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][15] ),
    .S(_03068_),
    .Z(_03069_));
 INV_X1 _16620_ (.A(_03069_),
    .ZN(_03070_));
 NAND2_X1 _16621_ (.A1(_02941_),
    .A2(_03070_),
    .ZN(_03071_));
 MUX2_X1 _16622_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][15] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][15] ),
    .S(_07246_),
    .Z(_03072_));
 OAI21_X4 _16623_ (.A(_03071_),
    .B1(_03072_),
    .B2(_02769_),
    .ZN(_03073_));
 MUX2_X1 _16624_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][15] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][15] ),
    .S(_02792_),
    .Z(_03074_));
 OR2_X1 _16625_ (.A1(_02791_),
    .A2(_03074_),
    .ZN(_03075_));
 MUX2_X1 _16626_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][15] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][15] ),
    .S(_02795_),
    .Z(_03076_));
 OAI21_X4 _16627_ (.A(_03075_),
    .B1(_03076_),
    .B2(_02797_),
    .ZN(_03077_));
 OAI22_X1 _16628_ (.A1(_02780_),
    .A2(_03073_),
    .B1(_03077_),
    .B2(_02801_),
    .ZN(_03078_));
 MUX2_X1 _16629_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][15] ),
    .S(_02808_),
    .Z(_03079_));
 MUX2_X1 _16630_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][15] ),
    .S(_02810_),
    .Z(_03080_));
 MUX2_X1 _16631_ (.A(_03079_),
    .B(_03080_),
    .S(_02812_),
    .Z(_03081_));
 NAND2_X1 _16632_ (.A1(_02806_),
    .A2(_03081_),
    .ZN(_03082_));
 MUX2_X1 _16633_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][15] ),
    .S(_02816_),
    .Z(_03083_));
 MUX2_X1 _16634_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][15] ),
    .S(_03042_),
    .Z(_03084_));
 MUX2_X1 _16635_ (.A(_03083_),
    .B(_03084_),
    .S(_02820_),
    .Z(_03085_));
 NAND2_X1 _16636_ (.A1(_02815_),
    .A2(_03085_),
    .ZN(_03086_));
 NAND3_X2 _16637_ (.A1(_03036_),
    .A2(_03082_),
    .A3(_03086_),
    .ZN(_03087_));
 MUX2_X1 _16638_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][15] ),
    .S(_03047_),
    .Z(_03088_));
 MUX2_X1 _16639_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][15] ),
    .S(_02826_),
    .Z(_03089_));
 MUX2_X1 _16640_ (.A(_03088_),
    .B(_03089_),
    .S(_02828_),
    .Z(_03090_));
 MUX2_X1 _16641_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][15] ),
    .S(_02830_),
    .Z(_03091_));
 MUX2_X1 _16642_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][15] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][15] ),
    .S(_02832_),
    .Z(_03092_));
 MUX2_X1 _16643_ (.A(_03091_),
    .B(_03092_),
    .S(_02834_),
    .Z(_03093_));
 MUX2_X1 _16644_ (.A(_03090_),
    .B(_03093_),
    .S(_02836_),
    .Z(_03094_));
 OAI21_X4 _16645_ (.A(_03087_),
    .B1(_03094_),
    .B2(_02839_),
    .ZN(_03095_));
 NOR2_X1 _16646_ (.A1(_02804_),
    .A2(_03095_),
    .ZN(_03096_));
 NOR3_X1 _16647_ (.A1(_03067_),
    .A2(_03078_),
    .A3(_03096_),
    .ZN(_03097_));
 NOR2_X1 _16648_ (.A1(_02760_),
    .A2(_03097_),
    .ZN(net306));
 MUX2_X1 _16649_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][16] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][16] ),
    .S(_02770_),
    .Z(_03098_));
 INV_X1 _16650_ (.A(_03098_),
    .ZN(_03099_));
 NAND2_X1 _16651_ (.A1(_02845_),
    .A2(_03099_),
    .ZN(_03100_));
 MUX2_X1 _16652_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][16] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][16] ),
    .S(_07250_),
    .Z(_03101_));
 OAI21_X4 _16653_ (.A(_03100_),
    .B1(_03101_),
    .B2(_07244_),
    .ZN(_03102_));
 MUX2_X1 _16654_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][16] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][16] ),
    .S(_02859_),
    .Z(_03103_));
 OR2_X1 _16655_ (.A1(_02858_),
    .A2(_03103_),
    .ZN(_03104_));
 MUX2_X1 _16656_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][16] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][16] ),
    .S(_07443_),
    .Z(_03105_));
 OAI21_X4 _16657_ (.A(_03104_),
    .B1(_03105_),
    .B2(_07446_),
    .ZN(_03106_));
 OAI22_X1 _16658_ (.A1(_02844_),
    .A2(_03102_),
    .B1(_03106_),
    .B2(_02906_),
    .ZN(_03107_));
 MUX2_X1 _16659_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][16] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][16] ),
    .S(_07520_),
    .Z(_03108_));
 OR2_X1 _16660_ (.A1(_07519_),
    .A2(_03108_),
    .ZN(_03109_));
 MUX2_X1 _16661_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][16] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][16] ),
    .S(_07523_),
    .Z(_03110_));
 OAI21_X4 _16662_ (.A(_03109_),
    .B1(_03110_),
    .B2(_07526_),
    .ZN(_03111_));
 MUX2_X1 _16663_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][16] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][16] ),
    .S(_02792_),
    .Z(_03112_));
 OR2_X1 _16664_ (.A1(_02991_),
    .A2(_03112_),
    .ZN(_03113_));
 MUX2_X1 _16665_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][16] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][16] ),
    .S(_07497_),
    .Z(_03114_));
 OAI21_X2 _16666_ (.A(_03113_),
    .B1(_03114_),
    .B2(_02995_),
    .ZN(_03115_));
 OAI22_X1 _16667_ (.A1(_02761_),
    .A2(_03111_),
    .B1(_03115_),
    .B2(_02869_),
    .ZN(_03116_));
 NOR2_X1 _16668_ (.A1(_03107_),
    .A2(_03116_),
    .ZN(_03117_));
 MUX2_X1 _16669_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][16] ),
    .S(_02810_),
    .Z(_03118_));
 MUX2_X1 _16670_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][16] ),
    .S(_02875_),
    .Z(_03119_));
 MUX2_X1 _16671_ (.A(_03118_),
    .B(_03119_),
    .S(_02812_),
    .Z(_03120_));
 MUX2_X1 _16672_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][16] ),
    .S(_02875_),
    .Z(_03121_));
 MUX2_X1 _16673_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][16] ),
    .S(_02882_),
    .Z(_03122_));
 MUX2_X1 _16674_ (.A(_03121_),
    .B(_03122_),
    .S(_02879_),
    .Z(_03123_));
 MUX2_X1 _16675_ (.A(_03120_),
    .B(_03123_),
    .S(_02885_),
    .Z(_03124_));
 MUX2_X1 _16676_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][16] ),
    .S(_02877_),
    .Z(_03125_));
 MUX2_X1 _16677_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][16] ),
    .S(_02929_),
    .Z(_03126_));
 MUX2_X1 _16678_ (.A(_03125_),
    .B(_03126_),
    .S(_02890_),
    .Z(_03127_));
 MUX2_X1 _16679_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][16] ),
    .S(_02929_),
    .Z(_03128_));
 MUX2_X1 _16680_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][16] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][16] ),
    .S(_02888_),
    .Z(_03129_));
 MUX2_X1 _16681_ (.A(_03128_),
    .B(_03129_),
    .S(_05711_),
    .Z(_03130_));
 MUX2_X1 _16682_ (.A(_03127_),
    .B(_03130_),
    .S(_02885_),
    .Z(_03131_));
 MUX2_X2 _16683_ (.A(_03124_),
    .B(_03131_),
    .S(_07393_),
    .Z(_03132_));
 NAND2_X1 _16684_ (.A1(_02874_),
    .A2(_03132_),
    .ZN(_03133_));
 AOI21_X2 _16685_ (.A(_02843_),
    .B1(_03117_),
    .B2(_03133_),
    .ZN(net307));
 MUX2_X1 _16686_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][17] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][17] ),
    .S(_02763_),
    .Z(_03134_));
 OR2_X1 _16687_ (.A1(_02762_),
    .A2(_03134_),
    .ZN(_03135_));
 MUX2_X1 _16688_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][17] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][17] ),
    .S(_07523_),
    .Z(_03136_));
 OAI21_X4 _16689_ (.A(_03135_),
    .B1(_03136_),
    .B2(_02767_),
    .ZN(_03137_));
 MUX2_X1 _16690_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][17] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][17] ),
    .S(_07440_),
    .Z(_03138_));
 OR2_X1 _16691_ (.A1(_07439_),
    .A2(_03138_),
    .ZN(_03139_));
 MUX2_X1 _16692_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][17] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][17] ),
    .S(_07443_),
    .Z(_03140_));
 OAI21_X4 _16693_ (.A(_03139_),
    .B1(_03140_),
    .B2(_07446_),
    .ZN(_03141_));
 OAI22_X2 _16694_ (.A1(_02761_),
    .A2(_03137_),
    .B1(_03141_),
    .B2(_02906_),
    .ZN(_03142_));
 MUX2_X1 _16695_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][17] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][17] ),
    .S(_07246_),
    .Z(_03143_));
 INV_X1 _16696_ (.A(_03143_),
    .ZN(_03144_));
 NAND2_X1 _16697_ (.A1(_02845_),
    .A2(_03144_),
    .ZN(_03145_));
 MUX2_X1 _16698_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][17] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][17] ),
    .S(_07250_),
    .Z(_03146_));
 OAI21_X4 _16699_ (.A(_03145_),
    .B1(_03146_),
    .B2(_07244_),
    .ZN(_03147_));
 MUX2_X1 _16700_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][17] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][17] ),
    .S(_02792_),
    .Z(_03148_));
 OR2_X1 _16701_ (.A1(_02991_),
    .A2(_03148_),
    .ZN(_03149_));
 MUX2_X1 _16702_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][17] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][17] ),
    .S(_07497_),
    .Z(_03150_));
 OAI21_X4 _16703_ (.A(_03149_),
    .B1(_03150_),
    .B2(_02995_),
    .ZN(_03151_));
 OAI22_X2 _16704_ (.A1(_02844_),
    .A2(_03147_),
    .B1(_03151_),
    .B2(_02869_),
    .ZN(_03152_));
 NOR2_X2 _16705_ (.A1(_03142_),
    .A2(_03152_),
    .ZN(_03153_));
 MUX2_X1 _16706_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][17] ),
    .S(_02810_),
    .Z(_03154_));
 MUX2_X1 _16707_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][17] ),
    .S(_02875_),
    .Z(_03155_));
 MUX2_X1 _16708_ (.A(_03154_),
    .B(_03155_),
    .S(_02812_),
    .Z(_03156_));
 MUX2_X1 _16709_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][17] ),
    .S(_02875_),
    .Z(_03157_));
 MUX2_X1 _16710_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][17] ),
    .S(_02882_),
    .Z(_03158_));
 MUX2_X1 _16711_ (.A(_03157_),
    .B(_03158_),
    .S(_02879_),
    .Z(_03159_));
 MUX2_X1 _16712_ (.A(_03156_),
    .B(_03159_),
    .S(_02836_),
    .Z(_03160_));
 MUX2_X1 _16713_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][17] ),
    .S(_02877_),
    .Z(_03161_));
 MUX2_X1 _16714_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][17] ),
    .S(_02929_),
    .Z(_03162_));
 MUX2_X1 _16715_ (.A(_03161_),
    .B(_03162_),
    .S(_02890_),
    .Z(_03163_));
 MUX2_X1 _16716_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][17] ),
    .S(_02929_),
    .Z(_03164_));
 MUX2_X1 _16717_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][17] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][17] ),
    .S(_02888_),
    .Z(_03165_));
 MUX2_X1 _16718_ (.A(_03164_),
    .B(_03165_),
    .S(_02890_),
    .Z(_03166_));
 MUX2_X1 _16719_ (.A(_03163_),
    .B(_03166_),
    .S(_02885_),
    .Z(_03167_));
 MUX2_X2 _16720_ (.A(_03160_),
    .B(_03167_),
    .S(_07393_),
    .Z(_03168_));
 NAND2_X1 _16721_ (.A1(_02874_),
    .A2(_03168_),
    .ZN(_03169_));
 AOI21_X4 _16722_ (.A(_02843_),
    .B1(_03153_),
    .B2(_03169_),
    .ZN(net308));
 MUX2_X1 _16723_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][18] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][18] ),
    .S(_02763_),
    .Z(_03170_));
 OR2_X1 _16724_ (.A1(_02762_),
    .A2(_03170_),
    .ZN(_03171_));
 MUX2_X1 _16725_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][18] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][18] ),
    .S(_02938_),
    .Z(_03172_));
 OAI21_X4 _16726_ (.A(_03171_),
    .B1(_03172_),
    .B2(_02767_),
    .ZN(_03173_));
 MUX2_X1 _16727_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][18] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][18] ),
    .S(_03068_),
    .Z(_03174_));
 INV_X1 _16728_ (.A(_03174_),
    .ZN(_03175_));
 NAND2_X1 _16729_ (.A1(_02941_),
    .A2(_03175_),
    .ZN(_03176_));
 MUX2_X1 _16730_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][18] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][18] ),
    .S(_02774_),
    .Z(_03177_));
 OAI21_X4 _16731_ (.A(_03176_),
    .B1(_03177_),
    .B2(_02769_),
    .ZN(_03178_));
 OAI22_X1 _16732_ (.A1(_03015_),
    .A2(_03173_),
    .B1(_03178_),
    .B2(_03025_),
    .ZN(_03179_));
 MUX2_X1 _16733_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][18] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][18] ),
    .S(_02785_),
    .Z(_03180_));
 OR2_X1 _16734_ (.A1(_02784_),
    .A2(_03180_),
    .ZN(_03181_));
 MUX2_X1 _16735_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][18] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][18] ),
    .S(_02950_),
    .Z(_03182_));
 OAI21_X4 _16736_ (.A(_03181_),
    .B1(_03182_),
    .B2(_02789_),
    .ZN(_03183_));
 BUF_X4 _16737_ (.A(_05314_),
    .Z(_03184_));
 MUX2_X1 _16738_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][18] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][18] ),
    .S(_03184_),
    .Z(_03185_));
 OR2_X1 _16739_ (.A1(_02791_),
    .A2(_03185_),
    .ZN(_03186_));
 MUX2_X1 _16740_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][18] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][18] ),
    .S(_02795_),
    .Z(_03187_));
 OAI21_X4 _16741_ (.A(_03186_),
    .B1(_03187_),
    .B2(_02797_),
    .ZN(_03188_));
 OAI22_X1 _16742_ (.A1(_02783_),
    .A2(_03183_),
    .B1(_03188_),
    .B2(_02801_),
    .ZN(_03189_));
 MUX2_X1 _16743_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][18] ),
    .S(_02808_),
    .Z(_03190_));
 BUF_X4 _16744_ (.A(_02807_),
    .Z(_03191_));
 MUX2_X1 _16745_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][18] ),
    .S(_03191_),
    .Z(_03192_));
 MUX2_X1 _16746_ (.A(_03190_),
    .B(_03192_),
    .S(_02812_),
    .Z(_03193_));
 NAND2_X1 _16747_ (.A1(_02806_),
    .A2(_03193_),
    .ZN(_03194_));
 MUX2_X1 _16748_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][18] ),
    .S(_02816_),
    .Z(_03195_));
 MUX2_X1 _16749_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][18] ),
    .S(_03042_),
    .Z(_03196_));
 MUX2_X1 _16750_ (.A(_03195_),
    .B(_03196_),
    .S(_02820_),
    .Z(_03197_));
 NAND2_X1 _16751_ (.A1(_02815_),
    .A2(_03197_),
    .ZN(_03198_));
 NAND3_X2 _16752_ (.A1(_03036_),
    .A2(_03194_),
    .A3(_03198_),
    .ZN(_03199_));
 MUX2_X1 _16753_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][18] ),
    .S(_03047_),
    .Z(_03200_));
 MUX2_X1 _16754_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][18] ),
    .S(_02826_),
    .Z(_03201_));
 MUX2_X1 _16755_ (.A(_03200_),
    .B(_03201_),
    .S(_02828_),
    .Z(_03202_));
 BUF_X4 _16756_ (.A(_05702_),
    .Z(_03203_));
 MUX2_X1 _16757_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][18] ),
    .S(_03203_),
    .Z(_03204_));
 MUX2_X1 _16758_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][18] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][18] ),
    .S(_02832_),
    .Z(_03205_));
 BUF_X4 _16759_ (.A(_05709_),
    .Z(_03206_));
 MUX2_X1 _16760_ (.A(_03204_),
    .B(_03205_),
    .S(_03206_),
    .Z(_03207_));
 MUX2_X1 _16761_ (.A(_03202_),
    .B(_03207_),
    .S(_02836_),
    .Z(_03208_));
 OAI21_X4 _16762_ (.A(_03199_),
    .B1(_03208_),
    .B2(_02839_),
    .ZN(_03209_));
 NOR2_X1 _16763_ (.A1(_02804_),
    .A2(_03209_),
    .ZN(_03210_));
 NOR3_X1 _16764_ (.A1(_03179_),
    .A2(_03189_),
    .A3(_03210_),
    .ZN(_03211_));
 NOR2_X1 _16765_ (.A1(_02760_),
    .A2(_03211_),
    .ZN(net309));
 BUF_X4 _16766_ (.A(_02800_),
    .Z(_03212_));
 MUX2_X1 _16767_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][19] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][19] ),
    .S(_07494_),
    .Z(_03213_));
 OR2_X1 _16768_ (.A1(_07493_),
    .A2(_03213_),
    .ZN(_03214_));
 MUX2_X1 _16769_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][19] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][19] ),
    .S(_07497_),
    .Z(_03215_));
 OAI21_X4 _16770_ (.A(_03214_),
    .B1(_03215_),
    .B2(_07499_),
    .ZN(_03216_));
 MUX2_X1 _16771_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][19] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][19] ),
    .S(_02859_),
    .Z(_03217_));
 OR2_X1 _16772_ (.A1(_02858_),
    .A2(_03217_),
    .ZN(_03218_));
 MUX2_X1 _16773_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][19] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][19] ),
    .S(_07443_),
    .Z(_03219_));
 OAI21_X4 _16774_ (.A(_03218_),
    .B1(_03219_),
    .B2(_02863_),
    .ZN(_03220_));
 OAI22_X2 _16775_ (.A1(_03212_),
    .A2(_03216_),
    .B1(_03220_),
    .B2(_02782_),
    .ZN(_03221_));
 BUF_X2 _16776_ (.A(_05468_),
    .Z(_03222_));
 BUF_X4 _16777_ (.A(_07286_),
    .Z(_03223_));
 MUX2_X1 _16778_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][19] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][19] ),
    .S(_03223_),
    .Z(_03224_));
 OR2_X1 _16779_ (.A1(_03222_),
    .A2(_03224_),
    .ZN(_03225_));
 MUX2_X1 _16780_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][19] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][19] ),
    .S(_07520_),
    .Z(_03226_));
 BUF_X8 _16781_ (.A(_07290_),
    .Z(_03227_));
 OAI21_X4 _16782_ (.A(_03225_),
    .B1(_03226_),
    .B2(_03227_),
    .ZN(_03228_));
 MUX2_X1 _16783_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][19] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][19] ),
    .S(_03068_),
    .Z(_03229_));
 INV_X1 _16784_ (.A(_03229_),
    .ZN(_03230_));
 NAND2_X1 _16785_ (.A1(_07244_),
    .A2(_03230_),
    .ZN(_03231_));
 MUX2_X1 _16786_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][19] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][19] ),
    .S(_07246_),
    .Z(_03232_));
 BUF_X8 _16787_ (.A(_05127_),
    .Z(_03233_));
 OAI21_X4 _16788_ (.A(_03231_),
    .B1(_03232_),
    .B2(_03233_),
    .ZN(_03234_));
 BUF_X4 _16789_ (.A(_02778_),
    .Z(_03235_));
 OAI22_X2 _16790_ (.A1(_02855_),
    .A2(_03228_),
    .B1(_03234_),
    .B2(_03235_),
    .ZN(_03236_));
 MUX2_X1 _16791_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][19] ),
    .S(_02808_),
    .Z(_03237_));
 MUX2_X1 _16792_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][19] ),
    .S(_03191_),
    .Z(_03238_));
 MUX2_X1 _16793_ (.A(_03237_),
    .B(_03238_),
    .S(_02812_),
    .Z(_03239_));
 NAND2_X1 _16794_ (.A1(_02806_),
    .A2(_03239_),
    .ZN(_03240_));
 MUX2_X1 _16795_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][19] ),
    .S(_02816_),
    .Z(_03241_));
 MUX2_X1 _16796_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][19] ),
    .S(_03042_),
    .Z(_03242_));
 MUX2_X1 _16797_ (.A(_03241_),
    .B(_03242_),
    .S(_02820_),
    .Z(_03243_));
 NAND2_X1 _16798_ (.A1(_02815_),
    .A2(_03243_),
    .ZN(_03244_));
 NAND3_X2 _16799_ (.A1(_03036_),
    .A2(_03240_),
    .A3(_03244_),
    .ZN(_03245_));
 MUX2_X1 _16800_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][19] ),
    .S(_03047_),
    .Z(_03246_));
 MUX2_X1 _16801_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][19] ),
    .S(_02826_),
    .Z(_03247_));
 MUX2_X1 _16802_ (.A(_03246_),
    .B(_03247_),
    .S(_02828_),
    .Z(_03248_));
 MUX2_X1 _16803_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][19] ),
    .S(_03203_),
    .Z(_03249_));
 MUX2_X1 _16804_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][19] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][19] ),
    .S(_02832_),
    .Z(_03250_));
 MUX2_X1 _16805_ (.A(_03249_),
    .B(_03250_),
    .S(_03206_),
    .Z(_03251_));
 MUX2_X1 _16806_ (.A(_03248_),
    .B(_03251_),
    .S(_02836_),
    .Z(_03252_));
 OAI21_X4 _16807_ (.A(_03245_),
    .B1(_03252_),
    .B2(_02839_),
    .ZN(_03253_));
 NOR2_X1 _16808_ (.A1(_02804_),
    .A2(_03253_),
    .ZN(_03254_));
 NOR3_X2 _16809_ (.A1(_03221_),
    .A2(_03236_),
    .A3(_03254_),
    .ZN(_03255_));
 NOR2_X2 _16810_ (.A1(_02760_),
    .A2(_03255_),
    .ZN(net310));
 MUX2_X1 _16811_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][1] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][1] ),
    .S(_02763_),
    .Z(_03256_));
 OR2_X1 _16812_ (.A1(_02762_),
    .A2(_03256_),
    .ZN(_03257_));
 MUX2_X1 _16813_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][1] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][1] ),
    .S(_02938_),
    .Z(_03258_));
 OAI21_X4 _16814_ (.A(_03257_),
    .B1(_03258_),
    .B2(_02767_),
    .ZN(_03259_));
 MUX2_X1 _16815_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][1] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][1] ),
    .S(_03068_),
    .Z(_03260_));
 INV_X1 _16816_ (.A(_03260_),
    .ZN(_03261_));
 NAND2_X1 _16817_ (.A1(_02769_),
    .A2(_03261_),
    .ZN(_03262_));
 MUX2_X1 _16818_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][1] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][1] ),
    .S(_02774_),
    .Z(_03263_));
 OAI21_X4 _16819_ (.A(_03262_),
    .B1(_03263_),
    .B2(_02776_),
    .ZN(_03264_));
 OAI22_X1 _16820_ (.A1(_03015_),
    .A2(_03259_),
    .B1(_03264_),
    .B2(_03025_),
    .ZN(_03265_));
 MUX2_X1 _16821_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][1] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][1] ),
    .S(_02785_),
    .Z(_03266_));
 OR2_X1 _16822_ (.A1(_02784_),
    .A2(_03266_),
    .ZN(_03267_));
 MUX2_X1 _16823_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][1] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][1] ),
    .S(_07440_),
    .Z(_03268_));
 OAI21_X4 _16824_ (.A(_03267_),
    .B1(_03268_),
    .B2(_02789_),
    .ZN(_03269_));
 MUX2_X1 _16825_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][1] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][1] ),
    .S(_03184_),
    .Z(_03270_));
 OR2_X1 _16826_ (.A1(_02791_),
    .A2(_03270_),
    .ZN(_03271_));
 MUX2_X1 _16827_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][1] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][1] ),
    .S(_02795_),
    .Z(_03272_));
 OAI21_X4 _16828_ (.A(_03271_),
    .B1(_03272_),
    .B2(_02797_),
    .ZN(_03273_));
 OAI22_X1 _16829_ (.A1(_02783_),
    .A2(_03269_),
    .B1(_03273_),
    .B2(_02801_),
    .ZN(_03274_));
 MUX2_X1 _16830_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][1] ),
    .S(_02808_),
    .Z(_03275_));
 MUX2_X1 _16831_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][1] ),
    .S(_03191_),
    .Z(_03276_));
 BUF_X4 _16832_ (.A(_05710_),
    .Z(_03277_));
 MUX2_X1 _16833_ (.A(_03275_),
    .B(_03276_),
    .S(_03277_),
    .Z(_03278_));
 NAND2_X1 _16834_ (.A1(_02806_),
    .A2(_03278_),
    .ZN(_03279_));
 BUF_X4 _16835_ (.A(_02807_),
    .Z(_03280_));
 MUX2_X1 _16836_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][1] ),
    .S(_03280_),
    .Z(_03281_));
 MUX2_X1 _16837_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][1] ),
    .S(_03042_),
    .Z(_03282_));
 MUX2_X1 _16838_ (.A(_03281_),
    .B(_03282_),
    .S(_02820_),
    .Z(_03283_));
 NAND2_X1 _16839_ (.A1(_02815_),
    .A2(_03283_),
    .ZN(_03284_));
 NAND3_X2 _16840_ (.A1(_03036_),
    .A2(_03279_),
    .A3(_03284_),
    .ZN(_03285_));
 MUX2_X1 _16841_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][1] ),
    .S(_03047_),
    .Z(_03286_));
 MUX2_X1 _16842_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][1] ),
    .S(_02826_),
    .Z(_03287_));
 MUX2_X1 _16843_ (.A(_03286_),
    .B(_03287_),
    .S(_02828_),
    .Z(_03288_));
 MUX2_X1 _16844_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][1] ),
    .S(_03203_),
    .Z(_03289_));
 MUX2_X1 _16845_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][1] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][1] ),
    .S(_02832_),
    .Z(_03290_));
 MUX2_X1 _16846_ (.A(_03289_),
    .B(_03290_),
    .S(_03206_),
    .Z(_03291_));
 BUF_X4 _16847_ (.A(_05720_),
    .Z(_03292_));
 MUX2_X1 _16848_ (.A(_03288_),
    .B(_03291_),
    .S(_03292_),
    .Z(_03293_));
 OAI21_X4 _16849_ (.A(_03285_),
    .B1(_03293_),
    .B2(_02839_),
    .ZN(_03294_));
 NOR2_X1 _16850_ (.A1(_02804_),
    .A2(_03294_),
    .ZN(_03295_));
 NOR3_X1 _16851_ (.A1(_03265_),
    .A2(_03274_),
    .A3(_03295_),
    .ZN(_03296_));
 NOR2_X1 _16852_ (.A1(_02760_),
    .A2(_03296_),
    .ZN(net311));
 MUX2_X1 _16853_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][20] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][20] ),
    .S(_02770_),
    .Z(_03297_));
 INV_X1 _16854_ (.A(_03297_),
    .ZN(_03298_));
 NAND2_X1 _16855_ (.A1(_02845_),
    .A2(_03298_),
    .ZN(_03299_));
 MUX2_X1 _16856_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][20] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][20] ),
    .S(_07250_),
    .Z(_03300_));
 OAI21_X4 _16857_ (.A(_03299_),
    .B1(_03300_),
    .B2(_07244_),
    .ZN(_03301_));
 MUX2_X1 _16858_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][20] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][20] ),
    .S(_07440_),
    .Z(_03302_));
 OR2_X1 _16859_ (.A1(_07439_),
    .A2(_03302_),
    .ZN(_03303_));
 MUX2_X1 _16860_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][20] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][20] ),
    .S(_07443_),
    .Z(_03304_));
 OAI21_X4 _16861_ (.A(_03303_),
    .B1(_03304_),
    .B2(_07446_),
    .ZN(_03305_));
 OAI22_X1 _16862_ (.A1(_02844_),
    .A2(_03301_),
    .B1(_03305_),
    .B2(_02906_),
    .ZN(_03306_));
 MUX2_X1 _16863_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][20] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][20] ),
    .S(_02763_),
    .Z(_03307_));
 OR2_X1 _16864_ (.A1(_07519_),
    .A2(_03307_),
    .ZN(_03308_));
 MUX2_X1 _16865_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][20] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][20] ),
    .S(_07523_),
    .Z(_03309_));
 OAI21_X4 _16866_ (.A(_03308_),
    .B1(_03309_),
    .B2(_07526_),
    .ZN(_03310_));
 MUX2_X1 _16867_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][20] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][20] ),
    .S(_02792_),
    .Z(_03311_));
 OR2_X1 _16868_ (.A1(_02991_),
    .A2(_03311_),
    .ZN(_03312_));
 MUX2_X1 _16869_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][20] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][20] ),
    .S(_07497_),
    .Z(_03313_));
 OAI21_X4 _16870_ (.A(_03312_),
    .B1(_03313_),
    .B2(_02995_),
    .ZN(_03314_));
 OAI22_X1 _16871_ (.A1(_02761_),
    .A2(_03310_),
    .B1(_03314_),
    .B2(_02801_),
    .ZN(_03315_));
 NOR2_X1 _16872_ (.A1(_03306_),
    .A2(_03315_),
    .ZN(_03316_));
 MUX2_X1 _16873_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][20] ),
    .S(_02810_),
    .Z(_03317_));
 MUX2_X1 _16874_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][20] ),
    .S(_02875_),
    .Z(_03318_));
 MUX2_X1 _16875_ (.A(_03317_),
    .B(_03318_),
    .S(_02812_),
    .Z(_03319_));
 MUX2_X1 _16876_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][20] ),
    .S(_02875_),
    .Z(_03320_));
 MUX2_X1 _16877_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][20] ),
    .S(_02882_),
    .Z(_03321_));
 MUX2_X1 _16878_ (.A(_03320_),
    .B(_03321_),
    .S(_02879_),
    .Z(_03322_));
 MUX2_X1 _16879_ (.A(_03319_),
    .B(_03322_),
    .S(_02836_),
    .Z(_03323_));
 MUX2_X1 _16880_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][20] ),
    .S(_02877_),
    .Z(_03324_));
 MUX2_X1 _16881_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][20] ),
    .S(_02929_),
    .Z(_03325_));
 MUX2_X1 _16882_ (.A(_03324_),
    .B(_03325_),
    .S(_02890_),
    .Z(_03326_));
 MUX2_X1 _16883_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][20] ),
    .S(_02929_),
    .Z(_03327_));
 MUX2_X1 _16884_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][20] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][20] ),
    .S(_02888_),
    .Z(_03328_));
 MUX2_X1 _16885_ (.A(_03327_),
    .B(_03328_),
    .S(_02890_),
    .Z(_03329_));
 MUX2_X1 _16886_ (.A(_03326_),
    .B(_03329_),
    .S(_02885_),
    .Z(_03330_));
 MUX2_X2 _16887_ (.A(_03323_),
    .B(_03330_),
    .S(_07393_),
    .Z(_03331_));
 NAND2_X1 _16888_ (.A1(_02874_),
    .A2(_03331_),
    .ZN(_03332_));
 AOI21_X2 _16889_ (.A(_02843_),
    .B1(_03316_),
    .B2(_03332_),
    .ZN(net312));
 MUX2_X1 _16890_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][21] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][21] ),
    .S(_03223_),
    .Z(_03333_));
 OR2_X1 _16891_ (.A1(_02762_),
    .A2(_03333_),
    .ZN(_03334_));
 MUX2_X1 _16892_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][21] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][21] ),
    .S(_02938_),
    .Z(_03335_));
 OAI21_X4 _16893_ (.A(_03334_),
    .B1(_03335_),
    .B2(_02767_),
    .ZN(_03336_));
 MUX2_X1 _16894_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][21] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][21] ),
    .S(_03068_),
    .Z(_03337_));
 INV_X1 _16895_ (.A(_03337_),
    .ZN(_03338_));
 NAND2_X1 _16896_ (.A1(_02941_),
    .A2(_03338_),
    .ZN(_03339_));
 MUX2_X1 _16897_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][21] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][21] ),
    .S(_02774_),
    .Z(_03340_));
 OAI21_X4 _16898_ (.A(_03339_),
    .B1(_03340_),
    .B2(_02769_),
    .ZN(_03341_));
 OAI22_X1 _16899_ (.A1(_03015_),
    .A2(_03336_),
    .B1(_03341_),
    .B2(_03025_),
    .ZN(_03342_));
 MUX2_X1 _16900_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][21] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][21] ),
    .S(_02785_),
    .Z(_03343_));
 OR2_X1 _16901_ (.A1(_02784_),
    .A2(_03343_),
    .ZN(_03344_));
 MUX2_X1 _16902_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][21] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][21] ),
    .S(_02950_),
    .Z(_03345_));
 OAI21_X4 _16903_ (.A(_03344_),
    .B1(_03345_),
    .B2(_02789_),
    .ZN(_03346_));
 MUX2_X1 _16904_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][21] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][21] ),
    .S(_03184_),
    .Z(_03347_));
 OR2_X1 _16905_ (.A1(_02791_),
    .A2(_03347_),
    .ZN(_03348_));
 MUX2_X1 _16906_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][21] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][21] ),
    .S(_02795_),
    .Z(_03349_));
 OAI21_X4 _16907_ (.A(_03348_),
    .B1(_03349_),
    .B2(_02797_),
    .ZN(_03350_));
 CLKBUF_X3 _16908_ (.A(_02800_),
    .Z(_03351_));
 OAI22_X1 _16909_ (.A1(_02783_),
    .A2(_03346_),
    .B1(_03350_),
    .B2(_03351_),
    .ZN(_03352_));
 MUX2_X1 _16910_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][21] ),
    .S(_02808_),
    .Z(_03353_));
 MUX2_X1 _16911_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][21] ),
    .S(_03191_),
    .Z(_03354_));
 MUX2_X1 _16912_ (.A(_03353_),
    .B(_03354_),
    .S(_03277_),
    .Z(_03355_));
 NAND2_X1 _16913_ (.A1(_02806_),
    .A2(_03355_),
    .ZN(_03356_));
 MUX2_X1 _16914_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][21] ),
    .S(_03280_),
    .Z(_03357_));
 MUX2_X1 _16915_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][21] ),
    .S(_03042_),
    .Z(_03358_));
 MUX2_X1 _16916_ (.A(_03357_),
    .B(_03358_),
    .S(_02820_),
    .Z(_03359_));
 NAND2_X1 _16917_ (.A1(_02815_),
    .A2(_03359_),
    .ZN(_03360_));
 NAND3_X2 _16918_ (.A1(_03036_),
    .A2(_03356_),
    .A3(_03360_),
    .ZN(_03361_));
 MUX2_X1 _16919_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][21] ),
    .S(_03047_),
    .Z(_03362_));
 MUX2_X1 _16920_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][21] ),
    .S(_02826_),
    .Z(_03363_));
 MUX2_X1 _16921_ (.A(_03362_),
    .B(_03363_),
    .S(_02828_),
    .Z(_03364_));
 MUX2_X1 _16922_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][21] ),
    .S(_03203_),
    .Z(_03365_));
 MUX2_X1 _16923_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][21] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][21] ),
    .S(_02832_),
    .Z(_03366_));
 MUX2_X1 _16924_ (.A(_03365_),
    .B(_03366_),
    .S(_03206_),
    .Z(_03367_));
 MUX2_X1 _16925_ (.A(_03364_),
    .B(_03367_),
    .S(_03292_),
    .Z(_03368_));
 OAI21_X4 _16926_ (.A(_03361_),
    .B1(_03368_),
    .B2(_02839_),
    .ZN(_03369_));
 NOR2_X1 _16927_ (.A1(_02804_),
    .A2(_03369_),
    .ZN(_03370_));
 NOR3_X1 _16928_ (.A1(_03342_),
    .A2(_03352_),
    .A3(_03370_),
    .ZN(_03371_));
 NOR2_X1 _16929_ (.A1(_02760_),
    .A2(_03371_),
    .ZN(net313));
 INV_X4 _16930_ (.A(_02778_),
    .ZN(_03372_));
 AOI22_X1 _16931_ (.A1(_06996_),
    .A2(_05775_),
    .B1(_06080_),
    .B2(_03372_),
    .ZN(_03373_));
 INV_X2 _16932_ (.A(_05815_),
    .ZN(_03374_));
 OAI221_X1 _16933_ (.A(_03373_),
    .B1(_02494_),
    .B2(_03351_),
    .C1(_03066_),
    .C2(_03374_),
    .ZN(_03375_));
 BUF_X4 _16934_ (.A(_02872_),
    .Z(_03376_));
 AOI21_X1 _16935_ (.A(_03375_),
    .B1(_07132_),
    .B2(_03376_),
    .ZN(_03377_));
 NOR2_X1 _16936_ (.A1(_02760_),
    .A2(_03377_),
    .ZN(net314));
 INV_X2 _16937_ (.A(_02799_),
    .ZN(_03378_));
 BUF_X4 _16938_ (.A(_03378_),
    .Z(_03379_));
 BUF_X4 _16939_ (.A(_05157_),
    .Z(_03380_));
 AOI22_X1 _16940_ (.A1(_03379_),
    .A2(_05849_),
    .B1(_05796_),
    .B2(_03380_),
    .ZN(_03381_));
 INV_X2 _16941_ (.A(_06060_),
    .ZN(_03382_));
 INV_X2 _16942_ (.A(_05765_),
    .ZN(_03383_));
 OAI221_X1 _16943_ (.A(_03381_),
    .B1(_03382_),
    .B2(_02779_),
    .C1(_02855_),
    .C2(_03383_),
    .ZN(_03384_));
 AOI21_X1 _16944_ (.A(_03384_),
    .B1(_07156_),
    .B2(_03376_),
    .ZN(_03385_));
 NOR2_X1 _16945_ (.A1(_02760_),
    .A2(_03385_),
    .ZN(net315));
 CLKBUF_X3 _16946_ (.A(_05163_),
    .Z(_03386_));
 AOI22_X1 _16947_ (.A1(_03379_),
    .A2(_05839_),
    .B1(_05799_),
    .B2(_05157_),
    .ZN(_03387_));
 INV_X1 _16948_ (.A(_06064_),
    .ZN(_03388_));
 INV_X2 _16949_ (.A(_05771_),
    .ZN(_03389_));
 OAI221_X1 _16950_ (.A(_03387_),
    .B1(_03388_),
    .B2(_02779_),
    .C1(_02855_),
    .C2(_03389_),
    .ZN(_03390_));
 AOI21_X1 _16951_ (.A(_03390_),
    .B1(_05956_),
    .B2(_03376_),
    .ZN(_03391_));
 NOR2_X1 _16952_ (.A1(_03386_),
    .A2(_03391_),
    .ZN(net316));
 AOI22_X1 _16953_ (.A1(_03379_),
    .A2(_05829_),
    .B1(_05802_),
    .B2(_05157_),
    .ZN(_03392_));
 INV_X1 _16954_ (.A(_06067_),
    .ZN(_03393_));
 BUF_X4 _16955_ (.A(_06960_),
    .Z(_03394_));
 INV_X1 _16956_ (.A(_05768_),
    .ZN(_03395_));
 OAI221_X1 _16957_ (.A(_03392_),
    .B1(_03393_),
    .B2(_02779_),
    .C1(_03394_),
    .C2(_03395_),
    .ZN(_03396_));
 AOI21_X1 _16958_ (.A(_03396_),
    .B1(_05902_),
    .B2(_03376_),
    .ZN(_03397_));
 NOR2_X1 _16959_ (.A1(_03386_),
    .A2(_03397_),
    .ZN(net317));
 AOI22_X1 _16960_ (.A1(_03379_),
    .A2(_05832_),
    .B1(_05792_),
    .B2(_05157_),
    .ZN(_03398_));
 INV_X1 _16961_ (.A(_06056_),
    .ZN(_03399_));
 INV_X1 _16962_ (.A(_05760_),
    .ZN(_03400_));
 OAI221_X1 _16963_ (.A(_03398_),
    .B1(_03399_),
    .B2(_02779_),
    .C1(_03394_),
    .C2(_03400_),
    .ZN(_03401_));
 OR2_X1 _16964_ (.A1(_05922_),
    .A2(_05932_),
    .ZN(_03402_));
 OAI21_X4 _16965_ (.A(_03402_),
    .B1(_05918_),
    .B2(_07337_),
    .ZN(_03403_));
 AOI21_X1 _16966_ (.A(_03401_),
    .B1(_03403_),
    .B2(_03376_),
    .ZN(_03404_));
 NOR2_X1 _16967_ (.A1(_03386_),
    .A2(_03404_),
    .ZN(net318));
 OAI22_X2 _16968_ (.A1(_06959_),
    .A2(_07233_),
    .B1(_07196_),
    .B2(_02778_),
    .ZN(_03405_));
 AOI221_X2 _16969_ (.A(_03405_),
    .B1(_05836_),
    .B2(_03379_),
    .C1(_03380_),
    .C2(_05809_),
    .ZN(_03406_));
 NAND2_X1 _16970_ (.A1(_02874_),
    .A2(_05972_),
    .ZN(_03407_));
 AOI21_X2 _16971_ (.A(_02843_),
    .B1(_03406_),
    .B2(_03407_),
    .ZN(net319));
 OAI22_X2 _16972_ (.A1(_06959_),
    .A2(_07229_),
    .B1(_07192_),
    .B2(_02778_),
    .ZN(_03408_));
 AOI221_X2 _16973_ (.A(_03408_),
    .B1(_05843_),
    .B2(_03379_),
    .C1(_03380_),
    .C2(_05806_),
    .ZN(_03409_));
 NAND2_X1 _16974_ (.A1(_02874_),
    .A2(_06008_),
    .ZN(_03410_));
 AOI21_X2 _16975_ (.A(_02843_),
    .B1(_03409_),
    .B2(_03410_),
    .ZN(net320));
 AOI22_X1 _16976_ (.A1(_06724_),
    .A2(_05778_),
    .B1(_06071_),
    .B2(_03372_),
    .ZN(_03411_));
 INV_X2 _16977_ (.A(_05812_),
    .ZN(_03412_));
 OAI221_X1 _16978_ (.A(_03411_),
    .B1(_07105_),
    .B2(_03351_),
    .C1(_03066_),
    .C2(_03412_),
    .ZN(_03413_));
 AOI21_X1 _16979_ (.A(_03413_),
    .B1(_05993_),
    .B2(_03376_),
    .ZN(_03414_));
 NOR2_X1 _16980_ (.A1(_03386_),
    .A2(_03414_),
    .ZN(net321));
 MUX2_X1 _16981_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][2] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][2] ),
    .S(_03223_),
    .Z(_03415_));
 OR2_X1 _16982_ (.A1(_02762_),
    .A2(_03415_),
    .ZN(_03416_));
 MUX2_X1 _16983_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][2] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][2] ),
    .S(_02938_),
    .Z(_03417_));
 OAI21_X4 _16984_ (.A(_03416_),
    .B1(_03417_),
    .B2(_02767_),
    .ZN(_03418_));
 MUX2_X1 _16985_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][2] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][2] ),
    .S(_02859_),
    .Z(_03419_));
 OR2_X1 _16986_ (.A1(_02858_),
    .A2(_03419_),
    .ZN(_03420_));
 MUX2_X1 _16987_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][2] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][2] ),
    .S(_02950_),
    .Z(_03421_));
 OAI21_X4 _16988_ (.A(_03420_),
    .B1(_03421_),
    .B2(_02789_),
    .ZN(_03422_));
 OAI22_X1 _16989_ (.A1(_03015_),
    .A2(_03418_),
    .B1(_03422_),
    .B2(_02782_),
    .ZN(_03423_));
 MUX2_X1 _16990_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][2] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][2] ),
    .S(_03068_),
    .Z(_03424_));
 INV_X1 _16991_ (.A(_03424_),
    .ZN(_03425_));
 NAND2_X1 _16992_ (.A1(_02941_),
    .A2(_03425_),
    .ZN(_03426_));
 MUX2_X1 _16993_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][2] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][2] ),
    .S(_07246_),
    .Z(_03427_));
 OAI21_X4 _16994_ (.A(_03426_),
    .B1(_03427_),
    .B2(_02769_),
    .ZN(_03428_));
 MUX2_X1 _16995_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][2] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][2] ),
    .S(_03184_),
    .Z(_03429_));
 OR2_X1 _16996_ (.A1(_07488_),
    .A2(_03429_),
    .ZN(_03430_));
 MUX2_X1 _16997_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][2] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][2] ),
    .S(_02795_),
    .Z(_03431_));
 OAI21_X4 _16998_ (.A(_03430_),
    .B1(_03431_),
    .B2(_07499_),
    .ZN(_03432_));
 OAI22_X1 _16999_ (.A1(_02780_),
    .A2(_03428_),
    .B1(_03432_),
    .B2(_03351_),
    .ZN(_03433_));
 MUX2_X1 _17000_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][2] ),
    .S(_02818_),
    .Z(_03434_));
 MUX2_X1 _17001_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][2] ),
    .S(_03191_),
    .Z(_03435_));
 MUX2_X1 _17002_ (.A(_03434_),
    .B(_03435_),
    .S(_03277_),
    .Z(_03436_));
 NAND2_X1 _17003_ (.A1(_02806_),
    .A2(_03436_),
    .ZN(_03437_));
 MUX2_X1 _17004_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][2] ),
    .S(_03280_),
    .Z(_03438_));
 MUX2_X1 _17005_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][2] ),
    .S(_03042_),
    .Z(_03439_));
 MUX2_X1 _17006_ (.A(_03438_),
    .B(_03439_),
    .S(_02820_),
    .Z(_03440_));
 NAND2_X1 _17007_ (.A1(_02815_),
    .A2(_03440_),
    .ZN(_03441_));
 NAND3_X2 _17008_ (.A1(_03036_),
    .A2(_03437_),
    .A3(_03441_),
    .ZN(_03442_));
 MUX2_X1 _17009_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][2] ),
    .S(_03047_),
    .Z(_03443_));
 MUX2_X1 _17010_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][2] ),
    .S(_02824_),
    .Z(_03444_));
 MUX2_X1 _17011_ (.A(_03443_),
    .B(_03444_),
    .S(_07336_),
    .Z(_03445_));
 MUX2_X1 _17012_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][2] ),
    .S(_03203_),
    .Z(_03446_));
 MUX2_X1 _17013_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][2] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][2] ),
    .S(_02832_),
    .Z(_03447_));
 MUX2_X1 _17014_ (.A(_03446_),
    .B(_03447_),
    .S(_03206_),
    .Z(_03448_));
 MUX2_X1 _17015_ (.A(_03445_),
    .B(_03448_),
    .S(_03292_),
    .Z(_03449_));
 OAI21_X4 _17016_ (.A(_03442_),
    .B1(_02805_),
    .B2(_03449_),
    .ZN(_03450_));
 NOR2_X1 _17017_ (.A1(_02804_),
    .A2(_03450_),
    .ZN(_03451_));
 NOR3_X1 _17018_ (.A1(_03423_),
    .A2(_03433_),
    .A3(_03451_),
    .ZN(_03452_));
 NOR2_X1 _17019_ (.A1(_03386_),
    .A2(_03452_),
    .ZN(net322));
 AOI22_X2 _17020_ (.A1(_03379_),
    .A2(_06524_),
    .B1(_05492_),
    .B2(_06724_),
    .ZN(_03453_));
 OAI221_X2 _17021_ (.A(_03453_),
    .B1(_06099_),
    .B2(_02779_),
    .C1(_03066_),
    .C2(_05274_),
    .ZN(_03454_));
 AOI21_X1 _17022_ (.A(_03454_),
    .B1(_06179_),
    .B2(_03376_),
    .ZN(_03455_));
 NOR2_X1 _17023_ (.A1(_03386_),
    .A2(_03455_),
    .ZN(net323));
 AOI22_X1 _17024_ (.A1(_03380_),
    .A2(_06514_),
    .B1(_06100_),
    .B2(_03372_),
    .ZN(_03456_));
 OAI221_X1 _17025_ (.A(_03456_),
    .B1(_05376_),
    .B2(_02800_),
    .C1(_03394_),
    .C2(_06789_),
    .ZN(_03457_));
 AOI21_X1 _17026_ (.A(_03457_),
    .B1(_06146_),
    .B2(_03376_),
    .ZN(_03458_));
 NOR2_X1 _17027_ (.A1(_03386_),
    .A2(_03458_),
    .ZN(net324));
 OAI22_X2 _17028_ (.A1(_02782_),
    .A2(_06513_),
    .B1(_06098_),
    .B2(_02778_),
    .ZN(_03459_));
 AOI221_X2 _17029_ (.A(_03459_),
    .B1(_05370_),
    .B2(_03379_),
    .C1(_06996_),
    .C2(_05500_),
    .ZN(_03460_));
 NAND2_X1 _17030_ (.A1(_02874_),
    .A2(_06163_),
    .ZN(_03461_));
 AOI21_X2 _17031_ (.A(_02843_),
    .B1(_03460_),
    .B2(_03461_),
    .ZN(net325));
 MUX2_X1 _17032_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][33] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][33] ),
    .S(_03223_),
    .Z(_03462_));
 OR2_X1 _17033_ (.A1(_02762_),
    .A2(_03462_),
    .ZN(_03463_));
 MUX2_X1 _17034_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][33] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][33] ),
    .S(_02938_),
    .Z(_03464_));
 OAI21_X4 _17035_ (.A(_03463_),
    .B1(_03464_),
    .B2(_02767_),
    .ZN(_03465_));
 MUX2_X1 _17036_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][33] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][33] ),
    .S(_02770_),
    .Z(_03466_));
 INV_X1 _17037_ (.A(_03466_),
    .ZN(_03467_));
 NAND2_X1 _17038_ (.A1(_02776_),
    .A2(_03467_),
    .ZN(_03468_));
 MUX2_X1 _17039_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][33] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][33] ),
    .S(_02774_),
    .Z(_03469_));
 BUF_X8 _17040_ (.A(_07244_),
    .Z(_03470_));
 OAI21_X4 _17041_ (.A(_03468_),
    .B1(_03469_),
    .B2(_03470_),
    .ZN(_03471_));
 OAI22_X1 _17042_ (.A1(_03015_),
    .A2(_03465_),
    .B1(_03471_),
    .B2(_03025_),
    .ZN(_03472_));
 MUX2_X1 _17043_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][33] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][33] ),
    .S(_02785_),
    .Z(_03473_));
 OR2_X1 _17044_ (.A1(_05153_),
    .A2(_03473_),
    .ZN(_03474_));
 MUX2_X1 _17045_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][33] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][33] ),
    .S(_07440_),
    .Z(_03475_));
 OAI21_X4 _17046_ (.A(_03474_),
    .B1(_03475_),
    .B2(_07445_),
    .ZN(_03476_));
 MUX2_X1 _17047_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][33] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][33] ),
    .S(_03184_),
    .Z(_03477_));
 OR2_X1 _17048_ (.A1(_07488_),
    .A2(_03477_),
    .ZN(_03478_));
 MUX2_X1 _17049_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][33] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][33] ),
    .S(_02795_),
    .Z(_03479_));
 OAI21_X4 _17050_ (.A(_03478_),
    .B1(_03479_),
    .B2(_07499_),
    .ZN(_03480_));
 OAI22_X1 _17051_ (.A1(_02783_),
    .A2(_03476_),
    .B1(_03480_),
    .B2(_03351_),
    .ZN(_03481_));
 MUX2_X1 _17052_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][33] ),
    .S(_02818_),
    .Z(_03482_));
 MUX2_X1 _17053_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][33] ),
    .S(_03191_),
    .Z(_03483_));
 MUX2_X1 _17054_ (.A(_03482_),
    .B(_03483_),
    .S(_03277_),
    .Z(_03484_));
 NAND2_X1 _17055_ (.A1(_02806_),
    .A2(_03484_),
    .ZN(_03485_));
 MUX2_X1 _17056_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][33] ),
    .S(_03280_),
    .Z(_03486_));
 MUX2_X1 _17057_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][33] ),
    .S(_03042_),
    .Z(_03487_));
 MUX2_X1 _17058_ (.A(_03486_),
    .B(_03487_),
    .S(_02820_),
    .Z(_03488_));
 NAND2_X1 _17059_ (.A1(_07391_),
    .A2(_03488_),
    .ZN(_03489_));
 NAND3_X2 _17060_ (.A1(_03036_),
    .A2(_03485_),
    .A3(_03489_),
    .ZN(_03490_));
 MUX2_X1 _17061_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][33] ),
    .S(_03047_),
    .Z(_03491_));
 MUX2_X1 _17062_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][33] ),
    .S(_02824_),
    .Z(_03492_));
 MUX2_X1 _17063_ (.A(_03491_),
    .B(_03492_),
    .S(_07336_),
    .Z(_03493_));
 MUX2_X1 _17064_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][33] ),
    .S(_03203_),
    .Z(_03494_));
 MUX2_X1 _17065_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][33] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][33] ),
    .S(_02832_),
    .Z(_03495_));
 MUX2_X1 _17066_ (.A(_03494_),
    .B(_03495_),
    .S(_03206_),
    .Z(_03496_));
 MUX2_X1 _17067_ (.A(_03493_),
    .B(_03496_),
    .S(_03292_),
    .Z(_03497_));
 OAI21_X4 _17068_ (.A(_03490_),
    .B1(_03497_),
    .B2(_02805_),
    .ZN(_03498_));
 NOR2_X1 _17069_ (.A1(_02804_),
    .A2(_03498_),
    .ZN(_03499_));
 NOR3_X1 _17070_ (.A1(_03472_),
    .A2(_03481_),
    .A3(_03499_),
    .ZN(_03500_));
 NOR2_X1 _17071_ (.A1(_03386_),
    .A2(_03500_),
    .ZN(net326));
 BUF_X8 _17072_ (.A(_05163_),
    .Z(_03501_));
 INV_X2 _17073_ (.A(_10252_),
    .ZN(_03502_));
 OAI22_X2 _17074_ (.A1(_05156_),
    .A2(_03502_),
    .B1(_05327_),
    .B2(_02800_),
    .ZN(_03503_));
 AOI221_X2 _17075_ (.A(_03503_),
    .B1(_10225_),
    .B2(_03372_),
    .C1(_06996_),
    .C2(_10348_),
    .ZN(_03504_));
 NAND2_X1 _17076_ (.A1(_02874_),
    .A2(_10417_),
    .ZN(_03505_));
 AOI21_X4 _17077_ (.A(_03501_),
    .B1(_03504_),
    .B2(_03505_),
    .ZN(net327));
 AOI22_X1 _17078_ (.A1(_06724_),
    .A2(_07302_),
    .B1(net694),
    .B2(_03378_),
    .ZN(_03506_));
 OAI221_X1 _17079_ (.A(_03506_),
    .B1(_10221_),
    .B2(_02779_),
    .C1(_03066_),
    .C2(_10255_),
    .ZN(_03507_));
 AOI21_X1 _17080_ (.A(_03507_),
    .B1(_07676_),
    .B2(_02873_),
    .ZN(_03508_));
 NOR2_X1 _17081_ (.A1(_03386_),
    .A2(_03508_),
    .ZN(net328));
 OAI22_X2 _17082_ (.A1(_05156_),
    .A2(_10261_),
    .B1(_10315_),
    .B2(_02799_),
    .ZN(_03509_));
 INV_X1 _17083_ (.A(_10357_),
    .ZN(_03510_));
 AOI221_X2 _17084_ (.A(_03509_),
    .B1(_07434_),
    .B2(_03372_),
    .C1(_06996_),
    .C2(_03510_),
    .ZN(_03511_));
 CLKBUF_X3 _17085_ (.A(_02873_),
    .Z(_03512_));
 NAND2_X1 _17086_ (.A1(_03512_),
    .A2(_07661_),
    .ZN(_03513_));
 AOI21_X4 _17087_ (.A(_03501_),
    .B1(_03511_),
    .B2(_03513_),
    .ZN(net329));
 AOI22_X1 _17088_ (.A1(_03372_),
    .A2(net742),
    .B1(_07305_),
    .B2(_06724_),
    .ZN(_03514_));
 OAI221_X1 _17089_ (.A(_03514_),
    .B1(_10312_),
    .B2(_02800_),
    .C1(_03066_),
    .C2(_10258_),
    .ZN(_03515_));
 AOI21_X1 _17090_ (.A(_03515_),
    .B1(_07409_),
    .B2(_02873_),
    .ZN(_03516_));
 NOR2_X1 _17091_ (.A1(_03386_),
    .A2(_03516_),
    .ZN(net330));
 OAI22_X2 _17092_ (.A1(_05156_),
    .A2(_10273_),
    .B1(net697),
    .B2(_02799_),
    .ZN(_03517_));
 INV_X1 _17093_ (.A(_10369_),
    .ZN(_03518_));
 AOI221_X2 _17094_ (.A(_03517_),
    .B1(net674),
    .B2(_03372_),
    .C1(_06996_),
    .C2(_03518_),
    .ZN(_03519_));
 NAND2_X1 _17095_ (.A1(_03512_),
    .A2(_07646_),
    .ZN(_03520_));
 AOI21_X4 _17096_ (.A(_03501_),
    .B1(_03519_),
    .B2(_03520_),
    .ZN(net331));
 OAI22_X2 _17097_ (.A1(_05156_),
    .A2(_10270_),
    .B1(_10209_),
    .B2(_02778_),
    .ZN(_03521_));
 INV_X1 _17098_ (.A(_10366_),
    .ZN(_03522_));
 AOI221_X2 _17099_ (.A(_03521_),
    .B1(net665),
    .B2(_03379_),
    .C1(_06996_),
    .C2(_03522_),
    .ZN(_03523_));
 NAND2_X1 _17100_ (.A1(_03512_),
    .A2(_07631_),
    .ZN(_03524_));
 AOI21_X2 _17101_ (.A(_03501_),
    .B1(_03523_),
    .B2(_03524_),
    .ZN(net332));
 BUF_X4 _17102_ (.A(_05163_),
    .Z(_03525_));
 MUX2_X1 _17103_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][3] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][3] ),
    .S(_02770_),
    .Z(_03526_));
 INV_X1 _17104_ (.A(_03526_),
    .ZN(_03527_));
 NAND2_X1 _17105_ (.A1(_03470_),
    .A2(_03527_),
    .ZN(_03528_));
 MUX2_X1 _17106_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][3] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][3] ),
    .S(_07250_),
    .Z(_03529_));
 OAI21_X4 _17107_ (.A(_03528_),
    .B1(_03529_),
    .B2(_02845_),
    .ZN(_03530_));
 MUX2_X1 _17108_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][3] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][3] ),
    .S(_02859_),
    .Z(_03531_));
 OR2_X1 _17109_ (.A1(_02858_),
    .A2(_03531_),
    .ZN(_03532_));
 MUX2_X1 _17110_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][3] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][3] ),
    .S(_02950_),
    .Z(_03533_));
 OAI21_X4 _17111_ (.A(_03532_),
    .B1(_03533_),
    .B2(_02863_),
    .ZN(_03534_));
 OAI22_X1 _17112_ (.A1(_02780_),
    .A2(_03530_),
    .B1(_03534_),
    .B2(_02782_),
    .ZN(_03535_));
 MUX2_X1 _17113_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][3] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][3] ),
    .S(_03223_),
    .Z(_03536_));
 OR2_X1 _17114_ (.A1(_03222_),
    .A2(_03536_),
    .ZN(_03537_));
 MUX2_X1 _17115_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][3] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][3] ),
    .S(_07520_),
    .Z(_03538_));
 OAI21_X4 _17116_ (.A(_03537_),
    .B1(_03538_),
    .B2(_03227_),
    .ZN(_03539_));
 MUX2_X1 _17117_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][3] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][3] ),
    .S(_03184_),
    .Z(_03540_));
 OR2_X1 _17118_ (.A1(_07488_),
    .A2(_03540_),
    .ZN(_03541_));
 MUX2_X1 _17119_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][3] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][3] ),
    .S(_07494_),
    .Z(_03542_));
 OAI21_X4 _17120_ (.A(_03541_),
    .B1(_03542_),
    .B2(_07499_),
    .ZN(_03543_));
 OAI22_X1 _17121_ (.A1(_02855_),
    .A2(_03539_),
    .B1(_03543_),
    .B2(_03351_),
    .ZN(_03544_));
 CLKBUF_X3 _17122_ (.A(_02803_),
    .Z(_03545_));
 MUX2_X1 _17123_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][3] ),
    .S(_02818_),
    .Z(_03546_));
 MUX2_X1 _17124_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][3] ),
    .S(_03191_),
    .Z(_03547_));
 MUX2_X1 _17125_ (.A(_03546_),
    .B(_03547_),
    .S(_03277_),
    .Z(_03548_));
 NAND2_X1 _17126_ (.A1(_07130_),
    .A2(_03548_),
    .ZN(_03549_));
 MUX2_X1 _17127_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][3] ),
    .S(_03280_),
    .Z(_03550_));
 MUX2_X1 _17128_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][3] ),
    .S(_03042_),
    .Z(_03551_));
 MUX2_X1 _17129_ (.A(_03550_),
    .B(_03551_),
    .S(_02834_),
    .Z(_03552_));
 NAND2_X1 _17130_ (.A1(_07391_),
    .A2(_03552_),
    .ZN(_03553_));
 NAND3_X2 _17131_ (.A1(_03036_),
    .A2(_03549_),
    .A3(_03553_),
    .ZN(_03554_));
 MUX2_X1 _17132_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][3] ),
    .S(_03047_),
    .Z(_03555_));
 MUX2_X1 _17133_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][3] ),
    .S(_02824_),
    .Z(_03556_));
 MUX2_X1 _17134_ (.A(_03555_),
    .B(_03556_),
    .S(_07336_),
    .Z(_03557_));
 MUX2_X1 _17135_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][3] ),
    .S(_03203_),
    .Z(_03558_));
 MUX2_X1 _17136_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][3] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][3] ),
    .S(_02830_),
    .Z(_03559_));
 MUX2_X1 _17137_ (.A(_03558_),
    .B(_03559_),
    .S(_03206_),
    .Z(_03560_));
 MUX2_X1 _17138_ (.A(_03557_),
    .B(_03560_),
    .S(_03292_),
    .Z(_03561_));
 OAI21_X4 _17139_ (.A(_03554_),
    .B1(_03561_),
    .B2(_02805_),
    .ZN(_03562_));
 NOR2_X1 _17140_ (.A1(_03545_),
    .A2(_03562_),
    .ZN(_03563_));
 NOR3_X1 _17141_ (.A1(_03535_),
    .A2(_03544_),
    .A3(_03563_),
    .ZN(_03564_));
 NOR2_X2 _17142_ (.A1(_03525_),
    .A2(_03564_),
    .ZN(net333));
 OAI22_X2 _17143_ (.A1(_02778_),
    .A2(_10206_),
    .B1(_10303_),
    .B2(_02799_),
    .ZN(_03565_));
 INV_X1 _17144_ (.A(_10363_),
    .ZN(_03566_));
 AOI221_X2 _17145_ (.A(_03565_),
    .B1(_07473_),
    .B2(_03380_),
    .C1(_06996_),
    .C2(_03566_),
    .ZN(_03567_));
 NAND2_X1 _17146_ (.A1(_03512_),
    .A2(_07616_),
    .ZN(_03568_));
 AOI21_X2 _17147_ (.A(_03501_),
    .B1(_03567_),
    .B2(_03568_),
    .ZN(net334));
 OAI22_X2 _17148_ (.A1(_02857_),
    .A2(net640),
    .B1(net632),
    .B2(_03212_),
    .ZN(_03569_));
 OAI22_X2 _17149_ (.A1(_02844_),
    .A2(net650),
    .B1(net713),
    .B2(_02855_),
    .ZN(_03570_));
 NOR2_X2 _17150_ (.A1(_03569_),
    .A2(_03570_),
    .ZN(_03571_));
 NAND2_X1 _17151_ (.A1(_03512_),
    .A2(_07394_),
    .ZN(_03572_));
 AOI21_X4 _17152_ (.A(_03501_),
    .B1(_03571_),
    .B2(_03572_),
    .ZN(net335));
 AOI22_X1 _17153_ (.A1(_03380_),
    .A2(_10249_),
    .B1(_10276_),
    .B2(_03378_),
    .ZN(_03573_));
 INV_X1 _17154_ (.A(_10345_),
    .ZN(_03574_));
 OAI221_X1 _17155_ (.A(_03573_),
    .B1(net685),
    .B2(_02779_),
    .C1(_03394_),
    .C2(_03574_),
    .ZN(_03575_));
 AOI21_X1 _17156_ (.A(_03575_),
    .B1(_10372_),
    .B2(_02873_),
    .ZN(_03576_));
 NOR2_X2 _17157_ (.A1(_03525_),
    .A2(_03576_),
    .ZN(net336));
 INV_X1 _17158_ (.A(_10342_),
    .ZN(_03577_));
 INV_X1 _17159_ (.A(_10279_),
    .ZN(_03578_));
 AOI22_X1 _17160_ (.A1(_06724_),
    .A2(_03577_),
    .B1(_03578_),
    .B2(_03378_),
    .ZN(_03579_));
 OAI221_X1 _17161_ (.A(_03579_),
    .B1(net644),
    .B2(_02779_),
    .C1(_03066_),
    .C2(_10246_),
    .ZN(_03580_));
 AOI21_X1 _17162_ (.A(_03580_),
    .B1(_07556_),
    .B2(_02873_),
    .ZN(_03581_));
 NOR2_X2 _17163_ (.A1(_03525_),
    .A2(_03581_),
    .ZN(net337));
 OAI22_X2 _17164_ (.A1(_02778_),
    .A2(net645),
    .B1(net723),
    .B2(_06959_),
    .ZN(_03582_));
 INV_X2 _17165_ (.A(_10243_),
    .ZN(_03583_));
 AOI221_X2 _17166_ (.A(_03582_),
    .B1(net690),
    .B2(_03378_),
    .C1(_03380_),
    .C2(_03583_),
    .ZN(_03584_));
 NAND2_X1 _17167_ (.A1(_03512_),
    .A2(_07571_),
    .ZN(_03585_));
 AOI21_X4 _17168_ (.A(_03501_),
    .B1(_03584_),
    .B2(_03585_),
    .ZN(net338));
 INV_X1 _17169_ (.A(_10240_),
    .ZN(_03586_));
 AOI22_X1 _17170_ (.A1(_03380_),
    .A2(_03586_),
    .B1(_07296_),
    .B2(_06724_),
    .ZN(_03587_));
 OAI221_X1 _17171_ (.A(_03587_),
    .B1(_10285_),
    .B2(_02800_),
    .C1(_02780_),
    .C2(_10185_),
    .ZN(_03588_));
 AOI21_X1 _17172_ (.A(_03588_),
    .B1(_07342_),
    .B2(_02873_),
    .ZN(_03589_));
 NOR2_X1 _17173_ (.A1(_03525_),
    .A2(_03589_),
    .ZN(net339));
 INV_X2 _17174_ (.A(_10237_),
    .ZN(_03590_));
 AOI22_X1 _17175_ (.A1(_06724_),
    .A2(net651),
    .B1(_03590_),
    .B2(_05157_),
    .ZN(_03591_));
 OAI221_X1 _17176_ (.A(_03591_),
    .B1(_10288_),
    .B2(_02800_),
    .C1(_02780_),
    .C2(net648),
    .ZN(_03592_));
 AOI21_X1 _17177_ (.A(_03592_),
    .B1(_07376_),
    .B2(_02873_),
    .ZN(_03593_));
 NOR2_X1 _17178_ (.A1(_03525_),
    .A2(_03593_),
    .ZN(net340));
 OAI22_X1 _17179_ (.A1(_02844_),
    .A2(_10197_),
    .B1(_10234_),
    .B2(_02906_),
    .ZN(_03594_));
 OAI22_X1 _17180_ (.A1(_02761_),
    .A2(net704),
    .B1(_10291_),
    .B2(_02801_),
    .ZN(_03595_));
 NOR2_X1 _17181_ (.A1(_03594_),
    .A2(_03595_),
    .ZN(_03596_));
 NAND2_X1 _17182_ (.A1(_03512_),
    .A2(_07361_),
    .ZN(_03597_));
 AOI21_X2 _17183_ (.A(_03501_),
    .B1(_03596_),
    .B2(_03597_),
    .ZN(net341));
 OAI22_X2 _17184_ (.A1(_05156_),
    .A2(_10231_),
    .B1(_10294_),
    .B2(_02799_),
    .ZN(_03598_));
 INV_X2 _17185_ (.A(_10327_),
    .ZN(_03599_));
 AOI221_X2 _17186_ (.A(_03598_),
    .B1(net754),
    .B2(_03372_),
    .C1(_06996_),
    .C2(_03599_),
    .ZN(_03600_));
 NAND2_X1 _17187_ (.A1(_03512_),
    .A2(_07601_),
    .ZN(_03601_));
 AOI21_X4 _17188_ (.A(_03501_),
    .B1(_03600_),
    .B2(_03601_),
    .ZN(net342));
 OAI22_X1 _17189_ (.A1(_02857_),
    .A2(net731),
    .B1(_10297_),
    .B2(_03212_),
    .ZN(_03602_));
 OAI22_X1 _17190_ (.A1(_02844_),
    .A2(_10191_),
    .B1(net670),
    .B2(_02855_),
    .ZN(_03603_));
 NOR2_X1 _17191_ (.A1(_03602_),
    .A2(_03603_),
    .ZN(_03604_));
 NAND2_X1 _17192_ (.A1(_03512_),
    .A2(_07586_),
    .ZN(_03605_));
 AOI21_X2 _17193_ (.A(_03501_),
    .B1(_03604_),
    .B2(_03605_),
    .ZN(net343));
 MUX2_X1 _17194_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][4] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][4] ),
    .S(_02770_),
    .Z(_03606_));
 INV_X1 _17195_ (.A(_03606_),
    .ZN(_03607_));
 NAND2_X1 _17196_ (.A1(_02845_),
    .A2(_03607_),
    .ZN(_03608_));
 MUX2_X1 _17197_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][4] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][4] ),
    .S(_07250_),
    .Z(_03609_));
 OAI21_X4 _17198_ (.A(_03608_),
    .B1(_03609_),
    .B2(_02845_),
    .ZN(_03610_));
 MUX2_X1 _17199_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][4] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][4] ),
    .S(_07440_),
    .Z(_03611_));
 OR2_X1 _17200_ (.A1(_07439_),
    .A2(_03611_),
    .ZN(_03612_));
 MUX2_X1 _17201_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][4] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][4] ),
    .S(_07443_),
    .Z(_03613_));
 OAI21_X4 _17202_ (.A(_03612_),
    .B1(_03613_),
    .B2(_07446_),
    .ZN(_03614_));
 OAI22_X2 _17203_ (.A1(_02844_),
    .A2(_03610_),
    .B1(_03614_),
    .B2(_02906_),
    .ZN(_03615_));
 MUX2_X1 _17204_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][4] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][4] ),
    .S(_02763_),
    .Z(_03616_));
 OR2_X1 _17205_ (.A1(_07519_),
    .A2(_03616_),
    .ZN(_03617_));
 MUX2_X1 _17206_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][4] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][4] ),
    .S(_07523_),
    .Z(_03618_));
 OAI21_X4 _17207_ (.A(_03617_),
    .B1(_03618_),
    .B2(_07526_),
    .ZN(_03619_));
 MUX2_X1 _17208_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][4] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][4] ),
    .S(_02792_),
    .Z(_03620_));
 OR2_X1 _17209_ (.A1(_02991_),
    .A2(_03620_),
    .ZN(_03621_));
 MUX2_X1 _17210_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][4] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][4] ),
    .S(_02795_),
    .Z(_03622_));
 OAI21_X4 _17211_ (.A(_03621_),
    .B1(_03622_),
    .B2(_02995_),
    .ZN(_03623_));
 OAI22_X2 _17212_ (.A1(_02761_),
    .A2(_03619_),
    .B1(_03623_),
    .B2(_02801_),
    .ZN(_03624_));
 NOR2_X2 _17213_ (.A1(_03615_),
    .A2(_03624_),
    .ZN(_03625_));
 MUX2_X1 _17214_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][4] ),
    .S(_02810_),
    .Z(_03626_));
 MUX2_X1 _17215_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][4] ),
    .S(_02875_),
    .Z(_03627_));
 MUX2_X1 _17216_ (.A(_03626_),
    .B(_03627_),
    .S(_02812_),
    .Z(_03628_));
 MUX2_X1 _17217_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][4] ),
    .S(_02875_),
    .Z(_03629_));
 MUX2_X1 _17218_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][4] ),
    .S(_02882_),
    .Z(_03630_));
 MUX2_X1 _17219_ (.A(_03629_),
    .B(_03630_),
    .S(_02879_),
    .Z(_03631_));
 MUX2_X1 _17220_ (.A(_03628_),
    .B(_03631_),
    .S(_02836_),
    .Z(_03632_));
 MUX2_X1 _17221_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][4] ),
    .S(_02877_),
    .Z(_03633_));
 MUX2_X1 _17222_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][4] ),
    .S(_02929_),
    .Z(_03634_));
 MUX2_X1 _17223_ (.A(_03633_),
    .B(_03634_),
    .S(_02890_),
    .Z(_03635_));
 MUX2_X1 _17224_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][4] ),
    .S(_02882_),
    .Z(_03636_));
 MUX2_X1 _17225_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][4] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][4] ),
    .S(_02888_),
    .Z(_03637_));
 MUX2_X1 _17226_ (.A(_03636_),
    .B(_03637_),
    .S(_02890_),
    .Z(_03638_));
 MUX2_X1 _17227_ (.A(_03635_),
    .B(_03638_),
    .S(_02885_),
    .Z(_03639_));
 MUX2_X2 _17228_ (.A(_03632_),
    .B(_03639_),
    .S(_07393_),
    .Z(_03640_));
 NAND2_X1 _17229_ (.A1(_03512_),
    .A2(_03640_),
    .ZN(_03641_));
 AOI21_X4 _17230_ (.A(_05163_),
    .B1(_03625_),
    .B2(_03641_),
    .ZN(net344));
 OR2_X1 _17231_ (.A1(_07445_),
    .A2(_05248_),
    .ZN(_03642_));
 OAI21_X4 _17232_ (.A(_03642_),
    .B1(_05249_),
    .B2(_07439_),
    .ZN(_03643_));
 INV_X1 _17233_ (.A(_05682_),
    .ZN(_03644_));
 NAND2_X1 _17234_ (.A1(_02776_),
    .A2(_03644_),
    .ZN(_03645_));
 OAI21_X4 _17235_ (.A(_03645_),
    .B1(_05681_),
    .B2(_03470_),
    .ZN(_03646_));
 OAI22_X1 _17236_ (.A1(_02857_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(_03025_),
    .ZN(_03647_));
 OR2_X1 _17237_ (.A1(_02791_),
    .A2(_05429_),
    .ZN(_03648_));
 OAI21_X4 _17238_ (.A(_03648_),
    .B1(_05430_),
    .B2(_02797_),
    .ZN(_03649_));
 OR2_X1 _17239_ (.A1(_05465_),
    .A2(_05549_),
    .ZN(_03650_));
 OAI21_X4 _17240_ (.A(_03650_),
    .B1(_05551_),
    .B2(_07525_),
    .ZN(_03651_));
 OAI22_X1 _17241_ (.A1(_03212_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_06960_),
    .ZN(_03652_));
 AND2_X1 _17242_ (.A1(_02838_),
    .A2(_06448_),
    .ZN(_03653_));
 MUX2_X1 _17243_ (.A(_06272_),
    .B(_06462_),
    .S(_02836_),
    .Z(_03654_));
 AOI21_X4 _17244_ (.A(_03653_),
    .B1(_03654_),
    .B2(_05738_),
    .ZN(_03655_));
 NOR2_X1 _17245_ (.A1(_03545_),
    .A2(_03655_),
    .ZN(_03656_));
 NOR3_X1 _17246_ (.A1(_03647_),
    .A2(_03652_),
    .A3(_03656_),
    .ZN(_03657_));
 NOR2_X2 _17247_ (.A1(_03525_),
    .A2(_03657_),
    .ZN(net345));
 AOI22_X1 _17248_ (.A1(_03380_),
    .A2(_05189_),
    .B1(_05649_),
    .B2(_03372_),
    .ZN(_03658_));
 OR2_X1 _17249_ (.A1(_07488_),
    .A2(_05412_),
    .ZN(_03659_));
 OAI21_X4 _17250_ (.A(_03659_),
    .B1(_05413_),
    .B2(_07499_),
    .ZN(_03660_));
 OR2_X1 _17251_ (.A1(_05465_),
    .A2(_05530_),
    .ZN(_03661_));
 OAI21_X4 _17252_ (.A(_03661_),
    .B1(_05531_),
    .B2(_07525_),
    .ZN(_03662_));
 OAI221_X1 _17253_ (.A(_03658_),
    .B1(_03660_),
    .B2(_02800_),
    .C1(_03394_),
    .C2(_03662_),
    .ZN(_03663_));
 AOI21_X1 _17254_ (.A(_03663_),
    .B1(_06249_),
    .B2(_02873_),
    .ZN(_03664_));
 NOR2_X1 _17255_ (.A1(_03525_),
    .A2(_03664_),
    .ZN(net346));
 AND2_X1 _17256_ (.A1(_05153_),
    .A2(_05258_),
    .ZN(_03665_));
 AOI21_X4 _17257_ (.A(_03665_),
    .B1(_05259_),
    .B2(_07446_),
    .ZN(_03666_));
 INV_X1 _17258_ (.A(_05653_),
    .ZN(_03667_));
 NAND2_X1 _17259_ (.A1(_02776_),
    .A2(_03667_),
    .ZN(_03668_));
 OAI21_X4 _17260_ (.A(_03668_),
    .B1(_05652_),
    .B2(_03470_),
    .ZN(_03669_));
 OAI22_X1 _17261_ (.A1(_02857_),
    .A2(_03666_),
    .B1(_03669_),
    .B2(_03025_),
    .ZN(_03670_));
 OR2_X1 _17262_ (.A1(_02991_),
    .A2(_05416_),
    .ZN(_03671_));
 OAI21_X4 _17263_ (.A(_03671_),
    .B1(_05417_),
    .B2(_02995_),
    .ZN(_03672_));
 OR2_X1 _17264_ (.A1(_05465_),
    .A2(_05584_),
    .ZN(_03673_));
 OAI21_X4 _17265_ (.A(_03673_),
    .B1(_05585_),
    .B2(_07525_),
    .ZN(_03674_));
 OAI22_X1 _17266_ (.A1(_03212_),
    .A2(_03672_),
    .B1(_03674_),
    .B2(_06960_),
    .ZN(_03675_));
 AND2_X1 _17267_ (.A1(_05737_),
    .A2(_06428_),
    .ZN(_03676_));
 AOI21_X4 _17268_ (.A(_03676_),
    .B1(_06283_),
    .B2(_02839_),
    .ZN(_03677_));
 NOR2_X1 _17269_ (.A1(_03545_),
    .A2(_03677_),
    .ZN(_03678_));
 NOR3_X1 _17270_ (.A1(_03670_),
    .A2(_03675_),
    .A3(_03678_),
    .ZN(_03679_));
 NOR2_X2 _17271_ (.A1(_03525_),
    .A2(_03679_),
    .ZN(net347));
 AND2_X1 _17272_ (.A1(_05153_),
    .A2(_05243_),
    .ZN(_03680_));
 AOI21_X4 _17273_ (.A(_03680_),
    .B1(_05244_),
    .B2(_07446_),
    .ZN(_03681_));
 OR2_X1 _17274_ (.A1(_03222_),
    .A2(_05580_),
    .ZN(_03682_));
 OAI21_X4 _17275_ (.A(_03682_),
    .B1(_05581_),
    .B2(_03227_),
    .ZN(_03683_));
 OAI22_X1 _17276_ (.A1(_02857_),
    .A2(_03681_),
    .B1(_03683_),
    .B2(_03394_),
    .ZN(_03684_));
 OR2_X1 _17277_ (.A1(_02991_),
    .A2(_05446_),
    .ZN(_03685_));
 OAI21_X4 _17278_ (.A(_03685_),
    .B1(_05447_),
    .B2(_02995_),
    .ZN(_03686_));
 INV_X1 _17279_ (.A(_05642_),
    .ZN(_03687_));
 NAND2_X1 _17280_ (.A1(_03233_),
    .A2(_03687_),
    .ZN(_03688_));
 OAI21_X4 _17281_ (.A(_03688_),
    .B1(_05641_),
    .B2(_02941_),
    .ZN(_03689_));
 OAI22_X1 _17282_ (.A1(_02869_),
    .A2(_03686_),
    .B1(_03689_),
    .B2(_03235_),
    .ZN(_03690_));
 OR2_X1 _17283_ (.A1(_05922_),
    .A2(_06322_),
    .ZN(_03691_));
 OAI21_X4 _17284_ (.A(_03691_),
    .B1(_06329_),
    .B2(_07337_),
    .ZN(_03692_));
 NOR2_X1 _17285_ (.A1(_03545_),
    .A2(_03692_),
    .ZN(_03693_));
 NOR3_X1 _17286_ (.A1(_03684_),
    .A2(_03690_),
    .A3(_03693_),
    .ZN(_03694_));
 NOR2_X2 _17287_ (.A1(_03525_),
    .A2(_03694_),
    .ZN(net348));
 OR2_X1 _17288_ (.A1(_07445_),
    .A2(_05253_),
    .ZN(_03695_));
 OAI21_X4 _17289_ (.A(_03695_),
    .B1(_05254_),
    .B2(_07439_),
    .ZN(_03696_));
 INV_X1 _17290_ (.A(_05665_),
    .ZN(_03697_));
 NAND2_X1 _17291_ (.A1(_02776_),
    .A2(_03697_),
    .ZN(_03698_));
 OAI21_X4 _17292_ (.A(_03698_),
    .B1(_05664_),
    .B2(_03470_),
    .ZN(_03699_));
 OAI22_X2 _17293_ (.A1(_02906_),
    .A2(_03696_),
    .B1(_03699_),
    .B2(_03025_),
    .ZN(_03700_));
 OR2_X1 _17294_ (.A1(_02991_),
    .A2(_05407_),
    .ZN(_03701_));
 OAI21_X4 _17295_ (.A(_03701_),
    .B1(_05409_),
    .B2(_02995_),
    .ZN(_03702_));
 OR2_X1 _17296_ (.A1(_05465_),
    .A2(_05558_),
    .ZN(_03703_));
 OAI21_X4 _17297_ (.A(_03703_),
    .B1(_05559_),
    .B2(_07525_),
    .ZN(_03704_));
 OAI22_X2 _17298_ (.A1(_02869_),
    .A2(_03702_),
    .B1(_03704_),
    .B2(_06960_),
    .ZN(_03705_));
 NAND2_X1 _17299_ (.A1(_05738_),
    .A2(_06268_),
    .ZN(_03706_));
 OAI21_X4 _17300_ (.A(_03706_),
    .B1(_06488_),
    .B2(_05738_),
    .ZN(_03707_));
 NOR2_X1 _17301_ (.A1(_03545_),
    .A2(_03707_),
    .ZN(_03708_));
 NOR3_X2 _17302_ (.A1(_03700_),
    .A2(_03705_),
    .A3(_03708_),
    .ZN(_03709_));
 NOR2_X4 _17303_ (.A1(_03525_),
    .A2(_03709_),
    .ZN(net349));
 BUF_X4 _17304_ (.A(_05163_),
    .Z(_03710_));
 OR2_X1 _17305_ (.A1(_02791_),
    .A2(_05420_),
    .ZN(_03711_));
 OAI21_X4 _17306_ (.A(_03711_),
    .B1(_05421_),
    .B2(_02797_),
    .ZN(_03712_));
 OR2_X1 _17307_ (.A1(_05465_),
    .A2(_05571_),
    .ZN(_03713_));
 OAI21_X2 _17308_ (.A(_03713_),
    .B1(_05572_),
    .B2(_07525_),
    .ZN(_03714_));
 OAI22_X1 _17309_ (.A1(_03212_),
    .A2(_03712_),
    .B1(_03714_),
    .B2(_03394_),
    .ZN(_03715_));
 AND2_X1 _17310_ (.A1(_05153_),
    .A2(_05210_),
    .ZN(_03716_));
 AOI21_X4 _17311_ (.A(_03716_),
    .B1(_05212_),
    .B2(_02863_),
    .ZN(_03717_));
 INV_X1 _17312_ (.A(_05687_),
    .ZN(_03718_));
 NAND2_X1 _17313_ (.A1(_07244_),
    .A2(_03718_),
    .ZN(_03719_));
 OAI21_X4 _17314_ (.A(_03719_),
    .B1(_05686_),
    .B2(_03233_),
    .ZN(_03720_));
 OAI22_X1 _17315_ (.A1(_02783_),
    .A2(_03717_),
    .B1(_03720_),
    .B2(_03235_),
    .ZN(_03721_));
 AND2_X1 _17316_ (.A1(_02838_),
    .A2(_06397_),
    .ZN(_03722_));
 AOI21_X4 _17317_ (.A(_03722_),
    .B1(_06477_),
    .B2(_05738_),
    .ZN(_03723_));
 NOR2_X1 _17318_ (.A1(_03545_),
    .A2(_03723_),
    .ZN(_03724_));
 NOR3_X1 _17319_ (.A1(_03715_),
    .A2(_03721_),
    .A3(_03724_),
    .ZN(_03725_));
 NOR2_X2 _17320_ (.A1(_03710_),
    .A2(_03725_),
    .ZN(net350));
 OR2_X1 _17321_ (.A1(_07519_),
    .A2(_05545_),
    .ZN(_03726_));
 OAI21_X4 _17322_ (.A(_03726_),
    .B1(_05546_),
    .B2(_07526_),
    .ZN(_03727_));
 INV_X1 _17323_ (.A(_05657_),
    .ZN(_03728_));
 NAND2_X1 _17324_ (.A1(_03470_),
    .A2(_03728_),
    .ZN(_03729_));
 OAI21_X4 _17325_ (.A(_03729_),
    .B1(_05656_),
    .B2(_03470_),
    .ZN(_03730_));
 OAI22_X1 _17326_ (.A1(_02761_),
    .A2(_03727_),
    .B1(_03730_),
    .B2(_02780_),
    .ZN(_03731_));
 OR2_X1 _17327_ (.A1(_07445_),
    .A2(_05205_),
    .ZN(_03732_));
 OAI21_X2 _17328_ (.A(_03732_),
    .B1(_05206_),
    .B2(_07439_),
    .ZN(_03733_));
 OR2_X1 _17329_ (.A1(_07493_),
    .A2(_05398_),
    .ZN(_03734_));
 OAI21_X4 _17330_ (.A(_03734_),
    .B1(_05399_),
    .B2(_07499_),
    .ZN(_03735_));
 OAI22_X1 _17331_ (.A1(_02857_),
    .A2(_03733_),
    .B1(_03735_),
    .B2(_02801_),
    .ZN(_03736_));
 NOR2_X1 _17332_ (.A1(_03731_),
    .A2(_03736_),
    .ZN(_03737_));
 NOR2_X4 _17333_ (.A1(_06340_),
    .A2(_06347_),
    .ZN(_03738_));
 NAND2_X1 _17334_ (.A1(_03376_),
    .A2(_03738_),
    .ZN(_03739_));
 AOI21_X4 _17335_ (.A(_05163_),
    .B1(_03737_),
    .B2(_03739_),
    .ZN(net351));
 OR2_X1 _17336_ (.A1(_07493_),
    .A2(_05442_),
    .ZN(_03740_));
 OAI21_X4 _17337_ (.A(_03740_),
    .B1(_05443_),
    .B2(_07499_),
    .ZN(_03741_));
 OR2_X1 _17338_ (.A1(_03222_),
    .A2(_05535_),
    .ZN(_03742_));
 OAI21_X4 _17339_ (.A(_03742_),
    .B1(_05537_),
    .B2(_03227_),
    .ZN(_03743_));
 OAI22_X1 _17340_ (.A1(_03212_),
    .A2(_03741_),
    .B1(_03743_),
    .B2(_03394_),
    .ZN(_03744_));
 AND2_X1 _17341_ (.A1(_05153_),
    .A2(_05232_),
    .ZN(_03745_));
 AOI21_X4 _17342_ (.A(_03745_),
    .B1(_05233_),
    .B2(_02863_),
    .ZN(_03746_));
 INV_X1 _17343_ (.A(_05670_),
    .ZN(_03747_));
 NAND2_X1 _17344_ (.A1(_03233_),
    .A2(_03747_),
    .ZN(_03748_));
 OAI21_X4 _17345_ (.A(_03748_),
    .B1(_05669_),
    .B2(_03233_),
    .ZN(_03749_));
 OAI22_X1 _17346_ (.A1(_02783_),
    .A2(_03746_),
    .B1(_03749_),
    .B2(_03235_),
    .ZN(_03750_));
 AND2_X1 _17347_ (.A1(_05737_),
    .A2(_06294_),
    .ZN(_03751_));
 AOI21_X4 _17348_ (.A(_03751_),
    .B1(_06304_),
    .B2(_02839_),
    .ZN(_03752_));
 NOR2_X1 _17349_ (.A1(_03545_),
    .A2(_03752_),
    .ZN(_03753_));
 NOR3_X1 _17350_ (.A1(_03744_),
    .A2(_03750_),
    .A3(_03753_),
    .ZN(_03754_));
 NOR2_X2 _17351_ (.A1(_03710_),
    .A2(_03754_),
    .ZN(net352));
 OR2_X1 _17352_ (.A1(_07445_),
    .A2(_05216_),
    .ZN(_03755_));
 OAI21_X4 _17353_ (.A(_03755_),
    .B1(_05217_),
    .B2(_07439_),
    .ZN(_03756_));
 INV_X1 _17354_ (.A(_05691_),
    .ZN(_03757_));
 NAND2_X1 _17355_ (.A1(_02776_),
    .A2(_03757_),
    .ZN(_03758_));
 OAI21_X4 _17356_ (.A(_03758_),
    .B1(_05690_),
    .B2(_03470_),
    .ZN(_03759_));
 OAI22_X1 _17357_ (.A1(_02906_),
    .A2(_03756_),
    .B1(_03759_),
    .B2(_03025_),
    .ZN(_03760_));
 OR2_X1 _17358_ (.A1(_02991_),
    .A2(_05394_),
    .ZN(_03761_));
 OAI21_X2 _17359_ (.A(_03761_),
    .B1(_05395_),
    .B2(_02995_),
    .ZN(_03762_));
 OR2_X1 _17360_ (.A1(_05465_),
    .A2(_05526_),
    .ZN(_03763_));
 OAI21_X4 _17361_ (.A(_03763_),
    .B1(_05527_),
    .B2(_07525_),
    .ZN(_03764_));
 OAI22_X1 _17362_ (.A1(_02869_),
    .A2(_03762_),
    .B1(_03764_),
    .B2(_06960_),
    .ZN(_03765_));
 OR2_X1 _17363_ (.A1(_02838_),
    .A2(_06436_),
    .ZN(_03766_));
 OAI21_X4 _17364_ (.A(_03766_),
    .B1(_06456_),
    .B2(_05738_),
    .ZN(_03767_));
 NOR2_X1 _17365_ (.A1(_03545_),
    .A2(_03767_),
    .ZN(_03768_));
 NOR3_X1 _17366_ (.A1(_03760_),
    .A2(_03765_),
    .A3(_03768_),
    .ZN(_03769_));
 NOR2_X2 _17367_ (.A1(_03710_),
    .A2(_03769_),
    .ZN(net353));
 OR2_X1 _17368_ (.A1(_07493_),
    .A2(_05390_),
    .ZN(_03770_));
 OAI21_X2 _17369_ (.A(_03770_),
    .B1(_05391_),
    .B2(_07499_),
    .ZN(_03771_));
 OR2_X1 _17370_ (.A1(_03222_),
    .A2(_05567_),
    .ZN(_03772_));
 OAI21_X4 _17371_ (.A(_03772_),
    .B1(_05568_),
    .B2(_03227_),
    .ZN(_03773_));
 OAI22_X1 _17372_ (.A1(_03212_),
    .A2(_03771_),
    .B1(_03773_),
    .B2(_03394_),
    .ZN(_03774_));
 AND2_X1 _17373_ (.A1(_05153_),
    .A2(_05227_),
    .ZN(_03775_));
 AOI21_X4 _17374_ (.A(_03775_),
    .B1(_05228_),
    .B2(_02863_),
    .ZN(_03776_));
 INV_X1 _17375_ (.A(_05674_),
    .ZN(_03777_));
 NAND2_X1 _17376_ (.A1(_03233_),
    .A2(_03777_),
    .ZN(_03778_));
 OAI21_X4 _17377_ (.A(_03778_),
    .B1(_05673_),
    .B2(_03233_),
    .ZN(_03779_));
 OAI22_X1 _17378_ (.A1(_02783_),
    .A2(_03776_),
    .B1(_03779_),
    .B2(_03235_),
    .ZN(_03780_));
 OR2_X1 _17379_ (.A1(_02838_),
    .A2(_06417_),
    .ZN(_03781_));
 OAI21_X4 _17380_ (.A(_03781_),
    .B1(_06387_),
    .B2(_05738_),
    .ZN(_03782_));
 NOR2_X1 _17381_ (.A1(_03545_),
    .A2(_03782_),
    .ZN(_03783_));
 NOR3_X1 _17382_ (.A1(_03774_),
    .A2(_03780_),
    .A3(_03783_),
    .ZN(_03784_));
 NOR2_X2 _17383_ (.A1(_03710_),
    .A2(_03784_),
    .ZN(net354));
 MUX2_X1 _17384_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][5] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][5] ),
    .S(_03223_),
    .Z(_03785_));
 OR2_X1 _17385_ (.A1(_03222_),
    .A2(_03785_),
    .ZN(_03786_));
 MUX2_X1 _17386_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][5] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][5] ),
    .S(_02938_),
    .Z(_03787_));
 OAI21_X4 _17387_ (.A(_03786_),
    .B1(_03787_),
    .B2(_03227_),
    .ZN(_03788_));
 MUX2_X1 _17388_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][5] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][5] ),
    .S(_03068_),
    .Z(_03789_));
 INV_X1 _17389_ (.A(_03789_),
    .ZN(_03790_));
 NAND2_X1 _17390_ (.A1(_02941_),
    .A2(_03790_),
    .ZN(_03791_));
 MUX2_X1 _17391_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][5] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][5] ),
    .S(_07246_),
    .Z(_03792_));
 OAI21_X4 _17392_ (.A(_03791_),
    .B1(_03792_),
    .B2(_02769_),
    .ZN(_03793_));
 OAI22_X1 _17393_ (.A1(_03015_),
    .A2(_03788_),
    .B1(_03793_),
    .B2(_03025_),
    .ZN(_03794_));
 MUX2_X1 _17394_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][5] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][5] ),
    .S(_02859_),
    .Z(_03795_));
 OR2_X1 _17395_ (.A1(_02858_),
    .A2(_03795_),
    .ZN(_03796_));
 MUX2_X1 _17396_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][5] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][5] ),
    .S(_02950_),
    .Z(_03797_));
 OAI21_X4 _17397_ (.A(_03796_),
    .B1(_03797_),
    .B2(_02789_),
    .ZN(_03798_));
 MUX2_X1 _17398_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][5] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][5] ),
    .S(_03184_),
    .Z(_03799_));
 OR2_X1 _17399_ (.A1(_07488_),
    .A2(_03799_),
    .ZN(_03800_));
 MUX2_X1 _17400_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][5] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][5] ),
    .S(_07494_),
    .Z(_03801_));
 OAI21_X4 _17401_ (.A(_03800_),
    .B1(_03801_),
    .B2(_07499_),
    .ZN(_03802_));
 OAI22_X1 _17402_ (.A1(_03066_),
    .A2(_03798_),
    .B1(_03802_),
    .B2(_03351_),
    .ZN(_03803_));
 MUX2_X1 _17403_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][5] ),
    .S(_02818_),
    .Z(_03804_));
 MUX2_X1 _17404_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][5] ),
    .S(_03191_),
    .Z(_03805_));
 MUX2_X1 _17405_ (.A(_03804_),
    .B(_03805_),
    .S(_03277_),
    .Z(_03806_));
 NAND2_X1 _17406_ (.A1(_07130_),
    .A2(_03806_),
    .ZN(_03807_));
 MUX2_X1 _17407_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][5] ),
    .S(_03280_),
    .Z(_03808_));
 MUX2_X1 _17408_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][5] ),
    .S(_03042_),
    .Z(_03809_));
 MUX2_X1 _17409_ (.A(_03808_),
    .B(_03809_),
    .S(_02834_),
    .Z(_03810_));
 NAND2_X1 _17410_ (.A1(_07391_),
    .A2(_03810_),
    .ZN(_03811_));
 NAND3_X2 _17411_ (.A1(_03036_),
    .A2(_03807_),
    .A3(_03811_),
    .ZN(_03812_));
 MUX2_X1 _17412_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][5] ),
    .S(_03047_),
    .Z(_03813_));
 MUX2_X1 _17413_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][5] ),
    .S(_02824_),
    .Z(_03814_));
 MUX2_X1 _17414_ (.A(_03813_),
    .B(_03814_),
    .S(_07336_),
    .Z(_03815_));
 MUX2_X1 _17415_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][5] ),
    .S(_03203_),
    .Z(_03816_));
 MUX2_X1 _17416_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][5] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][5] ),
    .S(_02830_),
    .Z(_03817_));
 MUX2_X1 _17417_ (.A(_03816_),
    .B(_03817_),
    .S(_03206_),
    .Z(_03818_));
 MUX2_X1 _17418_ (.A(_03815_),
    .B(_03818_),
    .S(_03292_),
    .Z(_03819_));
 OAI21_X4 _17419_ (.A(_03812_),
    .B1(_03819_),
    .B2(_02805_),
    .ZN(_03820_));
 NOR2_X1 _17420_ (.A1(_03545_),
    .A2(_03820_),
    .ZN(_03821_));
 NOR3_X1 _17421_ (.A1(_03794_),
    .A2(_03803_),
    .A3(_03821_),
    .ZN(_03822_));
 NOR2_X2 _17422_ (.A1(_03710_),
    .A2(_03822_),
    .ZN(net355));
 NAND2_X1 _17423_ (.A1(_02857_),
    .A2(_05160_),
    .ZN(_03823_));
 AOI22_X1 _17424_ (.A1(_03379_),
    .A2(_05427_),
    .B1(_05556_),
    .B2(_06996_),
    .ZN(_03824_));
 AOI22_X1 _17425_ (.A1(_03380_),
    .A2(_05194_),
    .B1(_05639_),
    .B2(_03372_),
    .ZN(_03825_));
 MUX2_X1 _17426_ (.A(_06307_),
    .B(_06466_),
    .S(_05737_),
    .Z(_03826_));
 MUX2_X2 _17427_ (.A(_06258_),
    .B(_03826_),
    .S(_02815_),
    .Z(_03827_));
 NAND2_X1 _17428_ (.A1(_02873_),
    .A2(_03827_),
    .ZN(_03828_));
 NAND3_X1 _17429_ (.A1(_03824_),
    .A2(_03825_),
    .A3(_03828_),
    .ZN(_03829_));
 AND2_X1 _17430_ (.A1(_03823_),
    .A2(_03829_),
    .ZN(net356));
 AND2_X1 _17431_ (.A1(_05153_),
    .A2(_05237_),
    .ZN(_03830_));
 AOI21_X4 _17432_ (.A(_03830_),
    .B1(_05238_),
    .B2(_02863_),
    .ZN(_03831_));
 OR2_X1 _17433_ (.A1(_03222_),
    .A2(_05563_),
    .ZN(_03832_));
 OAI21_X4 _17434_ (.A(_03832_),
    .B1(_05564_),
    .B2(_03227_),
    .ZN(_03833_));
 OAI22_X1 _17435_ (.A1(_02906_),
    .A2(_03831_),
    .B1(_03833_),
    .B2(_03394_),
    .ZN(_03834_));
 OR2_X1 _17436_ (.A1(_02791_),
    .A2(_05437_),
    .ZN(_03835_));
 OAI21_X2 _17437_ (.A(_03835_),
    .B1(_05438_),
    .B2(_02797_),
    .ZN(_03836_));
 INV_X1 _17438_ (.A(_05678_),
    .ZN(_03837_));
 NAND2_X1 _17439_ (.A1(_07244_),
    .A2(_03837_),
    .ZN(_03838_));
 OAI21_X4 _17440_ (.A(_03838_),
    .B1(_05677_),
    .B2(_03233_),
    .ZN(_03839_));
 OAI22_X1 _17441_ (.A1(_02869_),
    .A2(_03836_),
    .B1(_03839_),
    .B2(_03235_),
    .ZN(_03840_));
 MUX2_X1 _17442_ (.A(_06370_),
    .B(_06374_),
    .S(_05946_),
    .Z(_03841_));
 NAND2_X1 _17443_ (.A1(_02838_),
    .A2(_03841_),
    .ZN(_03842_));
 MUX2_X1 _17444_ (.A(_06400_),
    .B(_06404_),
    .S(_05946_),
    .Z(_03843_));
 NAND2_X1 _17445_ (.A1(_05737_),
    .A2(_03843_),
    .ZN(_03844_));
 NAND3_X1 _17446_ (.A1(_05922_),
    .A2(_03842_),
    .A3(_03844_),
    .ZN(_03845_));
 MUX2_X1 _17447_ (.A(_06372_),
    .B(_06375_),
    .S(_07384_),
    .Z(_03846_));
 MUX2_X1 _17448_ (.A(_06402_),
    .B(_06405_),
    .S(_07384_),
    .Z(_03847_));
 MUX2_X1 _17449_ (.A(_03846_),
    .B(_03847_),
    .S(_05737_),
    .Z(_03848_));
 OAI21_X4 _17450_ (.A(_03845_),
    .B1(_03848_),
    .B2(_05922_),
    .ZN(_03849_));
 NOR2_X1 _17451_ (.A1(_02803_),
    .A2(_03849_),
    .ZN(_03850_));
 NOR3_X1 _17452_ (.A1(_03834_),
    .A2(_03840_),
    .A3(_03850_),
    .ZN(_03851_));
 NOR2_X2 _17453_ (.A1(_03710_),
    .A2(_03851_),
    .ZN(net357));
 AND2_X1 _17454_ (.A1(_02784_),
    .A2(_05198_),
    .ZN(_03852_));
 AOI21_X4 _17455_ (.A(_03852_),
    .B1(_05199_),
    .B2(_07446_),
    .ZN(_03853_));
 OR2_X1 _17456_ (.A1(_07493_),
    .A2(_05433_),
    .ZN(_03854_));
 OAI21_X4 _17457_ (.A(_03854_),
    .B1(_05434_),
    .B2(_07499_),
    .ZN(_03855_));
 OAI22_X1 _17458_ (.A1(_02857_),
    .A2(_03853_),
    .B1(_03855_),
    .B2(_03212_),
    .ZN(_03856_));
 OR2_X1 _17459_ (.A1(_07519_),
    .A2(_05540_),
    .ZN(_03857_));
 OAI21_X4 _17460_ (.A(_03857_),
    .B1(_05541_),
    .B2(_07526_),
    .ZN(_03858_));
 INV_X1 _17461_ (.A(_05661_),
    .ZN(_03859_));
 NAND2_X1 _17462_ (.A1(_02776_),
    .A2(_03859_),
    .ZN(_03860_));
 OAI21_X4 _17463_ (.A(_03860_),
    .B1(_05660_),
    .B2(_03470_),
    .ZN(_03861_));
 OAI22_X1 _17464_ (.A1(_02761_),
    .A2(_03858_),
    .B1(_03861_),
    .B2(_02780_),
    .ZN(_03862_));
 NOR2_X1 _17465_ (.A1(_03856_),
    .A2(_03862_),
    .ZN(_03863_));
 NOR2_X4 _17466_ (.A1(_06357_),
    .A2(_06365_),
    .ZN(_03864_));
 NAND2_X1 _17467_ (.A1(_03376_),
    .A2(_03864_),
    .ZN(_03865_));
 AOI21_X2 _17468_ (.A(_05163_),
    .B1(_03863_),
    .B2(_03865_),
    .ZN(net358));
 OR2_X1 _17469_ (.A1(_07445_),
    .A2(_05222_),
    .ZN(_03866_));
 OAI21_X4 _17470_ (.A(_03866_),
    .B1(_05223_),
    .B2(_07439_),
    .ZN(_03867_));
 OR2_X1 _17471_ (.A1(_05465_),
    .A2(_05575_),
    .ZN(_03868_));
 OAI21_X2 _17472_ (.A(_03868_),
    .B1(_05576_),
    .B2(_07525_),
    .ZN(_03869_));
 OAI22_X1 _17473_ (.A1(_02906_),
    .A2(_03867_),
    .B1(_03869_),
    .B2(_06960_),
    .ZN(_03870_));
 OR2_X1 _17474_ (.A1(_02991_),
    .A2(_05402_),
    .ZN(_03871_));
 OAI21_X2 _17475_ (.A(_03871_),
    .B1(_05403_),
    .B2(_02995_),
    .ZN(_03872_));
 INV_X1 _17476_ (.A(_05634_),
    .ZN(_03873_));
 NAND2_X1 _17477_ (.A1(_03233_),
    .A2(_03873_),
    .ZN(_03874_));
 OAI21_X4 _17478_ (.A(_03874_),
    .B1(_05633_),
    .B2(_02941_),
    .ZN(_03875_));
 OAI22_X1 _17479_ (.A1(_02869_),
    .A2(_03872_),
    .B1(_03875_),
    .B2(_03235_),
    .ZN(_03876_));
 NOR2_X1 _17480_ (.A1(_02803_),
    .A2(_06229_),
    .ZN(_03877_));
 NOR3_X1 _17481_ (.A1(_03870_),
    .A2(_03876_),
    .A3(_03877_),
    .ZN(_03878_));
 NOR2_X2 _17482_ (.A1(_03710_),
    .A2(_03878_),
    .ZN(net359));
 MUX2_X1 _17483_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][6] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][6] ),
    .S(_03223_),
    .Z(_03879_));
 OR2_X1 _17484_ (.A1(_03222_),
    .A2(_03879_),
    .ZN(_03880_));
 MUX2_X1 _17485_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][6] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][6] ),
    .S(_02938_),
    .Z(_03881_));
 OAI21_X4 _17486_ (.A(_03880_),
    .B1(_03881_),
    .B2(_03227_),
    .ZN(_03882_));
 MUX2_X1 _17487_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][6] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][6] ),
    .S(_03068_),
    .Z(_03883_));
 INV_X1 _17488_ (.A(_03883_),
    .ZN(_03884_));
 NAND2_X1 _17489_ (.A1(_02941_),
    .A2(_03884_),
    .ZN(_03885_));
 MUX2_X1 _17490_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][6] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][6] ),
    .S(_02774_),
    .Z(_03886_));
 OAI21_X4 _17491_ (.A(_03885_),
    .B1(_03886_),
    .B2(_02769_),
    .ZN(_03887_));
 OAI22_X1 _17492_ (.A1(_03015_),
    .A2(_03882_),
    .B1(_03887_),
    .B2(_03235_),
    .ZN(_03888_));
 MUX2_X1 _17493_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][6] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][6] ),
    .S(_02785_),
    .Z(_03889_));
 OR2_X1 _17494_ (.A1(_02784_),
    .A2(_03889_),
    .ZN(_03890_));
 MUX2_X1 _17495_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][6] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][6] ),
    .S(_02950_),
    .Z(_03891_));
 OAI21_X4 _17496_ (.A(_03890_),
    .B1(_03891_),
    .B2(_02789_),
    .ZN(_03892_));
 MUX2_X1 _17497_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][6] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][6] ),
    .S(_03184_),
    .Z(_03893_));
 OR2_X1 _17498_ (.A1(_07488_),
    .A2(_03893_),
    .ZN(_03894_));
 MUX2_X1 _17499_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][6] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][6] ),
    .S(_07494_),
    .Z(_03895_));
 OAI21_X4 _17500_ (.A(_03894_),
    .B1(_03895_),
    .B2(_07499_),
    .ZN(_03896_));
 OAI22_X1 _17501_ (.A1(_03066_),
    .A2(_03892_),
    .B1(_03896_),
    .B2(_03351_),
    .ZN(_03897_));
 MUX2_X1 _17502_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][6] ),
    .S(_02818_),
    .Z(_03898_));
 MUX2_X1 _17503_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][6] ),
    .S(_03191_),
    .Z(_03899_));
 MUX2_X1 _17504_ (.A(_03898_),
    .B(_03899_),
    .S(_03277_),
    .Z(_03900_));
 NAND2_X1 _17505_ (.A1(_07130_),
    .A2(_03900_),
    .ZN(_03901_));
 MUX2_X1 _17506_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][6] ),
    .S(_03280_),
    .Z(_03902_));
 MUX2_X1 _17507_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][6] ),
    .S(_02816_),
    .Z(_03903_));
 MUX2_X1 _17508_ (.A(_03902_),
    .B(_03903_),
    .S(_02834_),
    .Z(_03904_));
 NAND2_X1 _17509_ (.A1(_07391_),
    .A2(_03904_),
    .ZN(_03905_));
 NAND3_X2 _17510_ (.A1(_02838_),
    .A2(_03901_),
    .A3(_03905_),
    .ZN(_03906_));
 MUX2_X1 _17511_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][6] ),
    .S(_07325_),
    .Z(_03907_));
 MUX2_X1 _17512_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][6] ),
    .S(_02824_),
    .Z(_03908_));
 MUX2_X1 _17513_ (.A(_03907_),
    .B(_03908_),
    .S(_07336_),
    .Z(_03909_));
 MUX2_X1 _17514_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][6] ),
    .S(_03203_),
    .Z(_03910_));
 MUX2_X1 _17515_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][6] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][6] ),
    .S(_02830_),
    .Z(_03911_));
 MUX2_X1 _17516_ (.A(_03910_),
    .B(_03911_),
    .S(_03206_),
    .Z(_03912_));
 MUX2_X1 _17517_ (.A(_03909_),
    .B(_03912_),
    .S(_03292_),
    .Z(_03913_));
 OAI21_X4 _17518_ (.A(_03906_),
    .B1(_03913_),
    .B2(_02805_),
    .ZN(_03914_));
 NOR2_X1 _17519_ (.A1(_02803_),
    .A2(_03914_),
    .ZN(_03915_));
 NOR3_X1 _17520_ (.A1(_03888_),
    .A2(_03897_),
    .A3(_03915_),
    .ZN(_03916_));
 NOR2_X2 _17521_ (.A1(_03710_),
    .A2(_03916_),
    .ZN(net360));
 MUX2_X1 _17522_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][7] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][7] ),
    .S(_03223_),
    .Z(_03917_));
 OR2_X1 _17523_ (.A1(_03222_),
    .A2(_03917_),
    .ZN(_03918_));
 MUX2_X1 _17524_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][7] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][7] ),
    .S(_07520_),
    .Z(_03919_));
 OAI21_X4 _17525_ (.A(_03918_),
    .B1(_03919_),
    .B2(_03227_),
    .ZN(_03920_));
 MUX2_X1 _17526_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][7] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][7] ),
    .S(_03068_),
    .Z(_03921_));
 INV_X1 _17527_ (.A(_03921_),
    .ZN(_03922_));
 NAND2_X1 _17528_ (.A1(_02941_),
    .A2(_03922_),
    .ZN(_03923_));
 MUX2_X1 _17529_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][7] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][7] ),
    .S(_02774_),
    .Z(_03924_));
 OAI21_X4 _17530_ (.A(_03923_),
    .B1(_03924_),
    .B2(_02776_),
    .ZN(_03925_));
 OAI22_X1 _17531_ (.A1(_03015_),
    .A2(_03920_),
    .B1(_03925_),
    .B2(_03235_),
    .ZN(_03926_));
 MUX2_X1 _17532_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][7] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][7] ),
    .S(_02785_),
    .Z(_03927_));
 OR2_X1 _17533_ (.A1(_02784_),
    .A2(_03927_),
    .ZN(_03928_));
 MUX2_X1 _17534_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][7] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][7] ),
    .S(_07440_),
    .Z(_03929_));
 OAI21_X4 _17535_ (.A(_03928_),
    .B1(_03929_),
    .B2(_07445_),
    .ZN(_03930_));
 MUX2_X1 _17536_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][7] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][7] ),
    .S(_03184_),
    .Z(_03931_));
 OR2_X1 _17537_ (.A1(_07488_),
    .A2(_03931_),
    .ZN(_03932_));
 MUX2_X1 _17538_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][7] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][7] ),
    .S(_07494_),
    .Z(_03933_));
 OAI21_X4 _17539_ (.A(_03932_),
    .B1(_03933_),
    .B2(_07499_),
    .ZN(_03934_));
 OAI22_X1 _17540_ (.A1(_03066_),
    .A2(_03930_),
    .B1(_03934_),
    .B2(_03351_),
    .ZN(_03935_));
 MUX2_X1 _17541_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][7] ),
    .S(_02818_),
    .Z(_03936_));
 MUX2_X1 _17542_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][7] ),
    .S(_03191_),
    .Z(_03937_));
 MUX2_X1 _17543_ (.A(_03936_),
    .B(_03937_),
    .S(_03277_),
    .Z(_03938_));
 NAND2_X1 _17544_ (.A1(_07130_),
    .A2(_03938_),
    .ZN(_03939_));
 MUX2_X1 _17545_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][7] ),
    .S(_03280_),
    .Z(_03940_));
 MUX2_X1 _17546_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][7] ),
    .S(_02816_),
    .Z(_03941_));
 MUX2_X1 _17547_ (.A(_03940_),
    .B(_03941_),
    .S(_02834_),
    .Z(_03942_));
 NAND2_X1 _17548_ (.A1(_07391_),
    .A2(_03942_),
    .ZN(_03943_));
 NAND3_X2 _17549_ (.A1(_02838_),
    .A2(_03939_),
    .A3(_03943_),
    .ZN(_03944_));
 MUX2_X1 _17550_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][7] ),
    .S(_07325_),
    .Z(_03945_));
 MUX2_X1 _17551_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][7] ),
    .S(_02824_),
    .Z(_03946_));
 MUX2_X1 _17552_ (.A(_03945_),
    .B(_03946_),
    .S(_07336_),
    .Z(_03947_));
 MUX2_X1 _17553_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][7] ),
    .S(_03203_),
    .Z(_03948_));
 MUX2_X1 _17554_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][7] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][7] ),
    .S(_02830_),
    .Z(_03949_));
 MUX2_X1 _17555_ (.A(_03948_),
    .B(_03949_),
    .S(_03206_),
    .Z(_03950_));
 MUX2_X1 _17556_ (.A(_03947_),
    .B(_03950_),
    .S(_03292_),
    .Z(_03951_));
 OAI21_X4 _17557_ (.A(_03944_),
    .B1(_03951_),
    .B2(_02805_),
    .ZN(_03952_));
 NOR2_X1 _17558_ (.A1(_02803_),
    .A2(_03952_),
    .ZN(_03953_));
 NOR3_X1 _17559_ (.A1(_03926_),
    .A2(_03935_),
    .A3(_03953_),
    .ZN(_03954_));
 NOR2_X2 _17560_ (.A1(_03710_),
    .A2(_03954_),
    .ZN(net361));
 MUX2_X1 _17561_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][8] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][8] ),
    .S(_07494_),
    .Z(_03955_));
 OR2_X1 _17562_ (.A1(_07493_),
    .A2(_03955_),
    .ZN(_03956_));
 MUX2_X1 _17563_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][8] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][8] ),
    .S(_07497_),
    .Z(_03957_));
 OAI21_X4 _17564_ (.A(_03956_),
    .B1(_03957_),
    .B2(_07499_),
    .ZN(_03958_));
 MUX2_X1 _17565_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][8] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][8] ),
    .S(_02785_),
    .Z(_03959_));
 OR2_X1 _17566_ (.A1(_02784_),
    .A2(_03959_),
    .ZN(_03960_));
 MUX2_X1 _17567_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][8] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][8] ),
    .S(_02950_),
    .Z(_03961_));
 OAI21_X4 _17568_ (.A(_03960_),
    .B1(_03961_),
    .B2(_02789_),
    .ZN(_03962_));
 OAI22_X1 _17569_ (.A1(_03212_),
    .A2(_03958_),
    .B1(_03962_),
    .B2(_02782_),
    .ZN(_03963_));
 MUX2_X1 _17570_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][8] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][8] ),
    .S(_03223_),
    .Z(_03964_));
 OR2_X1 _17571_ (.A1(_03222_),
    .A2(_03964_),
    .ZN(_03965_));
 MUX2_X1 _17572_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][8] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][8] ),
    .S(_07520_),
    .Z(_03966_));
 OAI21_X4 _17573_ (.A(_03965_),
    .B1(_03966_),
    .B2(_03227_),
    .ZN(_03967_));
 MUX2_X1 _17574_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][8] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][8] ),
    .S(_03068_),
    .Z(_03968_));
 INV_X1 _17575_ (.A(_03968_),
    .ZN(_03969_));
 NAND2_X1 _17576_ (.A1(_07244_),
    .A2(_03969_),
    .ZN(_03970_));
 MUX2_X1 _17577_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][8] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][8] ),
    .S(_07246_),
    .Z(_03971_));
 OAI21_X4 _17578_ (.A(_03970_),
    .B1(_03971_),
    .B2(_03233_),
    .ZN(_03972_));
 OAI22_X1 _17579_ (.A1(_02855_),
    .A2(_03967_),
    .B1(_03972_),
    .B2(_03235_),
    .ZN(_03973_));
 MUX2_X1 _17580_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][8] ),
    .S(_02818_),
    .Z(_03974_));
 MUX2_X1 _17581_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][8] ),
    .S(_02808_),
    .Z(_03975_));
 MUX2_X1 _17582_ (.A(_03974_),
    .B(_03975_),
    .S(_03277_),
    .Z(_03976_));
 NAND2_X1 _17583_ (.A1(_07130_),
    .A2(_03976_),
    .ZN(_03977_));
 MUX2_X1 _17584_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][8] ),
    .S(_03280_),
    .Z(_03978_));
 MUX2_X1 _17585_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][8] ),
    .S(_02816_),
    .Z(_03979_));
 MUX2_X1 _17586_ (.A(_03978_),
    .B(_03979_),
    .S(_02834_),
    .Z(_03980_));
 NAND2_X1 _17587_ (.A1(_07391_),
    .A2(_03980_),
    .ZN(_03981_));
 NAND3_X2 _17588_ (.A1(_02838_),
    .A2(_03977_),
    .A3(_03981_),
    .ZN(_03982_));
 MUX2_X1 _17589_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][8] ),
    .S(_07325_),
    .Z(_03983_));
 MUX2_X1 _17590_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][8] ),
    .S(_02824_),
    .Z(_03984_));
 MUX2_X1 _17591_ (.A(_03983_),
    .B(_03984_),
    .S(_07336_),
    .Z(_03985_));
 MUX2_X1 _17592_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][8] ),
    .S(_02826_),
    .Z(_03986_));
 MUX2_X1 _17593_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][8] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][8] ),
    .S(_02830_),
    .Z(_03987_));
 MUX2_X1 _17594_ (.A(_03986_),
    .B(_03987_),
    .S(_02828_),
    .Z(_03988_));
 MUX2_X1 _17595_ (.A(_03985_),
    .B(_03988_),
    .S(_03292_),
    .Z(_03989_));
 OAI21_X4 _17596_ (.A(_03982_),
    .B1(_03989_),
    .B2(_02805_),
    .ZN(_03990_));
 NOR2_X1 _17597_ (.A1(_02803_),
    .A2(_03990_),
    .ZN(_03991_));
 NOR3_X1 _17598_ (.A1(_03963_),
    .A2(_03973_),
    .A3(_03991_),
    .ZN(_03992_));
 NOR2_X2 _17599_ (.A1(_03710_),
    .A2(_03992_),
    .ZN(net362));
 MUX2_X1 _17600_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[1][9] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[3][9] ),
    .S(_02770_),
    .Z(_03993_));
 INV_X1 _17601_ (.A(_03993_),
    .ZN(_03994_));
 NAND2_X1 _17602_ (.A1(_03470_),
    .A2(_03994_),
    .ZN(_03995_));
 MUX2_X1 _17603_ (.A(\dynamic_node_top.south_input.NIB.storage_data_f[0][9] ),
    .B(\dynamic_node_top.south_input.NIB.storage_data_f[2][9] ),
    .S(_02774_),
    .Z(_03996_));
 OAI21_X4 _17604_ (.A(_03995_),
    .B1(_03996_),
    .B2(_02845_),
    .ZN(_03997_));
 MUX2_X1 _17605_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[0][9] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[2][9] ),
    .S(_02859_),
    .Z(_03998_));
 OR2_X1 _17606_ (.A1(_02858_),
    .A2(_03998_),
    .ZN(_03999_));
 MUX2_X1 _17607_ (.A(\dynamic_node_top.west_input.NIB.storage_data_f[1][9] ),
    .B(\dynamic_node_top.west_input.NIB.storage_data_f[3][9] ),
    .S(_02950_),
    .Z(_04000_));
 OAI21_X4 _17608_ (.A(_03999_),
    .B1(_04000_),
    .B2(_02863_),
    .ZN(_04001_));
 OAI22_X1 _17609_ (.A1(_02780_),
    .A2(_03997_),
    .B1(_04001_),
    .B2(_02782_),
    .ZN(_04002_));
 MUX2_X1 _17610_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[0][9] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[2][9] ),
    .S(_03223_),
    .Z(_04003_));
 OR2_X1 _17611_ (.A1(_05465_),
    .A2(_04003_),
    .ZN(_04004_));
 MUX2_X1 _17612_ (.A(\dynamic_node_top.east_input.NIB.storage_data_f[1][9] ),
    .B(\dynamic_node_top.east_input.NIB.storage_data_f[3][9] ),
    .S(_07520_),
    .Z(_04005_));
 OAI21_X4 _17613_ (.A(_04004_),
    .B1(_04005_),
    .B2(_07525_),
    .ZN(_04006_));
 MUX2_X1 _17614_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[0][9] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[2][9] ),
    .S(_03184_),
    .Z(_04007_));
 OR2_X1 _17615_ (.A1(_07488_),
    .A2(_04007_),
    .ZN(_04008_));
 MUX2_X1 _17616_ (.A(\dynamic_node_top.north_input.NIB.storage_data_f[1][9] ),
    .B(\dynamic_node_top.north_input.NIB.storage_data_f[3][9] ),
    .S(_07494_),
    .Z(_04009_));
 OAI21_X4 _17617_ (.A(_04008_),
    .B1(_04009_),
    .B2(_07499_),
    .ZN(_04010_));
 OAI22_X1 _17618_ (.A1(_02855_),
    .A2(_04006_),
    .B1(_04010_),
    .B2(_03351_),
    .ZN(_04011_));
 MUX2_X1 _17619_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[8][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[10][9] ),
    .S(_02818_),
    .Z(_04012_));
 MUX2_X1 _17620_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[9][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[11][9] ),
    .S(_02808_),
    .Z(_04013_));
 MUX2_X1 _17621_ (.A(_04012_),
    .B(_04013_),
    .S(_03277_),
    .Z(_04014_));
 NAND2_X1 _17622_ (.A1(_07130_),
    .A2(_04014_),
    .ZN(_04015_));
 MUX2_X1 _17623_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[0][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[2][9] ),
    .S(_03280_),
    .Z(_04016_));
 MUX2_X1 _17624_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[1][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[3][9] ),
    .S(_02816_),
    .Z(_04017_));
 MUX2_X1 _17625_ (.A(_04016_),
    .B(_04017_),
    .S(_02834_),
    .Z(_04018_));
 NAND2_X1 _17626_ (.A1(_07391_),
    .A2(_04018_),
    .ZN(_04019_));
 NAND3_X2 _17627_ (.A1(_02838_),
    .A2(_04015_),
    .A3(_04019_),
    .ZN(_04020_));
 MUX2_X1 _17628_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[12][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[14][9] ),
    .S(_07325_),
    .Z(_04021_));
 MUX2_X1 _17629_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[13][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[15][9] ),
    .S(_02824_),
    .Z(_04022_));
 MUX2_X1 _17630_ (.A(_04021_),
    .B(_04022_),
    .S(_07336_),
    .Z(_04023_));
 MUX2_X1 _17631_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[4][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[6][9] ),
    .S(_02826_),
    .Z(_04024_));
 MUX2_X1 _17632_ (.A(\dynamic_node_top.proc_input.NIB.storage_data_f[5][9] ),
    .B(\dynamic_node_top.proc_input.NIB.storage_data_f[7][9] ),
    .S(_02830_),
    .Z(_04025_));
 MUX2_X1 _17633_ (.A(_04024_),
    .B(_04025_),
    .S(_02828_),
    .Z(_04026_));
 MUX2_X1 _17634_ (.A(_04023_),
    .B(_04026_),
    .S(_03292_),
    .Z(_04027_));
 OAI21_X4 _17635_ (.A(_04020_),
    .B1(_04027_),
    .B2(_02805_),
    .ZN(_04028_));
 NOR2_X1 _17636_ (.A1(_02803_),
    .A2(_04028_),
    .ZN(_04029_));
 NOR3_X1 _17637_ (.A1(_04002_),
    .A2(_04011_),
    .A3(_04029_),
    .ZN(_04030_));
 NOR2_X2 _17638_ (.A1(_02843_),
    .A2(_04030_),
    .ZN(net363));
 BUF_X4 _17639_ (.A(_06086_),
    .Z(_04031_));
 BUF_X4 _17640_ (.A(_04031_),
    .Z(_04032_));
 CLKBUF_X3 _17641_ (.A(_00071_),
    .Z(_04033_));
 BUF_X4 _17642_ (.A(_04033_),
    .Z(_04034_));
 BUF_X4 _17643_ (.A(_04034_),
    .Z(_04035_));
 BUF_X4 _17644_ (.A(_06085_),
    .Z(_04036_));
 OAI22_X1 _17645_ (.A1(_04035_),
    .A2(_02768_),
    .B1(_02777_),
    .B2(_04036_),
    .ZN(_04037_));
 BUF_X4 _17646_ (.A(_00073_),
    .Z(_04038_));
 BUF_X4 _17647_ (.A(_04038_),
    .Z(_04039_));
 BUF_X4 _17648_ (.A(_07022_),
    .Z(_04040_));
 CLKBUF_X3 _17649_ (.A(_04040_),
    .Z(_04041_));
 OAI22_X1 _17650_ (.A1(_04039_),
    .A2(_02790_),
    .B1(_02798_),
    .B2(_04041_),
    .ZN(_04042_));
 BUF_X4 _17651_ (.A(_00072_),
    .Z(_04043_));
 CLKBUF_X3 _17652_ (.A(_04043_),
    .Z(_04044_));
 NOR2_X1 _17653_ (.A1(_04044_),
    .A2(_02840_),
    .ZN(_04045_));
 NOR3_X1 _17654_ (.A1(_04037_),
    .A2(_04042_),
    .A3(_04045_),
    .ZN(_04046_));
 NOR2_X2 _17655_ (.A1(_04032_),
    .A2(_04046_),
    .ZN(net364));
 BUF_X4 _17656_ (.A(_04031_),
    .Z(_04047_));
 BUF_X4 _17657_ (.A(_04038_),
    .Z(_04048_));
 BUF_X4 _17658_ (.A(_04048_),
    .Z(_04049_));
 OAI22_X1 _17659_ (.A1(_04035_),
    .A2(_02854_),
    .B1(_02864_),
    .B2(_04049_),
    .ZN(_04050_));
 BUF_X4 _17660_ (.A(_06085_),
    .Z(_04051_));
 BUF_X4 _17661_ (.A(_04040_),
    .Z(_04052_));
 OAI22_X1 _17662_ (.A1(_04051_),
    .A2(_02850_),
    .B1(_02868_),
    .B2(_04052_),
    .ZN(_04053_));
 NOR2_X1 _17663_ (.A1(_04050_),
    .A2(_04053_),
    .ZN(_04054_));
 INV_X1 _17664_ (.A(_04043_),
    .ZN(_04055_));
 BUF_X4 _17665_ (.A(_04055_),
    .Z(_04056_));
 BUF_X4 _17666_ (.A(_04056_),
    .Z(_04057_));
 NAND2_X1 _17667_ (.A1(_04057_),
    .A2(_02896_),
    .ZN(_04058_));
 AOI21_X2 _17668_ (.A(_04047_),
    .B1(_04054_),
    .B2(_04058_),
    .ZN(net365));
 BUF_X4 _17669_ (.A(_04048_),
    .Z(_04059_));
 BUF_X4 _17670_ (.A(_06085_),
    .Z(_04060_));
 OAI22_X2 _17671_ (.A1(_04059_),
    .A2(_02905_),
    .B1(_02912_),
    .B2(_04060_),
    .ZN(_04061_));
 OAI22_X2 _17672_ (.A1(_04035_),
    .A2(_02901_),
    .B1(_02916_),
    .B2(_04052_),
    .ZN(_04062_));
 NOR2_X2 _17673_ (.A1(_04061_),
    .A2(_04062_),
    .ZN(_04063_));
 NAND2_X1 _17674_ (.A1(_04057_),
    .A2(_02934_),
    .ZN(_04064_));
 AOI21_X4 _17675_ (.A(_04047_),
    .B1(_04063_),
    .B2(_04064_),
    .ZN(net366));
 CLKBUF_X3 _17676_ (.A(_04034_),
    .Z(_04065_));
 OAI22_X1 _17677_ (.A1(_04065_),
    .A2(_02940_),
    .B1(_02946_),
    .B2(_04036_),
    .ZN(_04066_));
 OAI22_X1 _17678_ (.A1(_04039_),
    .A2(_02952_),
    .B1(_02956_),
    .B2(_04041_),
    .ZN(_04067_));
 NOR2_X1 _17679_ (.A1(_04044_),
    .A2(_02974_),
    .ZN(_04068_));
 NOR3_X1 _17680_ (.A1(_04066_),
    .A2(_04067_),
    .A3(_04068_),
    .ZN(_04069_));
 NOR2_X2 _17681_ (.A1(_04032_),
    .A2(_04069_),
    .ZN(net367));
 OAI22_X1 _17682_ (.A1(_04035_),
    .A2(_02985_),
    .B1(_02990_),
    .B2(_04049_),
    .ZN(_04070_));
 OAI22_X1 _17683_ (.A1(_04051_),
    .A2(_02981_),
    .B1(_02996_),
    .B2(_04052_),
    .ZN(_04071_));
 NOR2_X1 _17684_ (.A1(_04070_),
    .A2(_04071_),
    .ZN(_04072_));
 NAND2_X1 _17685_ (.A1(_04057_),
    .A2(_03013_),
    .ZN(_04073_));
 AOI21_X2 _17686_ (.A(_04047_),
    .B1(_04072_),
    .B2(_04073_),
    .ZN(net368));
 OAI22_X1 _17687_ (.A1(_04065_),
    .A2(_03019_),
    .B1(_03024_),
    .B2(_04036_),
    .ZN(_04074_));
 OAI22_X1 _17688_ (.A1(_04039_),
    .A2(_03030_),
    .B1(_03034_),
    .B2(_04041_),
    .ZN(_04075_));
 NOR2_X1 _17689_ (.A1(_04044_),
    .A2(_03055_),
    .ZN(_04076_));
 NOR3_X1 _17690_ (.A1(_04074_),
    .A2(_04075_),
    .A3(_04076_),
    .ZN(_04077_));
 NOR2_X2 _17691_ (.A1(_04032_),
    .A2(_04077_),
    .ZN(net369));
 BUF_X4 _17692_ (.A(_04038_),
    .Z(_04078_));
 OAI22_X1 _17693_ (.A1(_04065_),
    .A2(_03061_),
    .B1(_03065_),
    .B2(_04078_),
    .ZN(_04079_));
 OAI22_X1 _17694_ (.A1(_04060_),
    .A2(_03073_),
    .B1(_03077_),
    .B2(_04041_),
    .ZN(_04080_));
 NOR2_X1 _17695_ (.A1(_04044_),
    .A2(_03095_),
    .ZN(_04081_));
 NOR3_X1 _17696_ (.A1(_04079_),
    .A2(_04080_),
    .A3(_04081_),
    .ZN(_04082_));
 NOR2_X1 _17697_ (.A1(_04032_),
    .A2(_04082_),
    .ZN(net370));
 BUF_X8 _17698_ (.A(_04031_),
    .Z(_04083_));
 OAI22_X1 _17699_ (.A1(_04051_),
    .A2(_03102_),
    .B1(_03106_),
    .B2(_04049_),
    .ZN(_04084_));
 OAI22_X1 _17700_ (.A1(_04035_),
    .A2(_03111_),
    .B1(_03115_),
    .B2(_04052_),
    .ZN(_04085_));
 NOR2_X1 _17701_ (.A1(_04084_),
    .A2(_04085_),
    .ZN(_04086_));
 NAND2_X1 _17702_ (.A1(_04057_),
    .A2(_03132_),
    .ZN(_04087_));
 AOI21_X2 _17703_ (.A(_04083_),
    .B1(_04086_),
    .B2(_04087_),
    .ZN(net371));
 OAI22_X2 _17704_ (.A1(_04059_),
    .A2(_03141_),
    .B1(_03147_),
    .B2(_04060_),
    .ZN(_04088_));
 OAI22_X2 _17705_ (.A1(_04035_),
    .A2(_03137_),
    .B1(_03151_),
    .B2(_04052_),
    .ZN(_04089_));
 NOR2_X2 _17706_ (.A1(_04088_),
    .A2(_04089_),
    .ZN(_04090_));
 NAND2_X1 _17707_ (.A1(_04057_),
    .A2(_03168_),
    .ZN(_04091_));
 AOI21_X4 _17708_ (.A(_04083_),
    .B1(_04090_),
    .B2(_04091_),
    .ZN(net372));
 OAI22_X1 _17709_ (.A1(_04065_),
    .A2(_03173_),
    .B1(_03178_),
    .B2(_04036_),
    .ZN(_04092_));
 OAI22_X1 _17710_ (.A1(_04039_),
    .A2(_03183_),
    .B1(_03188_),
    .B2(_04041_),
    .ZN(_04093_));
 NOR2_X1 _17711_ (.A1(_04044_),
    .A2(_03209_),
    .ZN(_04094_));
 NOR3_X1 _17712_ (.A1(_04092_),
    .A2(_04093_),
    .A3(_04094_),
    .ZN(_04095_));
 NOR2_X1 _17713_ (.A1(_04032_),
    .A2(_04095_),
    .ZN(net373));
 BUF_X4 _17714_ (.A(_04040_),
    .Z(_04096_));
 OAI22_X1 _17715_ (.A1(_04096_),
    .A2(_03216_),
    .B1(_03220_),
    .B2(_04078_),
    .ZN(_04097_));
 BUF_X4 _17716_ (.A(_04034_),
    .Z(_04098_));
 CLKBUF_X3 _17717_ (.A(_06085_),
    .Z(_04099_));
 OAI22_X1 _17718_ (.A1(_04098_),
    .A2(_03228_),
    .B1(_03234_),
    .B2(_04099_),
    .ZN(_04100_));
 NOR2_X1 _17719_ (.A1(_04044_),
    .A2(_03253_),
    .ZN(_04101_));
 NOR3_X1 _17720_ (.A1(_04097_),
    .A2(_04100_),
    .A3(_04101_),
    .ZN(_04102_));
 NOR2_X2 _17721_ (.A1(_04032_),
    .A2(_04102_),
    .ZN(net374));
 OAI22_X1 _17722_ (.A1(_04065_),
    .A2(_03259_),
    .B1(_03264_),
    .B2(_04036_),
    .ZN(_04103_));
 OAI22_X1 _17723_ (.A1(_04039_),
    .A2(_03269_),
    .B1(_03273_),
    .B2(_04041_),
    .ZN(_04104_));
 NOR2_X1 _17724_ (.A1(_04044_),
    .A2(_03294_),
    .ZN(_04105_));
 NOR3_X1 _17725_ (.A1(_04103_),
    .A2(_04104_),
    .A3(_04105_),
    .ZN(_04106_));
 NOR2_X1 _17726_ (.A1(_04032_),
    .A2(_04106_),
    .ZN(net375));
 OAI22_X2 _17727_ (.A1(_04059_),
    .A2(_03305_),
    .B1(_03310_),
    .B2(_04098_),
    .ZN(_04107_));
 OAI22_X2 _17728_ (.A1(_04051_),
    .A2(_03301_),
    .B1(_03314_),
    .B2(_04052_),
    .ZN(_04108_));
 NOR2_X2 _17729_ (.A1(_04107_),
    .A2(_04108_),
    .ZN(_04109_));
 NAND2_X1 _17730_ (.A1(_04057_),
    .A2(_03331_),
    .ZN(_04110_));
 AOI21_X4 _17731_ (.A(_04083_),
    .B1(_04109_),
    .B2(_04110_),
    .ZN(net376));
 OAI22_X1 _17732_ (.A1(_04065_),
    .A2(_03336_),
    .B1(_03346_),
    .B2(_04078_),
    .ZN(_04111_));
 OAI22_X1 _17733_ (.A1(_04060_),
    .A2(_03341_),
    .B1(_03350_),
    .B2(_04041_),
    .ZN(_04112_));
 NOR2_X1 _17734_ (.A1(_04044_),
    .A2(_03369_),
    .ZN(_04113_));
 NOR3_X1 _17735_ (.A1(_04111_),
    .A2(_04112_),
    .A3(_04113_),
    .ZN(_04114_));
 NOR2_X1 _17736_ (.A1(_04032_),
    .A2(_04114_),
    .ZN(net377));
 INV_X2 _17737_ (.A(_04033_),
    .ZN(_04115_));
 INV_X1 _17738_ (.A(_06085_),
    .ZN(_04116_));
 BUF_X4 _17739_ (.A(_04116_),
    .Z(_04117_));
 AOI22_X1 _17740_ (.A1(_04115_),
    .A2(_05775_),
    .B1(_06080_),
    .B2(_04117_),
    .ZN(_04118_));
 BUF_X4 _17741_ (.A(_04040_),
    .Z(_04119_));
 OAI221_X1 _17742_ (.A(_04118_),
    .B1(_03374_),
    .B2(_04048_),
    .C1(_04119_),
    .C2(_02494_),
    .ZN(_04120_));
 BUF_X4 _17743_ (.A(_04055_),
    .Z(_04121_));
 AOI21_X1 _17744_ (.A(_04120_),
    .B1(_07132_),
    .B2(_04121_),
    .ZN(_04122_));
 NOR2_X1 _17745_ (.A1(_04032_),
    .A2(_04122_),
    .ZN(net378));
 INV_X1 _17746_ (.A(_04038_),
    .ZN(_04123_));
 BUF_X4 _17747_ (.A(_04123_),
    .Z(_04124_));
 AOI22_X2 _17748_ (.A1(_05754_),
    .A2(_05849_),
    .B1(_05796_),
    .B2(_04124_),
    .ZN(_04125_));
 BUF_X4 _17749_ (.A(_04033_),
    .Z(_04126_));
 CLKBUF_X3 _17750_ (.A(_06085_),
    .Z(_04127_));
 OAI221_X2 _17751_ (.A(_04125_),
    .B1(_03383_),
    .B2(_04126_),
    .C1(_04127_),
    .C2(_03382_),
    .ZN(_04128_));
 AOI21_X1 _17752_ (.A(_04128_),
    .B1(_07156_),
    .B2(_04121_),
    .ZN(_04129_));
 NOR2_X1 _17753_ (.A1(_04032_),
    .A2(_04129_),
    .ZN(net379));
 CLKBUF_X3 _17754_ (.A(_04031_),
    .Z(_04130_));
 AOI22_X1 _17755_ (.A1(_05754_),
    .A2(_05839_),
    .B1(_05799_),
    .B2(_04124_),
    .ZN(_04131_));
 OAI221_X1 _17756_ (.A(_04131_),
    .B1(_03389_),
    .B2(_04126_),
    .C1(_04127_),
    .C2(_03388_),
    .ZN(_04132_));
 AOI21_X1 _17757_ (.A(_04132_),
    .B1(_05956_),
    .B2(_04121_),
    .ZN(_04133_));
 NOR2_X1 _17758_ (.A1(_04130_),
    .A2(_04133_),
    .ZN(net380));
 AOI22_X1 _17759_ (.A1(_05754_),
    .A2(_05829_),
    .B1(_05802_),
    .B2(_04124_),
    .ZN(_04134_));
 OAI221_X1 _17760_ (.A(_04134_),
    .B1(_03395_),
    .B2(_04126_),
    .C1(_04127_),
    .C2(_03393_),
    .ZN(_04135_));
 BUF_X4 _17761_ (.A(_04056_),
    .Z(_04136_));
 AOI21_X1 _17762_ (.A(_04135_),
    .B1(_05902_),
    .B2(_04136_),
    .ZN(_04137_));
 NOR2_X1 _17763_ (.A1(_04130_),
    .A2(_04137_),
    .ZN(net381));
 AOI22_X1 _17764_ (.A1(_05754_),
    .A2(_05832_),
    .B1(_05792_),
    .B2(_04123_),
    .ZN(_04138_));
 OAI221_X1 _17765_ (.A(_04138_),
    .B1(_03400_),
    .B2(_04126_),
    .C1(_04127_),
    .C2(_03399_),
    .ZN(_04139_));
 AOI21_X1 _17766_ (.A(_04139_),
    .B1(_03403_),
    .B2(_04136_),
    .ZN(_04140_));
 NOR2_X1 _17767_ (.A1(_04130_),
    .A2(_04140_),
    .ZN(net382));
 AOI22_X1 _17768_ (.A1(_05754_),
    .A2(_05836_),
    .B1(_05809_),
    .B2(_04123_),
    .ZN(_04141_));
 OAI221_X1 _17769_ (.A(_04141_),
    .B1(_07233_),
    .B2(_04126_),
    .C1(_04127_),
    .C2(_07196_),
    .ZN(_04142_));
 AOI21_X1 _17770_ (.A(_04142_),
    .B1(_05972_),
    .B2(_04136_),
    .ZN(_04143_));
 NOR2_X1 _17771_ (.A1(_04130_),
    .A2(_04143_),
    .ZN(net383));
 AOI22_X1 _17772_ (.A1(_05754_),
    .A2(_05843_),
    .B1(_05806_),
    .B2(_04123_),
    .ZN(_04144_));
 OAI221_X1 _17773_ (.A(_04144_),
    .B1(_07229_),
    .B2(_04126_),
    .C1(_04127_),
    .C2(_07192_),
    .ZN(_04145_));
 AOI21_X1 _17774_ (.A(_04145_),
    .B1(_06008_),
    .B2(_04136_),
    .ZN(_04146_));
 NOR2_X1 _17775_ (.A1(_04130_),
    .A2(_04146_),
    .ZN(net384));
 AOI22_X1 _17776_ (.A1(_04115_),
    .A2(_05778_),
    .B1(_06071_),
    .B2(_04117_),
    .ZN(_04147_));
 OAI221_X1 _17777_ (.A(_04147_),
    .B1(_03412_),
    .B2(_04048_),
    .C1(_04119_),
    .C2(_07105_),
    .ZN(_04148_));
 AOI21_X1 _17778_ (.A(_04148_),
    .B1(_05993_),
    .B2(_04136_),
    .ZN(_04149_));
 NOR2_X1 _17779_ (.A1(_04130_),
    .A2(_04149_),
    .ZN(net385));
 OAI22_X1 _17780_ (.A1(_04065_),
    .A2(_03418_),
    .B1(_03422_),
    .B2(_04078_),
    .ZN(_04150_));
 OAI22_X1 _17781_ (.A1(_04060_),
    .A2(_03428_),
    .B1(_03432_),
    .B2(_04041_),
    .ZN(_04151_));
 NOR2_X1 _17782_ (.A1(_04044_),
    .A2(_03450_),
    .ZN(_04152_));
 NOR3_X1 _17783_ (.A1(_04150_),
    .A2(_04151_),
    .A3(_04152_),
    .ZN(_04153_));
 NOR2_X1 _17784_ (.A1(_04130_),
    .A2(_04153_),
    .ZN(net386));
 AOI22_X1 _17785_ (.A1(_06575_),
    .A2(_06524_),
    .B1(_05492_),
    .B2(_04115_),
    .ZN(_04154_));
 OAI221_X1 _17786_ (.A(_04154_),
    .B1(_05274_),
    .B2(_04048_),
    .C1(_04127_),
    .C2(_06099_),
    .ZN(_04155_));
 AOI21_X1 _17787_ (.A(_04155_),
    .B1(_06179_),
    .B2(_04136_),
    .ZN(_04156_));
 NOR2_X1 _17788_ (.A1(_04130_),
    .A2(_04156_),
    .ZN(net387));
 AOI22_X1 _17789_ (.A1(_04124_),
    .A2(_06514_),
    .B1(_06100_),
    .B2(_04117_),
    .ZN(_04157_));
 OAI221_X1 _17790_ (.A(_04157_),
    .B1(_06789_),
    .B2(_04126_),
    .C1(_04119_),
    .C2(_05376_),
    .ZN(_04158_));
 AOI21_X1 _17791_ (.A(_04158_),
    .B1(_06146_),
    .B2(_04136_),
    .ZN(_04159_));
 NOR2_X1 _17792_ (.A1(_04130_),
    .A2(_04159_),
    .ZN(net388));
 AOI22_X2 _17793_ (.A1(_06575_),
    .A2(_05370_),
    .B1(_05613_),
    .B2(_04117_),
    .ZN(_04160_));
 OAI221_X2 _17794_ (.A(_04160_),
    .B1(_06513_),
    .B2(_04048_),
    .C1(_04098_),
    .C2(_06548_),
    .ZN(_04161_));
 AOI21_X1 _17795_ (.A(_04161_),
    .B1(_06163_),
    .B2(_04136_),
    .ZN(_04162_));
 NOR2_X1 _17796_ (.A1(_04130_),
    .A2(_04162_),
    .ZN(net389));
 BUF_X4 _17797_ (.A(_04031_),
    .Z(_04163_));
 OAI22_X1 _17798_ (.A1(_04065_),
    .A2(_03465_),
    .B1(_03471_),
    .B2(_04036_),
    .ZN(_04164_));
 OAI22_X1 _17799_ (.A1(_04039_),
    .A2(_03476_),
    .B1(_03480_),
    .B2(_04040_),
    .ZN(_04165_));
 NOR2_X1 _17800_ (.A1(_04044_),
    .A2(_03498_),
    .ZN(_04166_));
 NOR3_X1 _17801_ (.A1(_04164_),
    .A2(_04165_),
    .A3(_04166_),
    .ZN(_04167_));
 NOR2_X1 _17802_ (.A1(_04163_),
    .A2(_04167_),
    .ZN(net390));
 AOI22_X1 _17803_ (.A1(_04117_),
    .A2(_10225_),
    .B1(_10348_),
    .B2(_04115_),
    .ZN(_04168_));
 OAI221_X1 _17804_ (.A(_04168_),
    .B1(_03502_),
    .B2(_04048_),
    .C1(_04119_),
    .C2(_05327_),
    .ZN(_04169_));
 AOI21_X1 _17805_ (.A(_04169_),
    .B1(_10417_),
    .B2(_04136_),
    .ZN(_04170_));
 NOR2_X1 _17806_ (.A1(_04163_),
    .A2(_04170_),
    .ZN(net391));
 AOI22_X1 _17807_ (.A1(_04115_),
    .A2(_07302_),
    .B1(net694),
    .B2(_06575_),
    .ZN(_04171_));
 OAI221_X1 _17808_ (.A(_04171_),
    .B1(_10255_),
    .B2(_04048_),
    .C1(_04127_),
    .C2(_10221_),
    .ZN(_04172_));
 AOI21_X1 _17809_ (.A(_04172_),
    .B1(_07676_),
    .B2(_04136_),
    .ZN(_04173_));
 NOR2_X2 _17810_ (.A1(_04163_),
    .A2(_04173_),
    .ZN(net392));
 OAI22_X2 _17811_ (.A1(_04038_),
    .A2(_10261_),
    .B1(_10357_),
    .B2(_04033_),
    .ZN(_04174_));
 INV_X1 _17812_ (.A(_10315_),
    .ZN(_04175_));
 AOI221_X2 _17813_ (.A(_04174_),
    .B1(_07434_),
    .B2(_04117_),
    .C1(_05754_),
    .C2(_04175_),
    .ZN(_04176_));
 NAND2_X1 _17814_ (.A1(_04057_),
    .A2(_07661_),
    .ZN(_04177_));
 AOI21_X2 _17815_ (.A(_04083_),
    .B1(_04176_),
    .B2(_04177_),
    .ZN(net393));
 OAI22_X2 _17816_ (.A1(_04038_),
    .A2(_10258_),
    .B1(_10354_),
    .B2(_04033_),
    .ZN(_04178_));
 INV_X1 _17817_ (.A(_10312_),
    .ZN(_04179_));
 AOI221_X2 _17818_ (.A(_04178_),
    .B1(net742),
    .B2(_04117_),
    .C1(_05754_),
    .C2(_04179_),
    .ZN(_04180_));
 NAND2_X1 _17819_ (.A1(_04057_),
    .A2(_07409_),
    .ZN(_04181_));
 AOI21_X2 _17820_ (.A(_04083_),
    .B1(_04180_),
    .B2(_04181_),
    .ZN(net394));
 OAI22_X2 _17821_ (.A1(_04038_),
    .A2(_10273_),
    .B1(net697),
    .B2(_07022_),
    .ZN(_04182_));
 AOI221_X2 _17822_ (.A(_04182_),
    .B1(_03518_),
    .B2(_04115_),
    .C1(_04117_),
    .C2(net675),
    .ZN(_04183_));
 NAND2_X1 _17823_ (.A1(_04057_),
    .A2(_07646_),
    .ZN(_04184_));
 AOI21_X2 _17824_ (.A(_04083_),
    .B1(_04183_),
    .B2(_04184_),
    .ZN(net395));
 AOI22_X1 _17825_ (.A1(_04124_),
    .A2(_07279_),
    .B1(net664),
    .B2(_06575_),
    .ZN(_04185_));
 OAI221_X1 _17826_ (.A(_04185_),
    .B1(_10366_),
    .B2(_04034_),
    .C1(_04127_),
    .C2(_10209_),
    .ZN(_04186_));
 AOI21_X1 _17827_ (.A(_04186_),
    .B1(_07631_),
    .B2(_04056_),
    .ZN(_04187_));
 NOR2_X1 _17828_ (.A1(_04163_),
    .A2(_04187_),
    .ZN(net396));
 OAI22_X1 _17829_ (.A1(_04060_),
    .A2(_03530_),
    .B1(_03534_),
    .B2(_04078_),
    .ZN(_04188_));
 OAI22_X1 _17830_ (.A1(_04098_),
    .A2(_03539_),
    .B1(_03543_),
    .B2(_04040_),
    .ZN(_04189_));
 CLKBUF_X3 _17831_ (.A(_04043_),
    .Z(_04190_));
 NOR2_X1 _17832_ (.A1(_04190_),
    .A2(_03562_),
    .ZN(_04191_));
 NOR3_X1 _17833_ (.A1(_04188_),
    .A2(_04189_),
    .A3(_04191_),
    .ZN(_04192_));
 NOR2_X2 _17834_ (.A1(_04163_),
    .A2(_04192_),
    .ZN(net397));
 AOI22_X1 _17835_ (.A1(_04124_),
    .A2(_07473_),
    .B1(_07506_),
    .B2(_06575_),
    .ZN(_04193_));
 OAI221_X1 _17836_ (.A(_04193_),
    .B1(_10363_),
    .B2(_04034_),
    .C1(_04127_),
    .C2(_10206_),
    .ZN(_04194_));
 AOI21_X1 _17837_ (.A(_04194_),
    .B1(_07616_),
    .B2(_04056_),
    .ZN(_04195_));
 NOR2_X1 _17838_ (.A1(_04163_),
    .A2(_04195_),
    .ZN(net398));
 OAI22_X1 _17839_ (.A1(_04059_),
    .A2(net640),
    .B1(net632),
    .B2(_04096_),
    .ZN(_04196_));
 OAI22_X1 _17840_ (.A1(_04051_),
    .A2(net650),
    .B1(net713),
    .B2(_04098_),
    .ZN(_04197_));
 NOR2_X1 _17841_ (.A1(_04196_),
    .A2(_04197_),
    .ZN(_04198_));
 NAND2_X1 _17842_ (.A1(_04057_),
    .A2(_07394_),
    .ZN(_04199_));
 AOI21_X2 _17843_ (.A(_04083_),
    .B1(_04198_),
    .B2(_04199_),
    .ZN(net399));
 AOI22_X1 _17844_ (.A1(_04124_),
    .A2(_10249_),
    .B1(_10276_),
    .B2(_06575_),
    .ZN(_04200_));
 OAI221_X1 _17845_ (.A(_04200_),
    .B1(_03574_),
    .B2(_04034_),
    .C1(_04036_),
    .C2(net685),
    .ZN(_04201_));
 AOI21_X1 _17846_ (.A(_04201_),
    .B1(_10372_),
    .B2(_04056_),
    .ZN(_04202_));
 NOR2_X1 _17847_ (.A1(_04163_),
    .A2(_04202_),
    .ZN(net400));
 OAI22_X1 _17848_ (.A1(_04035_),
    .A2(_10342_),
    .B1(net771),
    .B2(_04049_),
    .ZN(_04203_));
 OAI22_X1 _17849_ (.A1(_04051_),
    .A2(net643),
    .B1(_10279_),
    .B2(_04119_),
    .ZN(_04204_));
 NOR2_X1 _17850_ (.A1(_04203_),
    .A2(_04204_),
    .ZN(_04205_));
 NAND2_X1 _17851_ (.A1(_04121_),
    .A2(_07556_),
    .ZN(_04206_));
 AOI21_X2 _17852_ (.A(_04083_),
    .B1(_04205_),
    .B2(_04206_),
    .ZN(net401));
 AOI22_X1 _17853_ (.A1(_04124_),
    .A2(_03583_),
    .B1(net688),
    .B2(_06575_),
    .ZN(_04207_));
 OAI221_X1 _17854_ (.A(_04207_),
    .B1(net723),
    .B2(_04034_),
    .C1(_04036_),
    .C2(net646),
    .ZN(_04208_));
 AOI21_X1 _17855_ (.A(_04208_),
    .B1(_07571_),
    .B2(_04056_),
    .ZN(_04209_));
 NOR2_X2 _17856_ (.A1(_04163_),
    .A2(_04209_),
    .ZN(net402));
 INV_X2 _17857_ (.A(_10185_),
    .ZN(_04210_));
 INV_X1 _17858_ (.A(_10285_),
    .ZN(_04211_));
 AOI22_X1 _17859_ (.A1(_04117_),
    .A2(_04210_),
    .B1(_04211_),
    .B2(_06575_),
    .ZN(_04212_));
 BUF_X4 _17860_ (.A(_04034_),
    .Z(_04213_));
 OAI221_X1 _17861_ (.A(_04212_),
    .B1(_10240_),
    .B2(_04048_),
    .C1(_04213_),
    .C2(_10336_),
    .ZN(_04214_));
 AOI21_X1 _17862_ (.A(_04214_),
    .B1(_07342_),
    .B2(_04056_),
    .ZN(_04215_));
 NOR2_X1 _17863_ (.A1(_04163_),
    .A2(_04215_),
    .ZN(net403));
 OAI22_X1 _17864_ (.A1(_04051_),
    .A2(net647),
    .B1(_10237_),
    .B2(_04049_),
    .ZN(_04216_));
 OAI22_X1 _17865_ (.A1(_04035_),
    .A2(_10333_),
    .B1(_10288_),
    .B2(_04119_),
    .ZN(_04217_));
 NOR2_X1 _17866_ (.A1(_04216_),
    .A2(_04217_),
    .ZN(_04218_));
 NAND2_X1 _17867_ (.A1(_04121_),
    .A2(_07376_),
    .ZN(_04219_));
 AOI21_X2 _17868_ (.A(_04083_),
    .B1(_04218_),
    .B2(_04219_),
    .ZN(net404));
 INV_X2 _17869_ (.A(net686),
    .ZN(_04220_));
 AOI22_X1 _17870_ (.A1(_04117_),
    .A2(_04220_),
    .B1(_07489_),
    .B2(_06575_),
    .ZN(_04221_));
 OAI221_X1 _17871_ (.A(_04221_),
    .B1(net732),
    .B2(_04048_),
    .C1(_04213_),
    .C2(net703),
    .ZN(_04222_));
 AOI21_X1 _17872_ (.A(_04222_),
    .B1(_07361_),
    .B2(_04056_),
    .ZN(_04223_));
 NOR2_X1 _17873_ (.A1(_04163_),
    .A2(_04223_),
    .ZN(net405));
 OAI22_X1 _17874_ (.A1(_04059_),
    .A2(net751),
    .B1(_10327_),
    .B2(_04098_),
    .ZN(_04224_));
 OAI22_X1 _17875_ (.A1(_04051_),
    .A2(_10194_),
    .B1(_10294_),
    .B2(_04119_),
    .ZN(_04225_));
 NOR2_X1 _17876_ (.A1(_04224_),
    .A2(_04225_),
    .ZN(_04226_));
 NAND2_X1 _17877_ (.A1(_04121_),
    .A2(_07601_),
    .ZN(_04227_));
 AOI21_X2 _17878_ (.A(_04083_),
    .B1(_04226_),
    .B2(_04227_),
    .ZN(net406));
 OAI22_X1 _17879_ (.A1(_04051_),
    .A2(_10191_),
    .B1(net670),
    .B2(_04098_),
    .ZN(_04228_));
 OAI22_X1 _17880_ (.A1(_04059_),
    .A2(_10228_),
    .B1(_10297_),
    .B2(_04119_),
    .ZN(_04229_));
 NOR2_X1 _17881_ (.A1(_04228_),
    .A2(_04229_),
    .ZN(_04230_));
 NAND2_X1 _17882_ (.A1(_04121_),
    .A2(_07586_),
    .ZN(_04231_));
 AOI21_X4 _17883_ (.A(_04031_),
    .B1(_04230_),
    .B2(_04231_),
    .ZN(net407));
 OAI22_X1 _17884_ (.A1(_04059_),
    .A2(_03614_),
    .B1(_03619_),
    .B2(_04098_),
    .ZN(_04232_));
 OAI22_X1 _17885_ (.A1(_04051_),
    .A2(_03610_),
    .B1(_03623_),
    .B2(_04119_),
    .ZN(_04233_));
 NOR2_X1 _17886_ (.A1(_04232_),
    .A2(_04233_),
    .ZN(_04234_));
 NAND2_X1 _17887_ (.A1(_04121_),
    .A2(_03640_),
    .ZN(_04235_));
 AOI21_X2 _17888_ (.A(_04031_),
    .B1(_04234_),
    .B2(_04235_),
    .ZN(net408));
 BUF_X4 _17889_ (.A(_04031_),
    .Z(_04236_));
 OAI22_X1 _17890_ (.A1(_04059_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(_04036_),
    .ZN(_04237_));
 OAI22_X1 _17891_ (.A1(_04096_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_04213_),
    .ZN(_04238_));
 NOR2_X1 _17892_ (.A1(_04190_),
    .A2(_03655_),
    .ZN(_04239_));
 NOR3_X1 _17893_ (.A1(_04237_),
    .A2(_04238_),
    .A3(_04239_),
    .ZN(_04240_));
 NOR2_X2 _17894_ (.A1(_04236_),
    .A2(_04240_),
    .ZN(net409));
 AOI22_X1 _17895_ (.A1(_04124_),
    .A2(_05189_),
    .B1(_05649_),
    .B2(_04116_),
    .ZN(_04241_));
 OAI221_X1 _17896_ (.A(_04241_),
    .B1(_03662_),
    .B2(_04034_),
    .C1(_04041_),
    .C2(_03660_),
    .ZN(_04242_));
 AOI21_X1 _17897_ (.A(_04242_),
    .B1(_06249_),
    .B2(_04056_),
    .ZN(_04243_));
 NOR2_X1 _17898_ (.A1(_04236_),
    .A2(_04243_),
    .ZN(net410));
 OAI22_X1 _17899_ (.A1(_04049_),
    .A2(_03666_),
    .B1(_03669_),
    .B2(_04036_),
    .ZN(_04244_));
 OAI22_X1 _17900_ (.A1(_04096_),
    .A2(_03672_),
    .B1(_03674_),
    .B2(_04213_),
    .ZN(_04245_));
 NOR2_X1 _17901_ (.A1(_04190_),
    .A2(_03677_),
    .ZN(_04246_));
 NOR3_X1 _17902_ (.A1(_04244_),
    .A2(_04245_),
    .A3(_04246_),
    .ZN(_04247_));
 NOR2_X2 _17903_ (.A1(_04236_),
    .A2(_04247_),
    .ZN(net411));
 OAI22_X1 _17904_ (.A1(_04049_),
    .A2(_03681_),
    .B1(_03683_),
    .B2(_04213_),
    .ZN(_04248_));
 OAI22_X1 _17905_ (.A1(_04052_),
    .A2(_03686_),
    .B1(_03689_),
    .B2(_04099_),
    .ZN(_04249_));
 NOR2_X1 _17906_ (.A1(_04190_),
    .A2(_03692_),
    .ZN(_04250_));
 NOR3_X1 _17907_ (.A1(_04248_),
    .A2(_04249_),
    .A3(_04250_),
    .ZN(_04251_));
 NOR2_X2 _17908_ (.A1(_04236_),
    .A2(_04251_),
    .ZN(net412));
 OAI22_X1 _17909_ (.A1(_04049_),
    .A2(_03696_),
    .B1(_03699_),
    .B2(_04099_),
    .ZN(_04252_));
 OAI22_X1 _17910_ (.A1(_04052_),
    .A2(_03702_),
    .B1(_03704_),
    .B2(_04126_),
    .ZN(_04253_));
 NOR2_X1 _17911_ (.A1(_04190_),
    .A2(_03707_),
    .ZN(_04254_));
 NOR3_X1 _17912_ (.A1(_04252_),
    .A2(_04253_),
    .A3(_04254_),
    .ZN(_04255_));
 NOR2_X2 _17913_ (.A1(_04236_),
    .A2(_04255_),
    .ZN(net413));
 OAI22_X1 _17914_ (.A1(_04096_),
    .A2(_03712_),
    .B1(_03714_),
    .B2(_04213_),
    .ZN(_04256_));
 OAI22_X1 _17915_ (.A1(_04039_),
    .A2(_03717_),
    .B1(_03720_),
    .B2(_04099_),
    .ZN(_04257_));
 NOR2_X1 _17916_ (.A1(_04190_),
    .A2(_03723_),
    .ZN(_04258_));
 NOR3_X1 _17917_ (.A1(_04256_),
    .A2(_04257_),
    .A3(_04258_),
    .ZN(_04259_));
 NOR2_X2 _17918_ (.A1(_04236_),
    .A2(_04259_),
    .ZN(net414));
 OAI22_X1 _17919_ (.A1(_04035_),
    .A2(_03727_),
    .B1(_03730_),
    .B2(_04060_),
    .ZN(_04260_));
 OAI22_X1 _17920_ (.A1(_04059_),
    .A2(_03733_),
    .B1(_03735_),
    .B2(_04119_),
    .ZN(_04261_));
 NOR2_X1 _17921_ (.A1(_04260_),
    .A2(_04261_),
    .ZN(_04262_));
 NAND2_X1 _17922_ (.A1(_04121_),
    .A2(_03738_),
    .ZN(_04263_));
 AOI21_X2 _17923_ (.A(_04031_),
    .B1(_04262_),
    .B2(_04263_),
    .ZN(net415));
 OAI22_X1 _17924_ (.A1(_04096_),
    .A2(_03741_),
    .B1(_03743_),
    .B2(_04213_),
    .ZN(_04264_));
 OAI22_X1 _17925_ (.A1(_04039_),
    .A2(_03746_),
    .B1(_03749_),
    .B2(_04099_),
    .ZN(_04265_));
 NOR2_X1 _17926_ (.A1(_04190_),
    .A2(_03752_),
    .ZN(_04266_));
 NOR3_X1 _17927_ (.A1(_04264_),
    .A2(_04265_),
    .A3(_04266_),
    .ZN(_04267_));
 NOR2_X2 _17928_ (.A1(_04236_),
    .A2(_04267_),
    .ZN(net416));
 OAI22_X1 _17929_ (.A1(_04049_),
    .A2(_03756_),
    .B1(_03759_),
    .B2(_04099_),
    .ZN(_04268_));
 OAI22_X1 _17930_ (.A1(_04052_),
    .A2(_03762_),
    .B1(_03764_),
    .B2(_04126_),
    .ZN(_04269_));
 NOR2_X1 _17931_ (.A1(_04190_),
    .A2(_03767_),
    .ZN(_04270_));
 NOR3_X1 _17932_ (.A1(_04268_),
    .A2(_04269_),
    .A3(_04270_),
    .ZN(_04271_));
 NOR2_X2 _17933_ (.A1(_04236_),
    .A2(_04271_),
    .ZN(net417));
 OAI22_X1 _17934_ (.A1(_04096_),
    .A2(_03771_),
    .B1(_03773_),
    .B2(_04213_),
    .ZN(_04272_));
 OAI22_X1 _17935_ (.A1(_04039_),
    .A2(_03776_),
    .B1(_03779_),
    .B2(_04099_),
    .ZN(_04273_));
 NOR2_X1 _17936_ (.A1(_04190_),
    .A2(_03782_),
    .ZN(_04274_));
 NOR3_X1 _17937_ (.A1(_04272_),
    .A2(_04273_),
    .A3(_04274_),
    .ZN(_04275_));
 NOR2_X2 _17938_ (.A1(_04236_),
    .A2(_04275_),
    .ZN(net418));
 OAI22_X1 _17939_ (.A1(_04065_),
    .A2(_03788_),
    .B1(_03798_),
    .B2(_04078_),
    .ZN(_04276_));
 OAI22_X1 _17940_ (.A1(_04060_),
    .A2(_03793_),
    .B1(_03802_),
    .B2(_04040_),
    .ZN(_04277_));
 NOR2_X1 _17941_ (.A1(_04190_),
    .A2(_03820_),
    .ZN(_04278_));
 NOR3_X1 _17942_ (.A1(_04276_),
    .A2(_04277_),
    .A3(_04278_),
    .ZN(_04279_));
 NOR2_X2 _17943_ (.A1(_04236_),
    .A2(_04279_),
    .ZN(net419));
 AOI22_X1 _17944_ (.A1(_04124_),
    .A2(_05194_),
    .B1(_05639_),
    .B2(_04116_),
    .ZN(_04280_));
 INV_X1 _17945_ (.A(_05556_),
    .ZN(_04281_));
 INV_X1 _17946_ (.A(_05427_),
    .ZN(_04282_));
 OAI221_X1 _17947_ (.A(_04280_),
    .B1(_04281_),
    .B2(_04034_),
    .C1(_04041_),
    .C2(_04282_),
    .ZN(_04283_));
 AOI21_X1 _17948_ (.A(_04283_),
    .B1(_03827_),
    .B2(_04056_),
    .ZN(_04284_));
 NOR2_X2 _17949_ (.A1(_04047_),
    .A2(_04284_),
    .ZN(net420));
 OAI22_X1 _17950_ (.A1(_04096_),
    .A2(_03836_),
    .B1(_03833_),
    .B2(_04213_),
    .ZN(_04285_));
 OAI22_X1 _17951_ (.A1(_04039_),
    .A2(_03831_),
    .B1(_03839_),
    .B2(_06085_),
    .ZN(_04286_));
 NOR2_X1 _17952_ (.A1(_04043_),
    .A2(_03849_),
    .ZN(_04287_));
 NOR3_X1 _17953_ (.A1(_04285_),
    .A2(_04286_),
    .A3(_04287_),
    .ZN(_04288_));
 NOR2_X2 _17954_ (.A1(_04047_),
    .A2(_04288_),
    .ZN(net421));
 OAI22_X1 _17955_ (.A1(_04059_),
    .A2(_03853_),
    .B1(_03855_),
    .B2(_04096_),
    .ZN(_04289_));
 OAI22_X1 _17956_ (.A1(_04035_),
    .A2(_03858_),
    .B1(_03861_),
    .B2(_04060_),
    .ZN(_04290_));
 NOR2_X1 _17957_ (.A1(_04289_),
    .A2(_04290_),
    .ZN(_04291_));
 NAND2_X1 _17958_ (.A1(_04121_),
    .A2(_03864_),
    .ZN(_04292_));
 AOI21_X4 _17959_ (.A(_04031_),
    .B1(_04291_),
    .B2(_04292_),
    .ZN(net422));
 OAI22_X1 _17960_ (.A1(_04049_),
    .A2(_03867_),
    .B1(_03875_),
    .B2(_04099_),
    .ZN(_04293_));
 OAI22_X1 _17961_ (.A1(_04052_),
    .A2(_03872_),
    .B1(_03869_),
    .B2(_04126_),
    .ZN(_04294_));
 NOR2_X1 _17962_ (.A1(_04043_),
    .A2(_06229_),
    .ZN(_04295_));
 NOR3_X1 _17963_ (.A1(_04293_),
    .A2(_04294_),
    .A3(_04295_),
    .ZN(_04296_));
 NOR2_X2 _17964_ (.A1(_04047_),
    .A2(_04296_),
    .ZN(net423));
 OAI22_X1 _17965_ (.A1(_04065_),
    .A2(_03882_),
    .B1(_03887_),
    .B2(_04099_),
    .ZN(_04297_));
 OAI22_X1 _17966_ (.A1(_04078_),
    .A2(_03892_),
    .B1(_03896_),
    .B2(_04040_),
    .ZN(_04298_));
 NOR2_X1 _17967_ (.A1(_04043_),
    .A2(_03914_),
    .ZN(_04299_));
 NOR3_X1 _17968_ (.A1(_04297_),
    .A2(_04298_),
    .A3(_04299_),
    .ZN(_04300_));
 NOR2_X2 _17969_ (.A1(_04047_),
    .A2(_04300_),
    .ZN(net424));
 OAI22_X1 _17970_ (.A1(_04098_),
    .A2(_03920_),
    .B1(_03925_),
    .B2(_04099_),
    .ZN(_04301_));
 OAI22_X1 _17971_ (.A1(_04078_),
    .A2(_03930_),
    .B1(_03934_),
    .B2(_04040_),
    .ZN(_04302_));
 NOR2_X1 _17972_ (.A1(_04043_),
    .A2(_03952_),
    .ZN(_04303_));
 NOR3_X1 _17973_ (.A1(_04301_),
    .A2(_04302_),
    .A3(_04303_),
    .ZN(_04304_));
 NOR2_X2 _17974_ (.A1(_04047_),
    .A2(_04304_),
    .ZN(net425));
 OAI22_X2 _17975_ (.A1(_04096_),
    .A2(_03958_),
    .B1(_03967_),
    .B2(_04213_),
    .ZN(_04305_));
 OAI22_X2 _17976_ (.A1(_04078_),
    .A2(_03962_),
    .B1(_03972_),
    .B2(_06085_),
    .ZN(_04306_));
 NOR2_X1 _17977_ (.A1(_04043_),
    .A2(_03990_),
    .ZN(_04307_));
 NOR3_X2 _17978_ (.A1(_04305_),
    .A2(_04306_),
    .A3(_04307_),
    .ZN(_04308_));
 NOR2_X2 _17979_ (.A1(_04047_),
    .A2(_04308_),
    .ZN(net426));
 OAI22_X1 _17980_ (.A1(_04060_),
    .A2(_03997_),
    .B1(_04001_),
    .B2(_04078_),
    .ZN(_04309_));
 OAI22_X1 _17981_ (.A1(_04098_),
    .A2(_04006_),
    .B1(_04010_),
    .B2(_04040_),
    .ZN(_04310_));
 NOR2_X1 _17982_ (.A1(_04043_),
    .A2(_04028_),
    .ZN(_04311_));
 NOR3_X1 _17983_ (.A1(_04309_),
    .A2(_04310_),
    .A3(_04311_),
    .ZN(_04312_));
 NOR2_X2 _17984_ (.A1(_04047_),
    .A2(_04312_),
    .ZN(net427));
 BUF_X4 _17985_ (.A(_05599_),
    .Z(_04313_));
 BUF_X4 _17986_ (.A(_04313_),
    .Z(_04314_));
 BUF_X4 _17987_ (.A(_00065_),
    .Z(_04315_));
 BUF_X4 _17988_ (.A(_04315_),
    .Z(_04316_));
 BUF_X4 _17989_ (.A(_04316_),
    .Z(_04317_));
 BUF_X4 _17990_ (.A(_05592_),
    .Z(_04318_));
 BUF_X4 _17991_ (.A(_04318_),
    .Z(_04319_));
 OAI22_X1 _17992_ (.A1(_04317_),
    .A2(_02768_),
    .B1(_02777_),
    .B2(_04319_),
    .ZN(_04320_));
 BUF_X4 _17993_ (.A(_00067_),
    .Z(_04321_));
 BUF_X4 _17994_ (.A(_04321_),
    .Z(_04322_));
 BUF_X4 _17995_ (.A(_04322_),
    .Z(_04323_));
 BUF_X4 _17996_ (.A(_00066_),
    .Z(_04324_));
 BUF_X4 _17997_ (.A(_04324_),
    .Z(_04325_));
 OAI22_X1 _17998_ (.A1(_04323_),
    .A2(_02790_),
    .B1(_02798_),
    .B2(_04325_),
    .ZN(_04326_));
 CLKBUF_X3 _17999_ (.A(_07082_),
    .Z(_04327_));
 NOR2_X1 _18000_ (.A1(_04327_),
    .A2(_02840_),
    .ZN(_04328_));
 NOR3_X1 _18001_ (.A1(_04320_),
    .A2(_04326_),
    .A3(_04328_),
    .ZN(_04329_));
 NOR2_X2 _18002_ (.A1(_04314_),
    .A2(_04329_),
    .ZN(net428));
 BUF_X4 _18003_ (.A(_04313_),
    .Z(_04330_));
 BUF_X4 _18004_ (.A(_04318_),
    .Z(_04331_));
 BUF_X4 _18005_ (.A(_04315_),
    .Z(_04332_));
 OAI22_X1 _18006_ (.A1(_04331_),
    .A2(_02850_),
    .B1(_02854_),
    .B2(_04332_),
    .ZN(_04333_));
 BUF_X4 _18007_ (.A(_04322_),
    .Z(_04334_));
 BUF_X4 _18008_ (.A(_04324_),
    .Z(_04335_));
 OAI22_X1 _18009_ (.A1(_04334_),
    .A2(_02864_),
    .B1(_02868_),
    .B2(_04335_),
    .ZN(_04336_));
 NOR2_X1 _18010_ (.A1(_04333_),
    .A2(_04336_),
    .ZN(_04337_));
 NAND2_X1 _18011_ (.A1(_06977_),
    .A2(_02896_),
    .ZN(_04338_));
 AOI21_X2 _18012_ (.A(_04330_),
    .B1(_04337_),
    .B2(_04338_),
    .ZN(net429));
 OAI22_X1 _18013_ (.A1(_04317_),
    .A2(_02901_),
    .B1(_02905_),
    .B2(_04323_),
    .ZN(_04339_));
 OAI22_X1 _18014_ (.A1(_04331_),
    .A2(_02912_),
    .B1(_02916_),
    .B2(_04335_),
    .ZN(_04340_));
 NOR2_X1 _18015_ (.A1(_04339_),
    .A2(_04340_),
    .ZN(_04341_));
 NAND2_X1 _18016_ (.A1(_06977_),
    .A2(_02934_),
    .ZN(_04342_));
 AOI21_X2 _18017_ (.A(_04330_),
    .B1(_04341_),
    .B2(_04342_),
    .ZN(net430));
 BUF_X4 _18018_ (.A(_04322_),
    .Z(_04343_));
 OAI22_X2 _18019_ (.A1(_04317_),
    .A2(_02940_),
    .B1(_02952_),
    .B2(_04343_),
    .ZN(_04344_));
 BUF_X4 _18020_ (.A(_04318_),
    .Z(_04345_));
 OAI22_X2 _18021_ (.A1(_04345_),
    .A2(_02946_),
    .B1(_02956_),
    .B2(_04325_),
    .ZN(_04346_));
 NOR2_X1 _18022_ (.A1(_04327_),
    .A2(_02974_),
    .ZN(_04347_));
 NOR3_X2 _18023_ (.A1(_04344_),
    .A2(_04346_),
    .A3(_04347_),
    .ZN(_04348_));
 NOR2_X2 _18024_ (.A1(_04314_),
    .A2(_04348_),
    .ZN(net431));
 OAI22_X1 _18025_ (.A1(_04331_),
    .A2(_02981_),
    .B1(_02985_),
    .B2(_04332_),
    .ZN(_04349_));
 OAI22_X1 _18026_ (.A1(_04334_),
    .A2(_02990_),
    .B1(_02996_),
    .B2(_04335_),
    .ZN(_04350_));
 NOR2_X1 _18027_ (.A1(_04349_),
    .A2(_04350_),
    .ZN(_04351_));
 NAND2_X1 _18028_ (.A1(_06977_),
    .A2(_03013_),
    .ZN(_04352_));
 AOI21_X2 _18029_ (.A(_04330_),
    .B1(_04351_),
    .B2(_04352_),
    .ZN(net432));
 CLKBUF_X3 _18030_ (.A(_04315_),
    .Z(_04353_));
 BUF_X4 _18031_ (.A(_04318_),
    .Z(_04354_));
 OAI22_X1 _18032_ (.A1(_04353_),
    .A2(_03019_),
    .B1(_03024_),
    .B2(_04354_),
    .ZN(_04355_));
 OAI22_X1 _18033_ (.A1(_04323_),
    .A2(_03030_),
    .B1(_03034_),
    .B2(_04325_),
    .ZN(_04356_));
 NOR2_X1 _18034_ (.A1(_04327_),
    .A2(_03055_),
    .ZN(_04357_));
 NOR3_X1 _18035_ (.A1(_04355_),
    .A2(_04356_),
    .A3(_04357_),
    .ZN(_04358_));
 NOR2_X2 _18036_ (.A1(_04314_),
    .A2(_04358_),
    .ZN(net433));
 OAI22_X1 _18037_ (.A1(_04353_),
    .A2(_03061_),
    .B1(_03073_),
    .B2(_04354_),
    .ZN(_04359_));
 OAI22_X1 _18038_ (.A1(_04343_),
    .A2(_03065_),
    .B1(_03077_),
    .B2(_04325_),
    .ZN(_04360_));
 NOR2_X1 _18039_ (.A1(_04327_),
    .A2(_03095_),
    .ZN(_04361_));
 NOR3_X1 _18040_ (.A1(_04359_),
    .A2(_04360_),
    .A3(_04361_),
    .ZN(_04362_));
 NOR2_X2 _18041_ (.A1(_04314_),
    .A2(_04362_),
    .ZN(net434));
 OAI22_X1 _18042_ (.A1(_04331_),
    .A2(_03102_),
    .B1(_03106_),
    .B2(_04323_),
    .ZN(_04363_));
 OAI22_X1 _18043_ (.A1(_04317_),
    .A2(_03111_),
    .B1(_03115_),
    .B2(_04335_),
    .ZN(_04364_));
 NOR2_X1 _18044_ (.A1(_04363_),
    .A2(_04364_),
    .ZN(_04365_));
 NAND2_X1 _18045_ (.A1(_06977_),
    .A2(_03132_),
    .ZN(_04366_));
 AOI21_X2 _18046_ (.A(_04330_),
    .B1(_04365_),
    .B2(_04366_),
    .ZN(net435));
 OAI22_X2 _18047_ (.A1(_04317_),
    .A2(_03137_),
    .B1(_03141_),
    .B2(_04323_),
    .ZN(_04367_));
 OAI22_X2 _18048_ (.A1(_04331_),
    .A2(_03147_),
    .B1(_03151_),
    .B2(_04335_),
    .ZN(_04368_));
 NOR2_X2 _18049_ (.A1(_04367_),
    .A2(_04368_),
    .ZN(_04369_));
 NAND2_X1 _18050_ (.A1(_06977_),
    .A2(_03168_),
    .ZN(_04370_));
 AOI21_X4 _18051_ (.A(_04330_),
    .B1(_04369_),
    .B2(_04370_),
    .ZN(net436));
 OAI22_X1 _18052_ (.A1(_04353_),
    .A2(_03173_),
    .B1(_03183_),
    .B2(_04343_),
    .ZN(_04371_));
 CLKBUF_X3 _18053_ (.A(_04324_),
    .Z(_04372_));
 OAI22_X1 _18054_ (.A1(_04345_),
    .A2(_03178_),
    .B1(_03188_),
    .B2(_04372_),
    .ZN(_04373_));
 NOR2_X1 _18055_ (.A1(_04327_),
    .A2(_03209_),
    .ZN(_04374_));
 NOR3_X1 _18056_ (.A1(_04371_),
    .A2(_04373_),
    .A3(_04374_),
    .ZN(_04375_));
 NOR2_X1 _18057_ (.A1(_04314_),
    .A2(_04375_),
    .ZN(net437));
 BUF_X4 _18058_ (.A(_04324_),
    .Z(_04376_));
 OAI22_X2 _18059_ (.A1(_04376_),
    .A2(_03216_),
    .B1(_03220_),
    .B2(_04343_),
    .ZN(_04377_));
 OAI22_X2 _18060_ (.A1(_04332_),
    .A2(_03228_),
    .B1(_03234_),
    .B2(_04318_),
    .ZN(_04378_));
 NOR2_X1 _18061_ (.A1(_04327_),
    .A2(_03253_),
    .ZN(_04379_));
 NOR3_X2 _18062_ (.A1(_04377_),
    .A2(_04378_),
    .A3(_04379_),
    .ZN(_04380_));
 NOR2_X2 _18063_ (.A1(_04314_),
    .A2(_04380_),
    .ZN(net438));
 OAI22_X1 _18064_ (.A1(_04353_),
    .A2(_03259_),
    .B1(_03264_),
    .B2(_04354_),
    .ZN(_04381_));
 OAI22_X1 _18065_ (.A1(_04343_),
    .A2(_03269_),
    .B1(_03273_),
    .B2(_04372_),
    .ZN(_04382_));
 NOR2_X1 _18066_ (.A1(_04327_),
    .A2(_03294_),
    .ZN(_04383_));
 NOR3_X1 _18067_ (.A1(_04381_),
    .A2(_04382_),
    .A3(_04383_),
    .ZN(_04384_));
 NOR2_X1 _18068_ (.A1(_04314_),
    .A2(_04384_),
    .ZN(net439));
 OAI22_X1 _18069_ (.A1(_04331_),
    .A2(_03301_),
    .B1(_03305_),
    .B2(_04323_),
    .ZN(_04385_));
 OAI22_X1 _18070_ (.A1(_04317_),
    .A2(_03310_),
    .B1(_03314_),
    .B2(_04335_),
    .ZN(_04386_));
 NOR2_X1 _18071_ (.A1(_04385_),
    .A2(_04386_),
    .ZN(_04387_));
 NAND2_X1 _18072_ (.A1(_06977_),
    .A2(_03331_),
    .ZN(_04388_));
 AOI21_X2 _18073_ (.A(_04330_),
    .B1(_04387_),
    .B2(_04388_),
    .ZN(net440));
 BUF_X4 _18074_ (.A(_04321_),
    .Z(_04389_));
 OAI22_X1 _18075_ (.A1(_04353_),
    .A2(_03336_),
    .B1(_03346_),
    .B2(_04389_),
    .ZN(_04390_));
 OAI22_X1 _18076_ (.A1(_04345_),
    .A2(_03341_),
    .B1(_03350_),
    .B2(_04372_),
    .ZN(_04391_));
 NOR2_X1 _18077_ (.A1(_04327_),
    .A2(_03369_),
    .ZN(_04392_));
 NOR3_X1 _18078_ (.A1(_04390_),
    .A2(_04391_),
    .A3(_04392_),
    .ZN(_04393_));
 NOR2_X1 _18079_ (.A1(_04314_),
    .A2(_04393_),
    .ZN(net441));
 INV_X4 _18080_ (.A(_04315_),
    .ZN(_04394_));
 BUF_X4 _18081_ (.A(_05593_),
    .Z(_04395_));
 AOI22_X1 _18082_ (.A1(_04394_),
    .A2(_05775_),
    .B1(_06080_),
    .B2(_04395_),
    .ZN(_04396_));
 OAI221_X1 _18083_ (.A(_04396_),
    .B1(_03374_),
    .B2(_04389_),
    .C1(_04325_),
    .C2(_02494_),
    .ZN(_04397_));
 BUF_X4 _18084_ (.A(_06916_),
    .Z(_04398_));
 AOI21_X1 _18085_ (.A(_04397_),
    .B1(_07132_),
    .B2(_04398_),
    .ZN(_04399_));
 NOR2_X1 _18086_ (.A1(_04314_),
    .A2(_04399_),
    .ZN(net442));
 INV_X4 _18087_ (.A(_00066_),
    .ZN(_04400_));
 BUF_X4 _18088_ (.A(_04400_),
    .Z(_04401_));
 INV_X1 _18089_ (.A(_04321_),
    .ZN(_04402_));
 BUF_X4 _18090_ (.A(_04402_),
    .Z(_04403_));
 AOI22_X1 _18091_ (.A1(_04401_),
    .A2(_05849_),
    .B1(_05796_),
    .B2(_04403_),
    .ZN(_04404_));
 OAI221_X1 _18092_ (.A(_04404_),
    .B1(_03383_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_03382_),
    .ZN(_04405_));
 AOI21_X1 _18093_ (.A(_04405_),
    .B1(_07156_),
    .B2(_04398_),
    .ZN(_04406_));
 NOR2_X1 _18094_ (.A1(_04314_),
    .A2(_04406_),
    .ZN(net443));
 BUF_X4 _18095_ (.A(_04313_),
    .Z(_04407_));
 AOI22_X1 _18096_ (.A1(_04401_),
    .A2(_05839_),
    .B1(_05799_),
    .B2(_04403_),
    .ZN(_04408_));
 OAI221_X1 _18097_ (.A(_04408_),
    .B1(_03389_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_03388_),
    .ZN(_04409_));
 AOI21_X1 _18098_ (.A(_04409_),
    .B1(_05956_),
    .B2(_04398_),
    .ZN(_04410_));
 NOR2_X1 _18099_ (.A1(_04407_),
    .A2(_04410_),
    .ZN(net444));
 AOI22_X1 _18100_ (.A1(_04401_),
    .A2(_05829_),
    .B1(_05802_),
    .B2(_04402_),
    .ZN(_04411_));
 OAI221_X1 _18101_ (.A(_04411_),
    .B1(_03395_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_03393_),
    .ZN(_04412_));
 AOI21_X1 _18102_ (.A(_04412_),
    .B1(_05902_),
    .B2(_04398_),
    .ZN(_04413_));
 NOR2_X1 _18103_ (.A1(_04407_),
    .A2(_04413_),
    .ZN(net445));
 AOI22_X1 _18104_ (.A1(_04401_),
    .A2(_05832_),
    .B1(_05792_),
    .B2(_04402_),
    .ZN(_04414_));
 OAI221_X1 _18105_ (.A(_04414_),
    .B1(_03400_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_03399_),
    .ZN(_04415_));
 AOI21_X1 _18106_ (.A(_04415_),
    .B1(_03403_),
    .B2(_04398_),
    .ZN(_04416_));
 NOR2_X1 _18107_ (.A1(_04407_),
    .A2(_04416_),
    .ZN(net446));
 AOI22_X1 _18108_ (.A1(_04401_),
    .A2(_05836_),
    .B1(_05809_),
    .B2(_04402_),
    .ZN(_04417_));
 OAI221_X1 _18109_ (.A(_04417_),
    .B1(_07233_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_07196_),
    .ZN(_04418_));
 AOI21_X1 _18110_ (.A(_04418_),
    .B1(_05972_),
    .B2(_04398_),
    .ZN(_04419_));
 NOR2_X1 _18111_ (.A1(_04407_),
    .A2(_04419_),
    .ZN(net447));
 AOI22_X1 _18112_ (.A1(_04401_),
    .A2(_05843_),
    .B1(_05806_),
    .B2(_04402_),
    .ZN(_04420_));
 OAI221_X1 _18113_ (.A(_04420_),
    .B1(_07229_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_07192_),
    .ZN(_04421_));
 AOI21_X1 _18114_ (.A(_04421_),
    .B1(_06008_),
    .B2(_04398_),
    .ZN(_04422_));
 NOR2_X1 _18115_ (.A1(_04407_),
    .A2(_04422_),
    .ZN(net448));
 AOI22_X2 _18116_ (.A1(_04394_),
    .A2(_05778_),
    .B1(_06071_),
    .B2(_04395_),
    .ZN(_04423_));
 OAI221_X2 _18117_ (.A(_04423_),
    .B1(_03412_),
    .B2(_04389_),
    .C1(_04325_),
    .C2(_07105_),
    .ZN(_04424_));
 AOI21_X1 _18118_ (.A(_04424_),
    .B1(_05993_),
    .B2(_04398_),
    .ZN(_04425_));
 NOR2_X1 _18119_ (.A1(_04407_),
    .A2(_04425_),
    .ZN(net449));
 OAI22_X1 _18120_ (.A1(_04353_),
    .A2(_03418_),
    .B1(_03422_),
    .B2(_04389_),
    .ZN(_04426_));
 OAI22_X1 _18121_ (.A1(_04345_),
    .A2(_03428_),
    .B1(_03432_),
    .B2(_04372_),
    .ZN(_04427_));
 NOR2_X1 _18122_ (.A1(_04327_),
    .A2(_03450_),
    .ZN(_04428_));
 NOR3_X1 _18123_ (.A1(_04426_),
    .A2(_04427_),
    .A3(_04428_),
    .ZN(_04429_));
 NOR2_X1 _18124_ (.A1(_04407_),
    .A2(_04429_),
    .ZN(net450));
 AOI22_X1 _18125_ (.A1(_04401_),
    .A2(_06524_),
    .B1(_05492_),
    .B2(_04394_),
    .ZN(_04430_));
 OAI221_X1 _18126_ (.A(_04430_),
    .B1(_05274_),
    .B2(_04389_),
    .C1(_04319_),
    .C2(_06099_),
    .ZN(_04431_));
 BUF_X4 _18127_ (.A(_06916_),
    .Z(_04432_));
 AOI21_X1 _18128_ (.A(_04431_),
    .B1(_06179_),
    .B2(_04432_),
    .ZN(_04433_));
 NOR2_X1 _18129_ (.A1(_04407_),
    .A2(_04433_),
    .ZN(net451));
 AOI22_X2 _18130_ (.A1(_04403_),
    .A2(_06514_),
    .B1(_06100_),
    .B2(_05593_),
    .ZN(_04434_));
 OAI221_X2 _18131_ (.A(_04434_),
    .B1(_05376_),
    .B2(_04324_),
    .C1(_04332_),
    .C2(_06789_),
    .ZN(_04435_));
 AOI21_X2 _18132_ (.A(_04435_),
    .B1(_06146_),
    .B2(_04432_),
    .ZN(_04436_));
 NOR2_X2 _18133_ (.A1(_04407_),
    .A2(_04436_),
    .ZN(net452));
 AOI22_X1 _18134_ (.A1(_04401_),
    .A2(_05370_),
    .B1(_05500_),
    .B2(_04394_),
    .ZN(_04437_));
 OAI221_X1 _18135_ (.A(_04437_),
    .B1(_06513_),
    .B2(_04322_),
    .C1(_04319_),
    .C2(_06098_),
    .ZN(_04438_));
 AOI21_X1 _18136_ (.A(_04438_),
    .B1(_06163_),
    .B2(_04432_),
    .ZN(_04439_));
 NOR2_X1 _18137_ (.A1(_04407_),
    .A2(_04439_),
    .ZN(net453));
 BUF_X4 _18138_ (.A(_04313_),
    .Z(_04440_));
 OAI22_X1 _18139_ (.A1(_04353_),
    .A2(_03465_),
    .B1(_03471_),
    .B2(_04354_),
    .ZN(_04441_));
 OAI22_X1 _18140_ (.A1(_04343_),
    .A2(_03476_),
    .B1(_03480_),
    .B2(_04372_),
    .ZN(_04442_));
 NOR2_X1 _18141_ (.A1(_04327_),
    .A2(_03498_),
    .ZN(_04443_));
 NOR3_X1 _18142_ (.A1(_04441_),
    .A2(_04442_),
    .A3(_04443_),
    .ZN(_04444_));
 NOR2_X1 _18143_ (.A1(_04440_),
    .A2(_04444_),
    .ZN(net454));
 AOI22_X1 _18144_ (.A1(_04395_),
    .A2(_10225_),
    .B1(_10321_),
    .B2(_04400_),
    .ZN(_04445_));
 INV_X1 _18145_ (.A(_10348_),
    .ZN(_04446_));
 OAI221_X1 _18146_ (.A(_04445_),
    .B1(_03502_),
    .B2(_04322_),
    .C1(_04332_),
    .C2(_04446_),
    .ZN(_04447_));
 AOI21_X1 _18147_ (.A(_04447_),
    .B1(_10417_),
    .B2(_04432_),
    .ZN(_04448_));
 NOR2_X2 _18148_ (.A1(_04440_),
    .A2(_04448_),
    .ZN(net455));
 OAI22_X2 _18149_ (.A1(_04315_),
    .A2(_10351_),
    .B1(_10255_),
    .B2(_04321_),
    .ZN(_04449_));
 INV_X1 _18150_ (.A(_10221_),
    .ZN(_04450_));
 AOI221_X2 _18151_ (.A(_04449_),
    .B1(net694),
    .B2(_04400_),
    .C1(_04395_),
    .C2(_04450_),
    .ZN(_04451_));
 NAND2_X1 _18152_ (.A1(_06977_),
    .A2(_07676_),
    .ZN(_04452_));
 AOI21_X2 _18153_ (.A(_04330_),
    .B1(_04451_),
    .B2(_04452_),
    .ZN(net456));
 BUF_X8 _18154_ (.A(_04313_),
    .Z(_04453_));
 OAI22_X2 _18155_ (.A1(_04322_),
    .A2(_10261_),
    .B1(_10357_),
    .B2(_04315_),
    .ZN(_04454_));
 AOI221_X2 _18156_ (.A(_04454_),
    .B1(_04175_),
    .B2(_04400_),
    .C1(_04395_),
    .C2(_07434_),
    .ZN(_04455_));
 NAND2_X1 _18157_ (.A1(_06977_),
    .A2(_07661_),
    .ZN(_04456_));
 AOI21_X2 _18158_ (.A(_04453_),
    .B1(_04455_),
    .B2(_04456_),
    .ZN(net457));
 AOI22_X1 _18159_ (.A1(_04395_),
    .A2(net742),
    .B1(_07305_),
    .B2(_04394_),
    .ZN(_04457_));
 OAI221_X1 _18160_ (.A(_04457_),
    .B1(_10258_),
    .B2(_04322_),
    .C1(_04325_),
    .C2(_10312_),
    .ZN(_04458_));
 AOI21_X1 _18161_ (.A(_04458_),
    .B1(_07409_),
    .B2(_04432_),
    .ZN(_04459_));
 NOR2_X2 _18162_ (.A1(_04440_),
    .A2(_04459_),
    .ZN(net458));
 AOI22_X1 _18163_ (.A1(_04403_),
    .A2(_07282_),
    .B1(net673),
    .B2(_05593_),
    .ZN(_04460_));
 BUF_X4 _18164_ (.A(_04315_),
    .Z(_04461_));
 OAI221_X1 _18165_ (.A(_04460_),
    .B1(net697),
    .B2(_04324_),
    .C1(_04461_),
    .C2(_10369_),
    .ZN(_04462_));
 AOI21_X1 _18166_ (.A(_04462_),
    .B1(_07646_),
    .B2(_04432_),
    .ZN(_04463_));
 NOR2_X2 _18167_ (.A1(_04440_),
    .A2(_04463_),
    .ZN(net459));
 OAI22_X2 _18168_ (.A1(_04322_),
    .A2(_10270_),
    .B1(_10209_),
    .B2(_05592_),
    .ZN(_04464_));
 AOI221_X2 _18169_ (.A(_04464_),
    .B1(net665),
    .B2(_04400_),
    .C1(_04394_),
    .C2(_03522_),
    .ZN(_04465_));
 NAND2_X1 _18170_ (.A1(_06977_),
    .A2(_07631_),
    .ZN(_04466_));
 AOI21_X2 _18171_ (.A(_04453_),
    .B1(_04465_),
    .B2(_04466_),
    .ZN(net460));
 OAI22_X1 _18172_ (.A1(_04331_),
    .A2(_03530_),
    .B1(_03534_),
    .B2(_04389_),
    .ZN(_04467_));
 OAI22_X1 _18173_ (.A1(_04332_),
    .A2(_03539_),
    .B1(_03543_),
    .B2(_04372_),
    .ZN(_04468_));
 CLKBUF_X3 _18174_ (.A(_07082_),
    .Z(_04469_));
 NOR2_X1 _18175_ (.A1(_04469_),
    .A2(_03562_),
    .ZN(_04470_));
 NOR3_X1 _18176_ (.A1(_04467_),
    .A2(_04468_),
    .A3(_04470_),
    .ZN(_04471_));
 NOR2_X2 _18177_ (.A1(_04440_),
    .A2(_04471_),
    .ZN(net461));
 AOI22_X1 _18178_ (.A1(_04403_),
    .A2(_07473_),
    .B1(_07506_),
    .B2(_04400_),
    .ZN(_04472_));
 OAI221_X1 _18179_ (.A(_04472_),
    .B1(_10363_),
    .B2(_04316_),
    .C1(_04319_),
    .C2(_10206_),
    .ZN(_04473_));
 AOI21_X1 _18180_ (.A(_04473_),
    .B1(_07616_),
    .B2(_04432_),
    .ZN(_04474_));
 NOR2_X1 _18181_ (.A1(_04440_),
    .A2(_04474_),
    .ZN(net462));
 OAI22_X1 _18182_ (.A1(_04334_),
    .A2(net640),
    .B1(net713),
    .B2(_04332_),
    .ZN(_04475_));
 OAI22_X1 _18183_ (.A1(_04331_),
    .A2(net650),
    .B1(net632),
    .B2(_04335_),
    .ZN(_04476_));
 NOR2_X1 _18184_ (.A1(_04475_),
    .A2(_04476_),
    .ZN(_04477_));
 CLKBUF_X3 _18185_ (.A(_06916_),
    .Z(_04478_));
 NAND2_X1 _18186_ (.A1(_04478_),
    .A2(_07394_),
    .ZN(_04479_));
 AOI21_X2 _18187_ (.A(_04453_),
    .B1(_04477_),
    .B2(_04479_),
    .ZN(net463));
 AOI22_X1 _18188_ (.A1(_04403_),
    .A2(_10249_),
    .B1(_10345_),
    .B2(_04394_),
    .ZN(_04480_));
 AOI22_X1 _18189_ (.A1(_04395_),
    .A2(_10179_),
    .B1(_10276_),
    .B2(_04401_),
    .ZN(_04481_));
 NAND2_X1 _18190_ (.A1(_04480_),
    .A2(_04481_),
    .ZN(_04482_));
 AOI21_X1 _18191_ (.A(_04482_),
    .B1(_10372_),
    .B2(_04432_),
    .ZN(_04483_));
 NOR2_X2 _18192_ (.A1(_04440_),
    .A2(_04483_),
    .ZN(net464));
 OAI22_X2 _18193_ (.A1(_05592_),
    .A2(net643),
    .B1(_10246_),
    .B2(_04321_),
    .ZN(_04484_));
 AOI221_X2 _18194_ (.A(_04484_),
    .B1(_03578_),
    .B2(_04400_),
    .C1(_04394_),
    .C2(_03577_),
    .ZN(_04485_));
 NAND2_X1 _18195_ (.A1(_04478_),
    .A2(_07556_),
    .ZN(_04486_));
 AOI21_X4 _18196_ (.A(_04453_),
    .B1(_04485_),
    .B2(_04486_),
    .ZN(net465));
 OAI22_X2 _18197_ (.A1(_05592_),
    .A2(net645),
    .B1(net723),
    .B2(_04315_),
    .ZN(_04487_));
 AOI221_X2 _18198_ (.A(_04487_),
    .B1(_03583_),
    .B2(_04403_),
    .C1(_04401_),
    .C2(net690),
    .ZN(_04488_));
 NAND2_X1 _18199_ (.A1(_04478_),
    .A2(_07571_),
    .ZN(_04489_));
 AOI21_X4 _18200_ (.A(_04453_),
    .B1(_04488_),
    .B2(_04489_),
    .ZN(net466));
 OAI22_X2 _18201_ (.A1(_04322_),
    .A2(_10240_),
    .B1(_10336_),
    .B2(_04315_),
    .ZN(_04490_));
 AOI221_X2 _18202_ (.A(_04490_),
    .B1(_04211_),
    .B2(_04400_),
    .C1(_04395_),
    .C2(_04210_),
    .ZN(_04491_));
 NAND2_X1 _18203_ (.A1(_04478_),
    .A2(_07342_),
    .ZN(_04492_));
 AOI21_X4 _18204_ (.A(_04453_),
    .B1(_04491_),
    .B2(_04492_),
    .ZN(net467));
 OAI22_X2 _18205_ (.A1(_05592_),
    .A2(net647),
    .B1(_10288_),
    .B2(_04324_),
    .ZN(_04493_));
 AOI221_X2 _18206_ (.A(_04493_),
    .B1(_03590_),
    .B2(_04403_),
    .C1(_04394_),
    .C2(net652),
    .ZN(_04494_));
 NAND2_X1 _18207_ (.A1(_04478_),
    .A2(_07376_),
    .ZN(_04495_));
 AOI21_X2 _18208_ (.A(_04453_),
    .B1(_04494_),
    .B2(_04495_),
    .ZN(net468));
 OAI22_X2 _18209_ (.A1(_04315_),
    .A2(net703),
    .B1(net732),
    .B2(_04321_),
    .ZN(_04496_));
 AOI221_X2 _18210_ (.A(_04496_),
    .B1(_07489_),
    .B2(_04400_),
    .C1(_04395_),
    .C2(_04220_),
    .ZN(_04497_));
 NAND2_X1 _18211_ (.A1(_04478_),
    .A2(_07361_),
    .ZN(_04498_));
 AOI21_X4 _18212_ (.A(_04453_),
    .B1(_04497_),
    .B2(_04498_),
    .ZN(net469));
 OAI22_X2 _18213_ (.A1(_04322_),
    .A2(net750),
    .B1(_10294_),
    .B2(_04324_),
    .ZN(_04499_));
 AOI221_X2 _18214_ (.A(_04499_),
    .B1(_03599_),
    .B2(_04394_),
    .C1(_04395_),
    .C2(net752),
    .ZN(_04500_));
 NAND2_X1 _18215_ (.A1(_04478_),
    .A2(_07601_),
    .ZN(_04501_));
 AOI21_X2 _18216_ (.A(_04453_),
    .B1(_04500_),
    .B2(_04501_),
    .ZN(net470));
 OAI22_X1 _18217_ (.A1(_04334_),
    .A2(_10228_),
    .B1(net671),
    .B2(_04332_),
    .ZN(_04502_));
 OAI22_X1 _18218_ (.A1(_04331_),
    .A2(_10191_),
    .B1(_10297_),
    .B2(_04325_),
    .ZN(_04503_));
 NOR2_X1 _18219_ (.A1(_04502_),
    .A2(_04503_),
    .ZN(_04504_));
 NAND2_X1 _18220_ (.A1(_04478_),
    .A2(_07586_),
    .ZN(_04505_));
 AOI21_X2 _18221_ (.A(_04453_),
    .B1(_04504_),
    .B2(_04505_),
    .ZN(net471));
 OAI22_X1 _18222_ (.A1(_04331_),
    .A2(_03610_),
    .B1(_03614_),
    .B2(_04323_),
    .ZN(_04506_));
 OAI22_X1 _18223_ (.A1(_04317_),
    .A2(_03619_),
    .B1(_03623_),
    .B2(_04325_),
    .ZN(_04507_));
 NOR2_X1 _18224_ (.A1(_04506_),
    .A2(_04507_),
    .ZN(_04508_));
 NAND2_X1 _18225_ (.A1(_04478_),
    .A2(_03640_),
    .ZN(_04509_));
 AOI21_X2 _18226_ (.A(_04313_),
    .B1(_04508_),
    .B2(_04509_),
    .ZN(net472));
 OAI22_X1 _18227_ (.A1(_04334_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(_04354_),
    .ZN(_04510_));
 OAI22_X1 _18228_ (.A1(_04376_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_04461_),
    .ZN(_04511_));
 NOR2_X1 _18229_ (.A1(_04469_),
    .A2(_03655_),
    .ZN(_04512_));
 NOR3_X1 _18230_ (.A1(_04510_),
    .A2(_04511_),
    .A3(_04512_),
    .ZN(_04513_));
 NOR2_X1 _18231_ (.A1(_04440_),
    .A2(_04513_),
    .ZN(net473));
 AOI22_X1 _18232_ (.A1(_04403_),
    .A2(_05189_),
    .B1(_05649_),
    .B2(_05593_),
    .ZN(_04514_));
 OAI221_X1 _18233_ (.A(_04514_),
    .B1(_03660_),
    .B2(_04324_),
    .C1(_04461_),
    .C2(_03662_),
    .ZN(_04515_));
 AOI21_X1 _18234_ (.A(_04515_),
    .B1(_06249_),
    .B2(_04432_),
    .ZN(_04516_));
 NOR2_X2 _18235_ (.A1(_04440_),
    .A2(_04516_),
    .ZN(net474));
 OAI22_X1 _18236_ (.A1(_04334_),
    .A2(_03666_),
    .B1(_03669_),
    .B2(_04354_),
    .ZN(_04517_));
 OAI22_X1 _18237_ (.A1(_04376_),
    .A2(_03672_),
    .B1(_03674_),
    .B2(_04461_),
    .ZN(_04518_));
 NOR2_X1 _18238_ (.A1(_04469_),
    .A2(_03677_),
    .ZN(_04519_));
 NOR3_X1 _18239_ (.A1(_04517_),
    .A2(_04518_),
    .A3(_04519_),
    .ZN(_04520_));
 NOR2_X1 _18240_ (.A1(_04440_),
    .A2(_04520_),
    .ZN(net475));
 OAI22_X2 _18241_ (.A1(_04334_),
    .A2(_03681_),
    .B1(_03686_),
    .B2(_04376_),
    .ZN(_04521_));
 OAI22_X2 _18242_ (.A1(_04317_),
    .A2(_03683_),
    .B1(_03689_),
    .B2(_04345_),
    .ZN(_04522_));
 NOR2_X2 _18243_ (.A1(_04521_),
    .A2(_04522_),
    .ZN(_04523_));
 NAND2_X1 _18244_ (.A1(_04478_),
    .A2(_06330_),
    .ZN(_04524_));
 AOI21_X4 _18245_ (.A(_04313_),
    .B1(_04523_),
    .B2(_04524_),
    .ZN(net476));
 BUF_X4 _18246_ (.A(_04313_),
    .Z(_04525_));
 OAI22_X2 _18247_ (.A1(_04334_),
    .A2(_03696_),
    .B1(_03699_),
    .B2(_04354_),
    .ZN(_04526_));
 OAI22_X2 _18248_ (.A1(_04376_),
    .A2(_03702_),
    .B1(_03704_),
    .B2(_04461_),
    .ZN(_04527_));
 NOR2_X1 _18249_ (.A1(_04469_),
    .A2(_03707_),
    .ZN(_04528_));
 NOR3_X2 _18250_ (.A1(_04526_),
    .A2(_04527_),
    .A3(_04528_),
    .ZN(_04529_));
 NOR2_X4 _18251_ (.A1(_04525_),
    .A2(_04529_),
    .ZN(net477));
 OAI22_X1 _18252_ (.A1(_04323_),
    .A2(_03717_),
    .B1(_03720_),
    .B2(_04354_),
    .ZN(_04530_));
 OAI22_X1 _18253_ (.A1(_04335_),
    .A2(_03712_),
    .B1(_03714_),
    .B2(_04461_),
    .ZN(_04531_));
 NOR2_X1 _18254_ (.A1(_04469_),
    .A2(_03723_),
    .ZN(_04532_));
 NOR3_X1 _18255_ (.A1(_04530_),
    .A2(_04531_),
    .A3(_04532_),
    .ZN(_04533_));
 NOR2_X2 _18256_ (.A1(_04525_),
    .A2(_04533_),
    .ZN(net478));
 OAI22_X1 _18257_ (.A1(_04317_),
    .A2(_03727_),
    .B1(_03730_),
    .B2(_04345_),
    .ZN(_04534_));
 OAI22_X1 _18258_ (.A1(_04334_),
    .A2(_03733_),
    .B1(_03735_),
    .B2(_04325_),
    .ZN(_04535_));
 NOR2_X1 _18259_ (.A1(_04534_),
    .A2(_04535_),
    .ZN(_04536_));
 NAND2_X1 _18260_ (.A1(_04398_),
    .A2(_03738_),
    .ZN(_04537_));
 AOI21_X2 _18261_ (.A(_04313_),
    .B1(_04536_),
    .B2(_04537_),
    .ZN(net479));
 OAI22_X1 _18262_ (.A1(_04376_),
    .A2(_03741_),
    .B1(_03743_),
    .B2(_04461_),
    .ZN(_04538_));
 OAI22_X1 _18263_ (.A1(_04343_),
    .A2(_03746_),
    .B1(_03749_),
    .B2(_04318_),
    .ZN(_04539_));
 NOR2_X1 _18264_ (.A1(_04469_),
    .A2(_03752_),
    .ZN(_04540_));
 NOR3_X1 _18265_ (.A1(_04538_),
    .A2(_04539_),
    .A3(_04540_),
    .ZN(_04541_));
 NOR2_X2 _18266_ (.A1(_04525_),
    .A2(_04541_),
    .ZN(net480));
 OAI22_X1 _18267_ (.A1(_04323_),
    .A2(_03756_),
    .B1(_03759_),
    .B2(_04354_),
    .ZN(_04542_));
 OAI22_X1 _18268_ (.A1(_04335_),
    .A2(_03762_),
    .B1(_03764_),
    .B2(_04316_),
    .ZN(_04543_));
 NOR2_X1 _18269_ (.A1(_04469_),
    .A2(_03767_),
    .ZN(_04544_));
 NOR3_X1 _18270_ (.A1(_04542_),
    .A2(_04543_),
    .A3(_04544_),
    .ZN(_04545_));
 NOR2_X2 _18271_ (.A1(_04525_),
    .A2(_04545_),
    .ZN(net481));
 OAI22_X1 _18272_ (.A1(_04376_),
    .A2(_03771_),
    .B1(_03773_),
    .B2(_04461_),
    .ZN(_04546_));
 OAI22_X1 _18273_ (.A1(_04343_),
    .A2(_03776_),
    .B1(_03779_),
    .B2(_04318_),
    .ZN(_04547_));
 NOR2_X1 _18274_ (.A1(_04469_),
    .A2(_03782_),
    .ZN(_04548_));
 NOR3_X1 _18275_ (.A1(_04546_),
    .A2(_04547_),
    .A3(_04548_),
    .ZN(_04549_));
 NOR2_X2 _18276_ (.A1(_04525_),
    .A2(_04549_),
    .ZN(net482));
 OAI22_X1 _18277_ (.A1(_04353_),
    .A2(_03788_),
    .B1(_03798_),
    .B2(_04389_),
    .ZN(_04550_));
 OAI22_X1 _18278_ (.A1(_04345_),
    .A2(_03793_),
    .B1(_03802_),
    .B2(_04372_),
    .ZN(_04551_));
 NOR2_X1 _18279_ (.A1(_04469_),
    .A2(_03820_),
    .ZN(_04552_));
 NOR3_X1 _18280_ (.A1(_04550_),
    .A2(_04551_),
    .A3(_04552_),
    .ZN(_04553_));
 NOR2_X2 _18281_ (.A1(_04525_),
    .A2(_04553_),
    .ZN(net483));
 AOI22_X1 _18282_ (.A1(_04403_),
    .A2(_05194_),
    .B1(_05639_),
    .B2(_05593_),
    .ZN(_04554_));
 OAI221_X1 _18283_ (.A(_04554_),
    .B1(_04282_),
    .B2(_04324_),
    .C1(_04461_),
    .C2(_04281_),
    .ZN(_04555_));
 AOI21_X1 _18284_ (.A(_04555_),
    .B1(_03827_),
    .B2(_04432_),
    .ZN(_04556_));
 NOR2_X1 _18285_ (.A1(_04525_),
    .A2(_04556_),
    .ZN(net484));
 OAI22_X1 _18286_ (.A1(_04376_),
    .A2(_03836_),
    .B1(_03833_),
    .B2(_04461_),
    .ZN(_04557_));
 OAI22_X1 _18287_ (.A1(_04343_),
    .A2(_03831_),
    .B1(_03839_),
    .B2(_04318_),
    .ZN(_04558_));
 NOR2_X1 _18288_ (.A1(_04469_),
    .A2(_03849_),
    .ZN(_04559_));
 NOR3_X1 _18289_ (.A1(_04557_),
    .A2(_04558_),
    .A3(_04559_),
    .ZN(_04560_));
 NOR2_X2 _18290_ (.A1(_04525_),
    .A2(_04560_),
    .ZN(net485));
 OAI22_X1 _18291_ (.A1(_04334_),
    .A2(_03853_),
    .B1(_03855_),
    .B2(_04376_),
    .ZN(_04561_));
 OAI22_X1 _18292_ (.A1(_04317_),
    .A2(_03858_),
    .B1(_03861_),
    .B2(_04345_),
    .ZN(_04562_));
 NOR2_X1 _18293_ (.A1(_04561_),
    .A2(_04562_),
    .ZN(_04563_));
 NAND2_X1 _18294_ (.A1(_04398_),
    .A2(_03864_),
    .ZN(_04564_));
 AOI21_X2 _18295_ (.A(_04313_),
    .B1(_04563_),
    .B2(_04564_),
    .ZN(net486));
 OAI22_X1 _18296_ (.A1(_04323_),
    .A2(_03867_),
    .B1(_03875_),
    .B2(_04354_),
    .ZN(_04565_));
 OAI22_X1 _18297_ (.A1(_04335_),
    .A2(_03872_),
    .B1(_03869_),
    .B2(_04316_),
    .ZN(_04566_));
 NOR2_X1 _18298_ (.A1(_07082_),
    .A2(_06229_),
    .ZN(_04567_));
 NOR3_X1 _18299_ (.A1(_04565_),
    .A2(_04566_),
    .A3(_04567_),
    .ZN(_04568_));
 NOR2_X2 _18300_ (.A1(_04525_),
    .A2(_04568_),
    .ZN(net487));
 OAI22_X1 _18301_ (.A1(_04353_),
    .A2(_03882_),
    .B1(_03892_),
    .B2(_04389_),
    .ZN(_04569_));
 OAI22_X1 _18302_ (.A1(_04345_),
    .A2(_03887_),
    .B1(_03896_),
    .B2(_04372_),
    .ZN(_04570_));
 NOR2_X1 _18303_ (.A1(_07082_),
    .A2(_03914_),
    .ZN(_04571_));
 NOR3_X1 _18304_ (.A1(_04569_),
    .A2(_04570_),
    .A3(_04571_),
    .ZN(_04572_));
 NOR2_X2 _18305_ (.A1(_04525_),
    .A2(_04572_),
    .ZN(net488));
 OAI22_X1 _18306_ (.A1(_04353_),
    .A2(_03920_),
    .B1(_03925_),
    .B2(_04318_),
    .ZN(_04573_));
 OAI22_X1 _18307_ (.A1(_04343_),
    .A2(_03930_),
    .B1(_03934_),
    .B2(_04372_),
    .ZN(_04574_));
 NOR2_X1 _18308_ (.A1(_07082_),
    .A2(_03952_),
    .ZN(_04575_));
 NOR3_X1 _18309_ (.A1(_04573_),
    .A2(_04574_),
    .A3(_04575_),
    .ZN(_04576_));
 NOR2_X2 _18310_ (.A1(_04330_),
    .A2(_04576_),
    .ZN(net489));
 OAI22_X1 _18311_ (.A1(_04376_),
    .A2(_03958_),
    .B1(_03962_),
    .B2(_04389_),
    .ZN(_04577_));
 OAI22_X1 _18312_ (.A1(_04332_),
    .A2(_03967_),
    .B1(_03972_),
    .B2(_04318_),
    .ZN(_04578_));
 NOR2_X1 _18313_ (.A1(_07082_),
    .A2(_03990_),
    .ZN(_04579_));
 NOR3_X1 _18314_ (.A1(_04577_),
    .A2(_04578_),
    .A3(_04579_),
    .ZN(_04580_));
 NOR2_X2 _18315_ (.A1(_04330_),
    .A2(_04580_),
    .ZN(net490));
 OAI22_X1 _18316_ (.A1(_04345_),
    .A2(_03997_),
    .B1(_04001_),
    .B2(_04389_),
    .ZN(_04581_));
 OAI22_X1 _18317_ (.A1(_04332_),
    .A2(_04006_),
    .B1(_04010_),
    .B2(_04372_),
    .ZN(_04582_));
 NOR2_X1 _18318_ (.A1(_07082_),
    .A2(_04028_),
    .ZN(_04583_));
 NOR3_X1 _18319_ (.A1(_04581_),
    .A2(_04582_),
    .A3(_04583_),
    .ZN(_04584_));
 NOR2_X2 _18320_ (.A1(_04330_),
    .A2(_04584_),
    .ZN(net491));
 BUF_X8 _18321_ (.A(_05334_),
    .Z(_04585_));
 BUF_X4 _18322_ (.A(_04585_),
    .Z(_04586_));
 BUF_X4 _18323_ (.A(_00070_),
    .Z(_04587_));
 BUF_X4 _18324_ (.A(_04587_),
    .Z(_04588_));
 BUF_X4 _18325_ (.A(_04588_),
    .Z(_04589_));
 BUF_X4 _18326_ (.A(_00069_),
    .Z(_04590_));
 BUF_X4 _18327_ (.A(_04590_),
    .Z(_04591_));
 BUF_X4 _18328_ (.A(_04591_),
    .Z(_04592_));
 OAI22_X1 _18329_ (.A1(_04589_),
    .A2(_02768_),
    .B1(_02790_),
    .B2(_04592_),
    .ZN(_04593_));
 BUF_X4 _18330_ (.A(_05328_),
    .Z(_04594_));
 BUF_X4 _18331_ (.A(_04594_),
    .Z(_04595_));
 OAI22_X1 _18332_ (.A1(_06860_),
    .A2(_02777_),
    .B1(_02798_),
    .B2(_04595_),
    .ZN(_04596_));
 BUF_X4 _18333_ (.A(_00068_),
    .Z(_04597_));
 CLKBUF_X3 _18334_ (.A(_04597_),
    .Z(_04598_));
 NOR2_X1 _18335_ (.A1(_04598_),
    .A2(_02840_),
    .ZN(_04599_));
 NOR3_X1 _18336_ (.A1(_04593_),
    .A2(_04596_),
    .A3(_04599_),
    .ZN(_04600_));
 NOR2_X2 _18337_ (.A1(_04586_),
    .A2(_04600_),
    .ZN(net492));
 BUF_X4 _18338_ (.A(_04585_),
    .Z(_04601_));
 BUF_X4 _18339_ (.A(_06859_),
    .Z(_04602_));
 BUF_X4 _18340_ (.A(_04588_),
    .Z(_04603_));
 OAI22_X1 _18341_ (.A1(_04602_),
    .A2(_02850_),
    .B1(_02854_),
    .B2(_04603_),
    .ZN(_04604_));
 BUF_X4 _18342_ (.A(_04591_),
    .Z(_04605_));
 BUF_X4 _18343_ (.A(_04594_),
    .Z(_04606_));
 OAI22_X1 _18344_ (.A1(_04605_),
    .A2(_02864_),
    .B1(_02868_),
    .B2(_04606_),
    .ZN(_04607_));
 NOR2_X1 _18345_ (.A1(_04604_),
    .A2(_04607_),
    .ZN(_04608_));
 INV_X1 _18346_ (.A(_04597_),
    .ZN(_04609_));
 BUF_X4 _18347_ (.A(_04609_),
    .Z(_04610_));
 BUF_X4 _18348_ (.A(_04610_),
    .Z(_04611_));
 NAND2_X1 _18349_ (.A1(_04611_),
    .A2(_02896_),
    .ZN(_04612_));
 AOI21_X2 _18350_ (.A(_04601_),
    .B1(_04608_),
    .B2(_04612_),
    .ZN(net493));
 OAI22_X1 _18351_ (.A1(_04605_),
    .A2(_02905_),
    .B1(_02912_),
    .B2(_06860_),
    .ZN(_04613_));
 OAI22_X1 _18352_ (.A1(_04589_),
    .A2(_02901_),
    .B1(_02916_),
    .B2(_04606_),
    .ZN(_04614_));
 NOR2_X1 _18353_ (.A1(_04613_),
    .A2(_04614_),
    .ZN(_04615_));
 NAND2_X1 _18354_ (.A1(_04611_),
    .A2(_02934_),
    .ZN(_04616_));
 AOI21_X2 _18355_ (.A(_04601_),
    .B1(_04615_),
    .B2(_04616_),
    .ZN(net494));
 BUF_X4 _18356_ (.A(_06858_),
    .Z(_04617_));
 OAI22_X2 _18357_ (.A1(_04589_),
    .A2(_02940_),
    .B1(_02946_),
    .B2(_04617_),
    .ZN(_04618_));
 BUF_X4 _18358_ (.A(_04591_),
    .Z(_04619_));
 OAI22_X2 _18359_ (.A1(_04619_),
    .A2(_02952_),
    .B1(_02956_),
    .B2(_04595_),
    .ZN(_04620_));
 NOR2_X1 _18360_ (.A1(_04598_),
    .A2(_02974_),
    .ZN(_04621_));
 NOR3_X2 _18361_ (.A1(_04618_),
    .A2(_04620_),
    .A3(_04621_),
    .ZN(_04622_));
 NOR2_X2 _18362_ (.A1(_04586_),
    .A2(_04622_),
    .ZN(net495));
 OAI22_X1 _18363_ (.A1(_04602_),
    .A2(_02981_),
    .B1(_02985_),
    .B2(_04603_),
    .ZN(_04623_));
 OAI22_X1 _18364_ (.A1(_04605_),
    .A2(_02990_),
    .B1(_02996_),
    .B2(_04606_),
    .ZN(_04624_));
 NOR2_X1 _18365_ (.A1(_04623_),
    .A2(_04624_),
    .ZN(_04625_));
 NAND2_X1 _18366_ (.A1(_04611_),
    .A2(_03013_),
    .ZN(_04626_));
 AOI21_X2 _18367_ (.A(_04601_),
    .B1(_04625_),
    .B2(_04626_),
    .ZN(net496));
 OAI22_X1 _18368_ (.A1(_04589_),
    .A2(_03019_),
    .B1(_03030_),
    .B2(_04592_),
    .ZN(_04627_));
 OAI22_X1 _18369_ (.A1(_06860_),
    .A2(_03024_),
    .B1(_03034_),
    .B2(_04595_),
    .ZN(_04628_));
 NOR2_X1 _18370_ (.A1(_04598_),
    .A2(_03055_),
    .ZN(_04629_));
 NOR3_X1 _18371_ (.A1(_04627_),
    .A2(_04628_),
    .A3(_04629_),
    .ZN(_04630_));
 NOR2_X2 _18372_ (.A1(_04586_),
    .A2(_04630_),
    .ZN(net497));
 OAI22_X1 _18373_ (.A1(_04589_),
    .A2(_03061_),
    .B1(_03065_),
    .B2(_04592_),
    .ZN(_04631_));
 OAI22_X1 _18374_ (.A1(_06860_),
    .A2(_03073_),
    .B1(_03077_),
    .B2(_04595_),
    .ZN(_04632_));
 NOR2_X1 _18375_ (.A1(_04598_),
    .A2(_03095_),
    .ZN(_04633_));
 NOR3_X1 _18376_ (.A1(_04631_),
    .A2(_04632_),
    .A3(_04633_),
    .ZN(_04634_));
 NOR2_X2 _18377_ (.A1(_04586_),
    .A2(_04634_),
    .ZN(net498));
 BUF_X4 _18378_ (.A(_04588_),
    .Z(_04635_));
 OAI22_X1 _18379_ (.A1(_04605_),
    .A2(_03106_),
    .B1(_03111_),
    .B2(_04635_),
    .ZN(_04636_));
 OAI22_X1 _18380_ (.A1(_04602_),
    .A2(_03102_),
    .B1(_03115_),
    .B2(_04606_),
    .ZN(_04637_));
 NOR2_X1 _18381_ (.A1(_04636_),
    .A2(_04637_),
    .ZN(_04638_));
 NAND2_X1 _18382_ (.A1(_04611_),
    .A2(_03132_),
    .ZN(_04639_));
 AOI21_X2 _18383_ (.A(_04601_),
    .B1(_04638_),
    .B2(_04639_),
    .ZN(net499));
 OAI22_X1 _18384_ (.A1(_04589_),
    .A2(_03137_),
    .B1(_03141_),
    .B2(_04619_),
    .ZN(_04640_));
 OAI22_X1 _18385_ (.A1(_04602_),
    .A2(_03147_),
    .B1(_03151_),
    .B2(_04606_),
    .ZN(_04641_));
 NOR2_X1 _18386_ (.A1(_04640_),
    .A2(_04641_),
    .ZN(_04642_));
 NAND2_X1 _18387_ (.A1(_04611_),
    .A2(_03168_),
    .ZN(_04643_));
 AOI21_X2 _18388_ (.A(_04601_),
    .B1(_04642_),
    .B2(_04643_),
    .ZN(net500));
 OAI22_X1 _18389_ (.A1(_04603_),
    .A2(_03173_),
    .B1(_03178_),
    .B2(_04617_),
    .ZN(_04644_));
 OAI22_X1 _18390_ (.A1(_04619_),
    .A2(_03183_),
    .B1(_03188_),
    .B2(_04595_),
    .ZN(_04645_));
 NOR2_X1 _18391_ (.A1(_04598_),
    .A2(_03209_),
    .ZN(_04646_));
 NOR3_X1 _18392_ (.A1(_04644_),
    .A2(_04645_),
    .A3(_04646_),
    .ZN(_04647_));
 NOR2_X1 _18393_ (.A1(_04586_),
    .A2(_04647_),
    .ZN(net501));
 BUF_X4 _18394_ (.A(_04594_),
    .Z(_04648_));
 BUF_X4 _18395_ (.A(_04590_),
    .Z(_04649_));
 OAI22_X1 _18396_ (.A1(_04648_),
    .A2(_03216_),
    .B1(_03220_),
    .B2(_04649_),
    .ZN(_04650_));
 OAI22_X1 _18397_ (.A1(_04635_),
    .A2(_03228_),
    .B1(_03234_),
    .B2(_06859_),
    .ZN(_04651_));
 NOR2_X1 _18398_ (.A1(_04598_),
    .A2(_03253_),
    .ZN(_04652_));
 NOR3_X1 _18399_ (.A1(_04650_),
    .A2(_04651_),
    .A3(_04652_),
    .ZN(_04653_));
 NOR2_X2 _18400_ (.A1(_04586_),
    .A2(_04653_),
    .ZN(net502));
 OAI22_X1 _18401_ (.A1(_04603_),
    .A2(_03259_),
    .B1(_03269_),
    .B2(_04649_),
    .ZN(_04654_));
 OAI22_X1 _18402_ (.A1(_06860_),
    .A2(_03264_),
    .B1(_03273_),
    .B2(_04595_),
    .ZN(_04655_));
 NOR2_X1 _18403_ (.A1(_04598_),
    .A2(_03294_),
    .ZN(_04656_));
 NOR3_X1 _18404_ (.A1(_04654_),
    .A2(_04655_),
    .A3(_04656_),
    .ZN(_04657_));
 NOR2_X1 _18405_ (.A1(_04586_),
    .A2(_04657_),
    .ZN(net503));
 OAI22_X1 _18406_ (.A1(_04602_),
    .A2(_03301_),
    .B1(_03305_),
    .B2(_04619_),
    .ZN(_04658_));
 OAI22_X1 _18407_ (.A1(_04589_),
    .A2(_03310_),
    .B1(_03314_),
    .B2(_04606_),
    .ZN(_04659_));
 NOR2_X1 _18408_ (.A1(_04658_),
    .A2(_04659_),
    .ZN(_04660_));
 NAND2_X1 _18409_ (.A1(_04611_),
    .A2(_03331_),
    .ZN(_04661_));
 AOI21_X2 _18410_ (.A(_04601_),
    .B1(_04660_),
    .B2(_04661_),
    .ZN(net504));
 OAI22_X1 _18411_ (.A1(_04603_),
    .A2(_03336_),
    .B1(_03341_),
    .B2(_04617_),
    .ZN(_04662_));
 OAI22_X1 _18412_ (.A1(_04592_),
    .A2(_03346_),
    .B1(_03350_),
    .B2(_04595_),
    .ZN(_04663_));
 NOR2_X1 _18413_ (.A1(_04598_),
    .A2(_03369_),
    .ZN(_04664_));
 NOR3_X1 _18414_ (.A1(_04662_),
    .A2(_04663_),
    .A3(_04664_),
    .ZN(_04665_));
 NOR2_X1 _18415_ (.A1(_04586_),
    .A2(_04665_),
    .ZN(net505));
 INV_X1 _18416_ (.A(_04587_),
    .ZN(_04666_));
 BUF_X4 _18417_ (.A(_04666_),
    .Z(_04667_));
 AOI22_X1 _18418_ (.A1(_04667_),
    .A2(_05775_),
    .B1(_06080_),
    .B2(_06806_),
    .ZN(_04668_));
 BUF_X4 _18419_ (.A(_04594_),
    .Z(_04669_));
 OAI221_X1 _18420_ (.A(_04668_),
    .B1(_03374_),
    .B2(_04649_),
    .C1(_04669_),
    .C2(_02494_),
    .ZN(_04670_));
 CLKBUF_X3 _18421_ (.A(_04609_),
    .Z(_04671_));
 AOI21_X1 _18422_ (.A(_04670_),
    .B1(_07132_),
    .B2(_04671_),
    .ZN(_04672_));
 NOR2_X1 _18423_ (.A1(_04586_),
    .A2(_04672_),
    .ZN(net506));
 INV_X2 _18424_ (.A(_05328_),
    .ZN(_04673_));
 BUF_X4 _18425_ (.A(_04673_),
    .Z(_04674_));
 INV_X1 _18426_ (.A(_04590_),
    .ZN(_04675_));
 BUF_X4 _18427_ (.A(_04675_),
    .Z(_04676_));
 AOI22_X1 _18428_ (.A1(_04674_),
    .A2(_05849_),
    .B1(_05796_),
    .B2(_04676_),
    .ZN(_04677_));
 BUF_X4 _18429_ (.A(_04587_),
    .Z(_04678_));
 BUF_X4 _18430_ (.A(_06858_),
    .Z(_04679_));
 OAI221_X1 _18431_ (.A(_04677_),
    .B1(_03383_),
    .B2(_04678_),
    .C1(_04679_),
    .C2(_03382_),
    .ZN(_04680_));
 AOI21_X1 _18432_ (.A(_04680_),
    .B1(_07156_),
    .B2(_04671_),
    .ZN(_04681_));
 NOR2_X1 _18433_ (.A1(_04586_),
    .A2(_04681_),
    .ZN(net507));
 BUF_X4 _18434_ (.A(_04585_),
    .Z(_04682_));
 AOI22_X2 _18435_ (.A1(_04674_),
    .A2(_05839_),
    .B1(_05799_),
    .B2(_04676_),
    .ZN(_04683_));
 OAI221_X2 _18436_ (.A(_04683_),
    .B1(_03389_),
    .B2(_04678_),
    .C1(_04679_),
    .C2(_03388_),
    .ZN(_04684_));
 AOI21_X1 _18437_ (.A(_04684_),
    .B1(_05956_),
    .B2(_04671_),
    .ZN(_04685_));
 NOR2_X1 _18438_ (.A1(_04682_),
    .A2(_04685_),
    .ZN(net508));
 AOI22_X1 _18439_ (.A1(_04674_),
    .A2(_05829_),
    .B1(_05802_),
    .B2(_04676_),
    .ZN(_04686_));
 OAI221_X1 _18440_ (.A(_04686_),
    .B1(_03395_),
    .B2(_04678_),
    .C1(_04679_),
    .C2(_03393_),
    .ZN(_04687_));
 AOI21_X1 _18441_ (.A(_04687_),
    .B1(_05902_),
    .B2(_04671_),
    .ZN(_04688_));
 NOR2_X1 _18442_ (.A1(_04682_),
    .A2(_04688_),
    .ZN(net509));
 AOI22_X1 _18443_ (.A1(_04674_),
    .A2(_05832_),
    .B1(_05792_),
    .B2(_04675_),
    .ZN(_04689_));
 OAI221_X1 _18444_ (.A(_04689_),
    .B1(_03400_),
    .B2(_04588_),
    .C1(_04679_),
    .C2(_03399_),
    .ZN(_04690_));
 AOI21_X1 _18445_ (.A(_04690_),
    .B1(_03403_),
    .B2(_04671_),
    .ZN(_04691_));
 NOR2_X1 _18446_ (.A1(_04682_),
    .A2(_04691_),
    .ZN(net510));
 AOI22_X1 _18447_ (.A1(_04674_),
    .A2(_05836_),
    .B1(_05809_),
    .B2(_04675_),
    .ZN(_04692_));
 OAI221_X1 _18448_ (.A(_04692_),
    .B1(_07233_),
    .B2(_04588_),
    .C1(_04679_),
    .C2(_07196_),
    .ZN(_04693_));
 AOI21_X1 _18449_ (.A(_04693_),
    .B1(_05972_),
    .B2(_04671_),
    .ZN(_04694_));
 NOR2_X2 _18450_ (.A1(_04682_),
    .A2(_04694_),
    .ZN(net511));
 AOI22_X1 _18451_ (.A1(_04674_),
    .A2(_05843_),
    .B1(_05806_),
    .B2(_04675_),
    .ZN(_04695_));
 OAI221_X1 _18452_ (.A(_04695_),
    .B1(_07229_),
    .B2(_04588_),
    .C1(_04679_),
    .C2(_07192_),
    .ZN(_04696_));
 AOI21_X1 _18453_ (.A(_04696_),
    .B1(_06008_),
    .B2(_04671_),
    .ZN(_04697_));
 NOR2_X1 _18454_ (.A1(_04682_),
    .A2(_04697_),
    .ZN(net512));
 AOI22_X2 _18455_ (.A1(_04667_),
    .A2(_05778_),
    .B1(_06071_),
    .B2(_06806_),
    .ZN(_04698_));
 OAI221_X2 _18456_ (.A(_04698_),
    .B1(_03412_),
    .B2(_04649_),
    .C1(_04669_),
    .C2(_07105_),
    .ZN(_04699_));
 AOI21_X2 _18457_ (.A(_04699_),
    .B1(_05993_),
    .B2(_04671_),
    .ZN(_04700_));
 NOR2_X2 _18458_ (.A1(_04682_),
    .A2(_04700_),
    .ZN(net513));
 OAI22_X1 _18459_ (.A1(_04603_),
    .A2(_03418_),
    .B1(_03422_),
    .B2(_04649_),
    .ZN(_04701_));
 OAI22_X1 _18460_ (.A1(_06860_),
    .A2(_03428_),
    .B1(_03432_),
    .B2(_04595_),
    .ZN(_04702_));
 NOR2_X1 _18461_ (.A1(_04598_),
    .A2(_03450_),
    .ZN(_04703_));
 NOR3_X1 _18462_ (.A1(_04701_),
    .A2(_04702_),
    .A3(_04703_),
    .ZN(_04704_));
 NOR2_X1 _18463_ (.A1(_04682_),
    .A2(_04704_),
    .ZN(net514));
 AOI22_X1 _18464_ (.A1(_04674_),
    .A2(_06524_),
    .B1(_05492_),
    .B2(_04667_),
    .ZN(_04705_));
 OAI221_X1 _18465_ (.A(_04705_),
    .B1(_05274_),
    .B2(_04649_),
    .C1(_04679_),
    .C2(_06099_),
    .ZN(_04706_));
 AOI21_X1 _18466_ (.A(_04706_),
    .B1(_06179_),
    .B2(_04671_),
    .ZN(_04707_));
 NOR2_X1 _18467_ (.A1(_04682_),
    .A2(_04707_),
    .ZN(net515));
 BUF_X4 _18468_ (.A(_04585_),
    .Z(_04708_));
 OAI22_X2 _18469_ (.A1(_04594_),
    .A2(_05376_),
    .B1(_06789_),
    .B2(_04587_),
    .ZN(_04709_));
 AOI221_X2 _18470_ (.A(_04709_),
    .B1(_06514_),
    .B2(_04676_),
    .C1(_06807_),
    .C2(_06100_),
    .ZN(_04710_));
 NAND2_X1 _18471_ (.A1(_04611_),
    .A2(_06146_),
    .ZN(_04711_));
 AOI21_X2 _18472_ (.A(_04708_),
    .B1(_04710_),
    .B2(_04711_),
    .ZN(net516));
 AOI22_X1 _18473_ (.A1(_04674_),
    .A2(_05370_),
    .B1(_05500_),
    .B2(_04667_),
    .ZN(_04712_));
 OAI221_X1 _18474_ (.A(_04712_),
    .B1(_06513_),
    .B2(_04591_),
    .C1(_04679_),
    .C2(_06098_),
    .ZN(_04713_));
 AOI21_X1 _18475_ (.A(_04713_),
    .B1(_06163_),
    .B2(_04671_),
    .ZN(_04714_));
 NOR2_X1 _18476_ (.A1(_04682_),
    .A2(_04714_),
    .ZN(net517));
 OAI22_X1 _18477_ (.A1(_04603_),
    .A2(_03465_),
    .B1(_03471_),
    .B2(_04617_),
    .ZN(_04715_));
 OAI22_X1 _18478_ (.A1(_04592_),
    .A2(_03476_),
    .B1(_03480_),
    .B2(_04595_),
    .ZN(_04716_));
 NOR2_X1 _18479_ (.A1(_04598_),
    .A2(_03498_),
    .ZN(_04717_));
 NOR3_X1 _18480_ (.A1(_04715_),
    .A2(_04716_),
    .A3(_04717_),
    .ZN(_04718_));
 NOR2_X1 _18481_ (.A1(_04682_),
    .A2(_04718_),
    .ZN(net518));
 OAI22_X2 _18482_ (.A1(_04591_),
    .A2(_03502_),
    .B1(_05327_),
    .B2(_05328_),
    .ZN(_04719_));
 AOI221_X2 _18483_ (.A(_04719_),
    .B1(_10348_),
    .B2(_04667_),
    .C1(_06807_),
    .C2(_10225_),
    .ZN(_04720_));
 NAND2_X1 _18484_ (.A1(_04611_),
    .A2(_10417_),
    .ZN(_04721_));
 AOI21_X4 _18485_ (.A(_04708_),
    .B1(_04720_),
    .B2(_04721_),
    .ZN(net519));
 OAI22_X2 _18486_ (.A1(_04587_),
    .A2(_10351_),
    .B1(_10255_),
    .B2(_04590_),
    .ZN(_04722_));
 AOI221_X2 _18487_ (.A(_04722_),
    .B1(net694),
    .B2(_04674_),
    .C1(_06807_),
    .C2(_04450_),
    .ZN(_04723_));
 NAND2_X1 _18488_ (.A1(_04611_),
    .A2(_07676_),
    .ZN(_04724_));
 AOI21_X2 _18489_ (.A(_04708_),
    .B1(_04723_),
    .B2(_04724_),
    .ZN(net520));
 BUF_X4 _18490_ (.A(_04585_),
    .Z(_04725_));
 AOI22_X1 _18491_ (.A1(_06807_),
    .A2(_07434_),
    .B1(_03510_),
    .B2(_04667_),
    .ZN(_04726_));
 OAI221_X1 _18492_ (.A(_04726_),
    .B1(_10261_),
    .B2(_04591_),
    .C1(_04669_),
    .C2(_10315_),
    .ZN(_04727_));
 AOI21_X1 _18493_ (.A(_04727_),
    .B1(_07661_),
    .B2(_04610_),
    .ZN(_04728_));
 NOR2_X1 _18494_ (.A1(_04725_),
    .A2(_04728_),
    .ZN(net521));
 AOI22_X1 _18495_ (.A1(_06807_),
    .A2(_07267_),
    .B1(_07305_),
    .B2(_04666_),
    .ZN(_04729_));
 OAI221_X1 _18496_ (.A(_04729_),
    .B1(_10258_),
    .B2(_04591_),
    .C1(_04669_),
    .C2(_10312_),
    .ZN(_04730_));
 AOI21_X1 _18497_ (.A(_04730_),
    .B1(_07409_),
    .B2(_04610_),
    .ZN(_04731_));
 NOR2_X2 _18498_ (.A1(_04725_),
    .A2(_04731_),
    .ZN(net522));
 AOI22_X1 _18499_ (.A1(_04676_),
    .A2(_07282_),
    .B1(_07431_),
    .B2(_06806_),
    .ZN(_04732_));
 OAI221_X1 _18500_ (.A(_04732_),
    .B1(_10369_),
    .B2(_04588_),
    .C1(_04669_),
    .C2(net697),
    .ZN(_04733_));
 AOI21_X1 _18501_ (.A(_04733_),
    .B1(_07646_),
    .B2(_04610_),
    .ZN(_04734_));
 NOR2_X1 _18502_ (.A1(_04725_),
    .A2(_04734_),
    .ZN(net523));
 OAI22_X2 _18503_ (.A1(_04591_),
    .A2(_10270_),
    .B1(_10209_),
    .B2(_06858_),
    .ZN(_04735_));
 AOI221_X2 _18504_ (.A(_04735_),
    .B1(_03522_),
    .B2(_04667_),
    .C1(_04674_),
    .C2(net665),
    .ZN(_04736_));
 NAND2_X1 _18505_ (.A1(_04611_),
    .A2(_07631_),
    .ZN(_04737_));
 AOI21_X2 _18506_ (.A(_04708_),
    .B1(_04736_),
    .B2(_04737_),
    .ZN(net524));
 OAI22_X1 _18507_ (.A1(_04602_),
    .A2(_03530_),
    .B1(_03539_),
    .B2(_04635_),
    .ZN(_04738_));
 OAI22_X1 _18508_ (.A1(_04592_),
    .A2(_03534_),
    .B1(_03543_),
    .B2(_04594_),
    .ZN(_04739_));
 CLKBUF_X3 _18509_ (.A(_04597_),
    .Z(_04740_));
 NOR2_X1 _18510_ (.A1(_04740_),
    .A2(_03562_),
    .ZN(_04741_));
 NOR3_X1 _18511_ (.A1(_04738_),
    .A2(_04739_),
    .A3(_04741_),
    .ZN(_04742_));
 NOR2_X2 _18512_ (.A1(_04725_),
    .A2(_04742_),
    .ZN(net525));
 OAI22_X2 _18513_ (.A1(_06858_),
    .A2(_10206_),
    .B1(_10303_),
    .B2(_05328_),
    .ZN(_04743_));
 AOI221_X2 _18514_ (.A(_04743_),
    .B1(_03566_),
    .B2(_04667_),
    .C1(_04676_),
    .C2(_07473_),
    .ZN(_04744_));
 BUF_X4 _18515_ (.A(_04610_),
    .Z(_04745_));
 NAND2_X1 _18516_ (.A1(_04745_),
    .A2(_07616_),
    .ZN(_04746_));
 AOI21_X4 _18517_ (.A(_04708_),
    .B1(_04744_),
    .B2(_04746_),
    .ZN(net526));
 OAI22_X2 _18518_ (.A1(_04605_),
    .A2(net640),
    .B1(net713),
    .B2(_04635_),
    .ZN(_04747_));
 OAI22_X2 _18519_ (.A1(_04602_),
    .A2(net650),
    .B1(net632),
    .B2(_04606_),
    .ZN(_04748_));
 NOR2_X2 _18520_ (.A1(_04747_),
    .A2(_04748_),
    .ZN(_04749_));
 NAND2_X1 _18521_ (.A1(_04745_),
    .A2(_07394_),
    .ZN(_04750_));
 AOI21_X4 _18522_ (.A(_04708_),
    .B1(_04749_),
    .B2(_04750_),
    .ZN(net527));
 AOI22_X1 _18523_ (.A1(_04676_),
    .A2(_10249_),
    .B1(_10276_),
    .B2(_04673_),
    .ZN(_04751_));
 OAI221_X1 _18524_ (.A(_04751_),
    .B1(_03574_),
    .B2(_04588_),
    .C1(_04679_),
    .C2(net685),
    .ZN(_04752_));
 AOI21_X1 _18525_ (.A(_04752_),
    .B1(_10372_),
    .B2(_04610_),
    .ZN(_04753_));
 NOR2_X1 _18526_ (.A1(_04725_),
    .A2(_04753_),
    .ZN(net528));
 OAI22_X1 _18527_ (.A1(_04587_),
    .A2(_10342_),
    .B1(_10279_),
    .B2(_05328_),
    .ZN(_04754_));
 INV_X1 _18528_ (.A(_04754_),
    .ZN(_04755_));
 OAI221_X1 _18529_ (.A(_04755_),
    .B1(net771),
    .B2(_04591_),
    .C1(_04617_),
    .C2(net643),
    .ZN(_04756_));
 AOI21_X1 _18530_ (.A(_04756_),
    .B1(_07556_),
    .B2(_04610_),
    .ZN(_04757_));
 NOR2_X1 _18531_ (.A1(_04725_),
    .A2(_04757_),
    .ZN(net529));
 OAI22_X2 _18532_ (.A1(_04590_),
    .A2(_10243_),
    .B1(net723),
    .B2(_04587_),
    .ZN(_04758_));
 INV_X1 _18533_ (.A(net645),
    .ZN(_04759_));
 AOI221_X2 _18534_ (.A(_04758_),
    .B1(net690),
    .B2(_04673_),
    .C1(_06807_),
    .C2(_04759_),
    .ZN(_04760_));
 NAND2_X1 _18535_ (.A1(_04745_),
    .A2(_07571_),
    .ZN(_04761_));
 AOI21_X2 _18536_ (.A(_04708_),
    .B1(_04760_),
    .B2(_04761_),
    .ZN(net530));
 OAI22_X2 _18537_ (.A1(_04590_),
    .A2(_10240_),
    .B1(_10285_),
    .B2(_05328_),
    .ZN(_04762_));
 AOI221_X2 _18538_ (.A(_04762_),
    .B1(_07296_),
    .B2(_04667_),
    .C1(_06807_),
    .C2(_04210_),
    .ZN(_04763_));
 NAND2_X1 _18539_ (.A1(_04745_),
    .A2(_07342_),
    .ZN(_04764_));
 AOI21_X2 _18540_ (.A(_04708_),
    .B1(_04763_),
    .B2(_04764_),
    .ZN(net531));
 OAI22_X2 _18541_ (.A1(_06858_),
    .A2(net647),
    .B1(_10288_),
    .B2(_05328_),
    .ZN(_04765_));
 AOI221_X2 _18542_ (.A(_04765_),
    .B1(net651),
    .B2(_04667_),
    .C1(_04676_),
    .C2(_03590_),
    .ZN(_04766_));
 NAND2_X1 _18543_ (.A1(_04745_),
    .A2(_07376_),
    .ZN(_04767_));
 AOI21_X2 _18544_ (.A(_04708_),
    .B1(_04766_),
    .B2(_04767_),
    .ZN(net532));
 OAI22_X2 _18545_ (.A1(_04587_),
    .A2(net703),
    .B1(_10234_),
    .B2(_04590_),
    .ZN(_04768_));
 AOI221_X2 _18546_ (.A(_04768_),
    .B1(_07489_),
    .B2(_04673_),
    .C1(_06807_),
    .C2(_04220_),
    .ZN(_04769_));
 NAND2_X1 _18547_ (.A1(_04745_),
    .A2(_07361_),
    .ZN(_04770_));
 AOI21_X2 _18548_ (.A(_04708_),
    .B1(_04769_),
    .B2(_04770_),
    .ZN(net533));
 AOI22_X1 _18549_ (.A1(_06806_),
    .A2(net752),
    .B1(_03599_),
    .B2(_04666_),
    .ZN(_04771_));
 OAI221_X1 _18550_ (.A(_04771_),
    .B1(net750),
    .B2(_04591_),
    .C1(_04669_),
    .C2(_10294_),
    .ZN(_04772_));
 AOI21_X1 _18551_ (.A(_04772_),
    .B1(_07601_),
    .B2(_04610_),
    .ZN(_04773_));
 NOR2_X2 _18552_ (.A1(_04725_),
    .A2(_04773_),
    .ZN(net534));
 OAI22_X1 _18553_ (.A1(_04605_),
    .A2(net731),
    .B1(net670),
    .B2(_04635_),
    .ZN(_04774_));
 OAI22_X1 _18554_ (.A1(_04602_),
    .A2(_10191_),
    .B1(_10297_),
    .B2(_04669_),
    .ZN(_04775_));
 NOR2_X1 _18555_ (.A1(_04774_),
    .A2(_04775_),
    .ZN(_04776_));
 NAND2_X1 _18556_ (.A1(_04745_),
    .A2(_07586_),
    .ZN(_04777_));
 AOI21_X4 _18557_ (.A(_04585_),
    .B1(_04776_),
    .B2(_04777_),
    .ZN(net535));
 OAI22_X1 _18558_ (.A1(_04602_),
    .A2(_03610_),
    .B1(_03614_),
    .B2(_04619_),
    .ZN(_04778_));
 OAI22_X1 _18559_ (.A1(_04589_),
    .A2(_03619_),
    .B1(_03623_),
    .B2(_04669_),
    .ZN(_04779_));
 NOR2_X1 _18560_ (.A1(_04778_),
    .A2(_04779_),
    .ZN(_04780_));
 NAND2_X1 _18561_ (.A1(_04745_),
    .A2(_03640_),
    .ZN(_04781_));
 AOI21_X4 _18562_ (.A(_04585_),
    .B1(_04780_),
    .B2(_04781_),
    .ZN(net536));
 OAI22_X2 _18563_ (.A1(_04605_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(_04617_),
    .ZN(_04782_));
 OAI22_X2 _18564_ (.A1(_04648_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_04678_),
    .ZN(_04783_));
 NOR2_X1 _18565_ (.A1(_04740_),
    .A2(_03655_),
    .ZN(_04784_));
 NOR3_X2 _18566_ (.A1(_04782_),
    .A2(_04783_),
    .A3(_04784_),
    .ZN(_04785_));
 NOR2_X4 _18567_ (.A1(_04725_),
    .A2(_04785_),
    .ZN(net537));
 AOI22_X1 _18568_ (.A1(_04676_),
    .A2(_05189_),
    .B1(_05649_),
    .B2(_06806_),
    .ZN(_04786_));
 OAI221_X1 _18569_ (.A(_04786_),
    .B1(_03662_),
    .B2(_04588_),
    .C1(_04669_),
    .C2(_03660_),
    .ZN(_04787_));
 AOI21_X1 _18570_ (.A(_04787_),
    .B1(_06249_),
    .B2(_04610_),
    .ZN(_04788_));
 NOR2_X2 _18571_ (.A1(_04725_),
    .A2(_04788_),
    .ZN(net538));
 OAI22_X2 _18572_ (.A1(_04605_),
    .A2(_03666_),
    .B1(_03669_),
    .B2(_04617_),
    .ZN(_04789_));
 OAI22_X2 _18573_ (.A1(_04648_),
    .A2(_03672_),
    .B1(_03674_),
    .B2(_04678_),
    .ZN(_04790_));
 NOR2_X1 _18574_ (.A1(_04740_),
    .A2(_03677_),
    .ZN(_04791_));
 NOR3_X2 _18575_ (.A1(_04789_),
    .A2(_04790_),
    .A3(_04791_),
    .ZN(_04792_));
 NOR2_X4 _18576_ (.A1(_04725_),
    .A2(_04792_),
    .ZN(net539));
 BUF_X4 _18577_ (.A(_04585_),
    .Z(_04793_));
 OAI22_X2 _18578_ (.A1(_04619_),
    .A2(_03681_),
    .B1(_03683_),
    .B2(_04635_),
    .ZN(_04794_));
 OAI22_X2 _18579_ (.A1(_04648_),
    .A2(_03686_),
    .B1(_03689_),
    .B2(_06859_),
    .ZN(_04795_));
 NOR2_X1 _18580_ (.A1(_04740_),
    .A2(_03692_),
    .ZN(_04796_));
 NOR3_X2 _18581_ (.A1(_04794_),
    .A2(_04795_),
    .A3(_04796_),
    .ZN(_04797_));
 NOR2_X2 _18582_ (.A1(_04793_),
    .A2(_04797_),
    .ZN(net540));
 OAI22_X2 _18583_ (.A1(_04619_),
    .A2(_03696_),
    .B1(_03699_),
    .B2(_04617_),
    .ZN(_04798_));
 OAI22_X2 _18584_ (.A1(_04648_),
    .A2(_03702_),
    .B1(_03704_),
    .B2(_04678_),
    .ZN(_04799_));
 NOR2_X1 _18585_ (.A1(_04740_),
    .A2(_03707_),
    .ZN(_04800_));
 NOR3_X2 _18586_ (.A1(_04798_),
    .A2(_04799_),
    .A3(_04800_),
    .ZN(_04801_));
 NOR2_X2 _18587_ (.A1(_04793_),
    .A2(_04801_),
    .ZN(net541));
 OAI22_X1 _18588_ (.A1(_04619_),
    .A2(_03717_),
    .B1(_03720_),
    .B2(_04617_),
    .ZN(_04802_));
 OAI22_X1 _18589_ (.A1(_04606_),
    .A2(_03712_),
    .B1(_03714_),
    .B2(_04678_),
    .ZN(_04803_));
 NOR2_X1 _18590_ (.A1(_04740_),
    .A2(_03723_),
    .ZN(_04804_));
 NOR3_X1 _18591_ (.A1(_04802_),
    .A2(_04803_),
    .A3(_04804_),
    .ZN(_04805_));
 NOR2_X2 _18592_ (.A1(_04793_),
    .A2(_04805_),
    .ZN(net542));
 OAI22_X1 _18593_ (.A1(_04589_),
    .A2(_03727_),
    .B1(_03730_),
    .B2(_06860_),
    .ZN(_04806_));
 OAI22_X1 _18594_ (.A1(_04605_),
    .A2(_03733_),
    .B1(_03735_),
    .B2(_04669_),
    .ZN(_04807_));
 NOR2_X1 _18595_ (.A1(_04806_),
    .A2(_04807_),
    .ZN(_04808_));
 NAND2_X1 _18596_ (.A1(_04745_),
    .A2(_03738_),
    .ZN(_04809_));
 AOI21_X4 _18597_ (.A(_04585_),
    .B1(_04808_),
    .B2(_04809_),
    .ZN(net543));
 OAI22_X2 _18598_ (.A1(_04648_),
    .A2(_03741_),
    .B1(_03743_),
    .B2(_04635_),
    .ZN(_04810_));
 OAI22_X2 _18599_ (.A1(_04592_),
    .A2(_03746_),
    .B1(_03749_),
    .B2(_06859_),
    .ZN(_04811_));
 NOR2_X1 _18600_ (.A1(_04740_),
    .A2(_03752_),
    .ZN(_04812_));
 NOR3_X2 _18601_ (.A1(_04810_),
    .A2(_04811_),
    .A3(_04812_),
    .ZN(_04813_));
 NOR2_X2 _18602_ (.A1(_04793_),
    .A2(_04813_),
    .ZN(net544));
 OAI22_X1 _18603_ (.A1(_04619_),
    .A2(_03756_),
    .B1(_03759_),
    .B2(_04617_),
    .ZN(_04814_));
 OAI22_X1 _18604_ (.A1(_04606_),
    .A2(_03762_),
    .B1(_03764_),
    .B2(_04678_),
    .ZN(_04815_));
 NOR2_X1 _18605_ (.A1(_04740_),
    .A2(_03767_),
    .ZN(_04816_));
 NOR3_X1 _18606_ (.A1(_04814_),
    .A2(_04815_),
    .A3(_04816_),
    .ZN(_04817_));
 NOR2_X2 _18607_ (.A1(_04793_),
    .A2(_04817_),
    .ZN(net545));
 OAI22_X1 _18608_ (.A1(_04648_),
    .A2(_03771_),
    .B1(_03773_),
    .B2(_04635_),
    .ZN(_04818_));
 OAI22_X1 _18609_ (.A1(_04592_),
    .A2(_03776_),
    .B1(_03779_),
    .B2(_06859_),
    .ZN(_04819_));
 NOR2_X1 _18610_ (.A1(_04740_),
    .A2(_03782_),
    .ZN(_04820_));
 NOR3_X1 _18611_ (.A1(_04818_),
    .A2(_04819_),
    .A3(_04820_),
    .ZN(_04821_));
 NOR2_X2 _18612_ (.A1(_04793_),
    .A2(_04821_),
    .ZN(net546));
 OAI22_X2 _18613_ (.A1(_04603_),
    .A2(_03788_),
    .B1(_03798_),
    .B2(_04649_),
    .ZN(_04822_));
 OAI22_X2 _18614_ (.A1(_06860_),
    .A2(_03793_),
    .B1(_03802_),
    .B2(_04594_),
    .ZN(_04823_));
 NOR2_X1 _18615_ (.A1(_04740_),
    .A2(_03820_),
    .ZN(_04824_));
 NOR3_X2 _18616_ (.A1(_04822_),
    .A2(_04823_),
    .A3(_04824_),
    .ZN(_04825_));
 NOR2_X2 _18617_ (.A1(_04793_),
    .A2(_04825_),
    .ZN(net547));
 AOI22_X2 _18618_ (.A1(_04676_),
    .A2(_05194_),
    .B1(_05639_),
    .B2(_06806_),
    .ZN(_04826_));
 OAI221_X2 _18619_ (.A(_04826_),
    .B1(_04281_),
    .B2(_04588_),
    .C1(_04595_),
    .C2(_04282_),
    .ZN(_04827_));
 AOI21_X2 _18620_ (.A(_04827_),
    .B1(_03827_),
    .B2(_04610_),
    .ZN(_04828_));
 NOR2_X2 _18621_ (.A1(_04793_),
    .A2(_04828_),
    .ZN(net548));
 OAI22_X2 _18622_ (.A1(_04648_),
    .A2(_03836_),
    .B1(_03833_),
    .B2(_04678_),
    .ZN(_04829_));
 OAI22_X2 _18623_ (.A1(_04592_),
    .A2(_03831_),
    .B1(_03839_),
    .B2(_06859_),
    .ZN(_04830_));
 NOR2_X1 _18624_ (.A1(_04597_),
    .A2(_03849_),
    .ZN(_04831_));
 NOR3_X2 _18625_ (.A1(_04829_),
    .A2(_04830_),
    .A3(_04831_),
    .ZN(_04832_));
 NOR2_X2 _18626_ (.A1(_04793_),
    .A2(_04832_),
    .ZN(net549));
 OAI22_X2 _18627_ (.A1(_04605_),
    .A2(_03853_),
    .B1(_03855_),
    .B2(_04648_),
    .ZN(_04833_));
 OAI22_X2 _18628_ (.A1(_04589_),
    .A2(_03858_),
    .B1(_03861_),
    .B2(_04679_),
    .ZN(_04834_));
 NOR2_X2 _18629_ (.A1(_04833_),
    .A2(_04834_),
    .ZN(_04835_));
 NAND2_X1 _18630_ (.A1(_04745_),
    .A2(_03864_),
    .ZN(_04836_));
 AOI21_X4 _18631_ (.A(_04585_),
    .B1(_04835_),
    .B2(_04836_),
    .ZN(net550));
 OAI22_X1 _18632_ (.A1(_04619_),
    .A2(_03867_),
    .B1(_03869_),
    .B2(_04678_),
    .ZN(_04837_));
 OAI22_X1 _18633_ (.A1(_04606_),
    .A2(_03872_),
    .B1(_03875_),
    .B2(_06859_),
    .ZN(_04838_));
 NOR2_X1 _18634_ (.A1(_04597_),
    .A2(_06229_),
    .ZN(_04839_));
 NOR3_X1 _18635_ (.A1(_04837_),
    .A2(_04838_),
    .A3(_04839_),
    .ZN(_04840_));
 NOR2_X2 _18636_ (.A1(_04793_),
    .A2(_04840_),
    .ZN(net551));
 OAI22_X2 _18637_ (.A1(_04603_),
    .A2(_03882_),
    .B1(_03887_),
    .B2(_06859_),
    .ZN(_04841_));
 OAI22_X2 _18638_ (.A1(_04592_),
    .A2(_03892_),
    .B1(_03896_),
    .B2(_04594_),
    .ZN(_04842_));
 NOR2_X1 _18639_ (.A1(_04597_),
    .A2(_03914_),
    .ZN(_04843_));
 NOR3_X2 _18640_ (.A1(_04841_),
    .A2(_04842_),
    .A3(_04843_),
    .ZN(_04844_));
 NOR2_X2 _18641_ (.A1(_04601_),
    .A2(_04844_),
    .ZN(net552));
 OAI22_X2 _18642_ (.A1(_04603_),
    .A2(_03920_),
    .B1(_03930_),
    .B2(_04649_),
    .ZN(_04845_));
 OAI22_X2 _18643_ (.A1(_06860_),
    .A2(_03925_),
    .B1(_03934_),
    .B2(_04594_),
    .ZN(_04846_));
 NOR2_X1 _18644_ (.A1(_04597_),
    .A2(_03952_),
    .ZN(_04847_));
 NOR3_X2 _18645_ (.A1(_04845_),
    .A2(_04846_),
    .A3(_04847_),
    .ZN(_04848_));
 NOR2_X2 _18646_ (.A1(_04601_),
    .A2(_04848_),
    .ZN(net553));
 OAI22_X2 _18647_ (.A1(_04648_),
    .A2(_03958_),
    .B1(_03962_),
    .B2(_04649_),
    .ZN(_04849_));
 OAI22_X2 _18648_ (.A1(_04635_),
    .A2(_03967_),
    .B1(_03972_),
    .B2(_06859_),
    .ZN(_04850_));
 NOR2_X1 _18649_ (.A1(_04597_),
    .A2(_03990_),
    .ZN(_04851_));
 NOR3_X2 _18650_ (.A1(_04849_),
    .A2(_04850_),
    .A3(_04851_),
    .ZN(_04852_));
 NOR2_X2 _18651_ (.A1(_04601_),
    .A2(_04852_),
    .ZN(net554));
 OAI22_X2 _18652_ (.A1(_04602_),
    .A2(_03997_),
    .B1(_04001_),
    .B2(_04649_),
    .ZN(_04853_));
 OAI22_X2 _18653_ (.A1(_04635_),
    .A2(_04006_),
    .B1(_04010_),
    .B2(_04594_),
    .ZN(_04854_));
 NOR2_X1 _18654_ (.A1(_04597_),
    .A2(_04028_),
    .ZN(_04855_));
 NOR3_X2 _18655_ (.A1(_04853_),
    .A2(_04854_),
    .A3(_04855_),
    .ZN(_04856_));
 NOR2_X2 _18656_ (.A1(_04601_),
    .A2(_04856_),
    .ZN(net555));
 BUF_X8 _18657_ (.A(_05474_),
    .Z(_04857_));
 BUF_X4 _18658_ (.A(_04857_),
    .Z(_04858_));
 BUF_X4 _18659_ (.A(_00051_),
    .Z(_04859_));
 BUF_X4 _18660_ (.A(_04859_),
    .Z(_04860_));
 BUF_X4 _18661_ (.A(_00064_),
    .Z(_04861_));
 BUF_X4 _18662_ (.A(_04861_),
    .Z(_04862_));
 BUF_X4 _18663_ (.A(_04862_),
    .Z(_04863_));
 OAI22_X1 _18664_ (.A1(_04860_),
    .A2(_02768_),
    .B1(_02777_),
    .B2(_04863_),
    .ZN(_04864_));
 BUF_X4 _18665_ (.A(_06611_),
    .Z(_04865_));
 BUF_X2 _18666_ (.A(_00062_),
    .Z(_04866_));
 BUF_X4 _18667_ (.A(_04866_),
    .Z(_04867_));
 BUF_X4 _18668_ (.A(_04867_),
    .Z(_04868_));
 OAI22_X1 _18669_ (.A1(_04865_),
    .A2(_02790_),
    .B1(_02798_),
    .B2(_04868_),
    .ZN(_04869_));
 BUF_X4 _18670_ (.A(_00063_),
    .Z(_04870_));
 CLKBUF_X3 _18671_ (.A(_04870_),
    .Z(_04871_));
 NOR2_X1 _18672_ (.A1(_04871_),
    .A2(_02840_),
    .ZN(_04872_));
 NOR3_X1 _18673_ (.A1(_04864_),
    .A2(_04869_),
    .A3(_04872_),
    .ZN(_04873_));
 NOR2_X2 _18674_ (.A1(_04858_),
    .A2(_04873_),
    .ZN(net556));
 BUF_X4 _18675_ (.A(_04857_),
    .Z(_04874_));
 BUF_X4 _18676_ (.A(_04862_),
    .Z(_04875_));
 BUF_X4 _18677_ (.A(_04859_),
    .Z(_04876_));
 OAI22_X1 _18678_ (.A1(_04875_),
    .A2(_02850_),
    .B1(_02854_),
    .B2(_04876_),
    .ZN(_04877_));
 CLKBUF_X3 _18679_ (.A(_04867_),
    .Z(_04878_));
 OAI22_X1 _18680_ (.A1(_06699_),
    .A2(_02864_),
    .B1(_02868_),
    .B2(_04878_),
    .ZN(_04879_));
 NOR2_X1 _18681_ (.A1(_04877_),
    .A2(_04879_),
    .ZN(_04880_));
 INV_X1 _18682_ (.A(_04870_),
    .ZN(_04881_));
 CLKBUF_X3 _18683_ (.A(_04881_),
    .Z(_04882_));
 BUF_X4 _18684_ (.A(_04882_),
    .Z(_04883_));
 NAND2_X1 _18685_ (.A1(_04883_),
    .A2(_02896_),
    .ZN(_04884_));
 AOI21_X2 _18686_ (.A(_04874_),
    .B1(_04880_),
    .B2(_04884_),
    .ZN(net557));
 OAI22_X1 _18687_ (.A1(_04860_),
    .A2(_02901_),
    .B1(_02905_),
    .B2(_06612_),
    .ZN(_04885_));
 OAI22_X1 _18688_ (.A1(_04875_),
    .A2(_02912_),
    .B1(_02916_),
    .B2(_04878_),
    .ZN(_04886_));
 NOR2_X1 _18689_ (.A1(_04885_),
    .A2(_04886_),
    .ZN(_04887_));
 NAND2_X1 _18690_ (.A1(_04883_),
    .A2(_02934_),
    .ZN(_04888_));
 AOI21_X2 _18691_ (.A(_04874_),
    .B1(_04887_),
    .B2(_04888_),
    .ZN(net558));
 OAI22_X1 _18692_ (.A1(_04860_),
    .A2(_02940_),
    .B1(_02946_),
    .B2(_04863_),
    .ZN(_04889_));
 OAI22_X1 _18693_ (.A1(_04865_),
    .A2(_02952_),
    .B1(_02956_),
    .B2(_04868_),
    .ZN(_04890_));
 NOR2_X1 _18694_ (.A1(_04871_),
    .A2(_02974_),
    .ZN(_04891_));
 NOR3_X1 _18695_ (.A1(_04889_),
    .A2(_04890_),
    .A3(_04891_),
    .ZN(_04892_));
 NOR2_X2 _18696_ (.A1(_04858_),
    .A2(_04892_),
    .ZN(net559));
 OAI22_X1 _18697_ (.A1(_04875_),
    .A2(_02981_),
    .B1(_02985_),
    .B2(_04876_),
    .ZN(_04893_));
 OAI22_X1 _18698_ (.A1(_06699_),
    .A2(_02990_),
    .B1(_02996_),
    .B2(_04878_),
    .ZN(_04894_));
 NOR2_X1 _18699_ (.A1(_04893_),
    .A2(_04894_),
    .ZN(_04895_));
 NAND2_X1 _18700_ (.A1(_04883_),
    .A2(_03013_),
    .ZN(_04896_));
 AOI21_X2 _18701_ (.A(_04874_),
    .B1(_04895_),
    .B2(_04896_),
    .ZN(net560));
 OAI22_X1 _18702_ (.A1(_04860_),
    .A2(_03019_),
    .B1(_03024_),
    .B2(_04863_),
    .ZN(_04897_));
 OAI22_X1 _18703_ (.A1(_04865_),
    .A2(_03030_),
    .B1(_03034_),
    .B2(_04868_),
    .ZN(_04898_));
 NOR2_X1 _18704_ (.A1(_04871_),
    .A2(_03055_),
    .ZN(_04899_));
 NOR3_X1 _18705_ (.A1(_04897_),
    .A2(_04898_),
    .A3(_04899_),
    .ZN(_04900_));
 NOR2_X2 _18706_ (.A1(_04858_),
    .A2(_04900_),
    .ZN(net561));
 OAI22_X1 _18707_ (.A1(_04860_),
    .A2(_03061_),
    .B1(_03065_),
    .B2(_06611_),
    .ZN(_04901_));
 OAI22_X1 _18708_ (.A1(_04863_),
    .A2(_03073_),
    .B1(_03077_),
    .B2(_04868_),
    .ZN(_04902_));
 NOR2_X1 _18709_ (.A1(_04871_),
    .A2(_03095_),
    .ZN(_04903_));
 NOR3_X1 _18710_ (.A1(_04901_),
    .A2(_04902_),
    .A3(_04903_),
    .ZN(_04904_));
 NOR2_X2 _18711_ (.A1(_04858_),
    .A2(_04904_),
    .ZN(net562));
 BUF_X4 _18712_ (.A(_04859_),
    .Z(_04905_));
 OAI22_X1 _18713_ (.A1(_06699_),
    .A2(_03106_),
    .B1(_03111_),
    .B2(_04905_),
    .ZN(_04906_));
 OAI22_X1 _18714_ (.A1(_04875_),
    .A2(_03102_),
    .B1(_03115_),
    .B2(_04878_),
    .ZN(_04907_));
 NOR2_X1 _18715_ (.A1(_04906_),
    .A2(_04907_),
    .ZN(_04908_));
 NAND2_X1 _18716_ (.A1(_04883_),
    .A2(_03132_),
    .ZN(_04909_));
 AOI21_X2 _18717_ (.A(_04874_),
    .B1(_04908_),
    .B2(_04909_),
    .ZN(net563));
 OAI22_X1 _18718_ (.A1(_04860_),
    .A2(_03137_),
    .B1(_03141_),
    .B2(_06612_),
    .ZN(_04910_));
 OAI22_X1 _18719_ (.A1(_04875_),
    .A2(_03147_),
    .B1(_03151_),
    .B2(_04878_),
    .ZN(_04911_));
 NOR2_X1 _18720_ (.A1(_04910_),
    .A2(_04911_),
    .ZN(_04912_));
 NAND2_X1 _18721_ (.A1(_04883_),
    .A2(_03168_),
    .ZN(_04913_));
 AOI21_X2 _18722_ (.A(_04874_),
    .B1(_04912_),
    .B2(_04913_),
    .ZN(net564));
 OAI22_X1 _18723_ (.A1(_04876_),
    .A2(_03173_),
    .B1(_03178_),
    .B2(_04863_),
    .ZN(_04914_));
 OAI22_X1 _18724_ (.A1(_04865_),
    .A2(_03183_),
    .B1(_03188_),
    .B2(_04868_),
    .ZN(_04915_));
 NOR2_X1 _18725_ (.A1(_04871_),
    .A2(_03209_),
    .ZN(_04916_));
 NOR3_X1 _18726_ (.A1(_04914_),
    .A2(_04915_),
    .A3(_04916_),
    .ZN(_04917_));
 NOR2_X1 _18727_ (.A1(_04858_),
    .A2(_04917_),
    .ZN(net565));
 CLKBUF_X3 _18728_ (.A(_04867_),
    .Z(_04918_));
 OAI22_X1 _18729_ (.A1(_04918_),
    .A2(_03216_),
    .B1(_03220_),
    .B2(_06611_),
    .ZN(_04919_));
 BUF_X4 _18730_ (.A(_04861_),
    .Z(_04920_));
 OAI22_X1 _18731_ (.A1(_04905_),
    .A2(_03228_),
    .B1(_03234_),
    .B2(_04920_),
    .ZN(_04921_));
 NOR2_X1 _18732_ (.A1(_04871_),
    .A2(_03253_),
    .ZN(_04922_));
 NOR3_X1 _18733_ (.A1(_04919_),
    .A2(_04921_),
    .A3(_04922_),
    .ZN(_04923_));
 NOR2_X1 _18734_ (.A1(_04858_),
    .A2(_04923_),
    .ZN(net566));
 OAI22_X1 _18735_ (.A1(_04876_),
    .A2(_03259_),
    .B1(_03264_),
    .B2(_04863_),
    .ZN(_04924_));
 OAI22_X1 _18736_ (.A1(_04865_),
    .A2(_03269_),
    .B1(_03273_),
    .B2(_04868_),
    .ZN(_04925_));
 NOR2_X1 _18737_ (.A1(_04871_),
    .A2(_03294_),
    .ZN(_04926_));
 NOR3_X1 _18738_ (.A1(_04924_),
    .A2(_04925_),
    .A3(_04926_),
    .ZN(_04927_));
 NOR2_X1 _18739_ (.A1(_04858_),
    .A2(_04927_),
    .ZN(net567));
 OAI22_X1 _18740_ (.A1(_04875_),
    .A2(_03301_),
    .B1(_03305_),
    .B2(_06612_),
    .ZN(_04928_));
 OAI22_X1 _18741_ (.A1(_04860_),
    .A2(_03310_),
    .B1(_03314_),
    .B2(_04878_),
    .ZN(_04929_));
 NOR2_X1 _18742_ (.A1(_04928_),
    .A2(_04929_),
    .ZN(_04930_));
 NAND2_X1 _18743_ (.A1(_04883_),
    .A2(_03331_),
    .ZN(_04931_));
 AOI21_X2 _18744_ (.A(_04874_),
    .B1(_04930_),
    .B2(_04931_),
    .ZN(net568));
 OAI22_X1 _18745_ (.A1(_04876_),
    .A2(_03336_),
    .B1(_03341_),
    .B2(_04863_),
    .ZN(_04932_));
 OAI22_X1 _18746_ (.A1(_04865_),
    .A2(_03346_),
    .B1(_03350_),
    .B2(_04868_),
    .ZN(_04933_));
 NOR2_X1 _18747_ (.A1(_04871_),
    .A2(_03369_),
    .ZN(_04934_));
 NOR3_X1 _18748_ (.A1(_04932_),
    .A2(_04933_),
    .A3(_04934_),
    .ZN(_04935_));
 NOR2_X1 _18749_ (.A1(_04858_),
    .A2(_04935_),
    .ZN(net569));
 INV_X2 _18750_ (.A(_04861_),
    .ZN(_04936_));
 BUF_X4 _18751_ (.A(_04936_),
    .Z(_04937_));
 AOI22_X1 _18752_ (.A1(_05469_),
    .A2(_05775_),
    .B1(_06080_),
    .B2(_04937_),
    .ZN(_04938_));
 BUF_X4 _18753_ (.A(_04867_),
    .Z(_04939_));
 OAI221_X1 _18754_ (.A(_04938_),
    .B1(_02494_),
    .B2(_04939_),
    .C1(_06691_),
    .C2(_03374_),
    .ZN(_04940_));
 BUF_X2 _18755_ (.A(_04881_),
    .Z(_04941_));
 AOI21_X1 _18756_ (.A(_04940_),
    .B1(_07132_),
    .B2(_04941_),
    .ZN(_04942_));
 NOR2_X2 _18757_ (.A1(_04858_),
    .A2(_04942_),
    .ZN(net570));
 INV_X4 _18758_ (.A(_04866_),
    .ZN(_04943_));
 BUF_X4 _18759_ (.A(_04943_),
    .Z(_04944_));
 AOI22_X2 _18760_ (.A1(_04944_),
    .A2(_05849_),
    .B1(_05796_),
    .B2(_06609_),
    .ZN(_04945_));
 OAI221_X2 _18761_ (.A(_04945_),
    .B1(_03382_),
    .B2(_04920_),
    .C1(_04905_),
    .C2(_03383_),
    .ZN(_04946_));
 AOI21_X1 _18762_ (.A(_04946_),
    .B1(_07156_),
    .B2(_04941_),
    .ZN(_04947_));
 NOR2_X1 _18763_ (.A1(_04858_),
    .A2(_04947_),
    .ZN(net571));
 BUF_X2 _18764_ (.A(_04857_),
    .Z(_04948_));
 AOI22_X1 _18765_ (.A1(_04944_),
    .A2(_05839_),
    .B1(_05799_),
    .B2(_06609_),
    .ZN(_04949_));
 OAI221_X1 _18766_ (.A(_04949_),
    .B1(_03388_),
    .B2(_04920_),
    .C1(_04905_),
    .C2(_03389_),
    .ZN(_04950_));
 AOI21_X1 _18767_ (.A(_04950_),
    .B1(_05956_),
    .B2(_04941_),
    .ZN(_04951_));
 NOR2_X1 _18768_ (.A1(_04948_),
    .A2(_04951_),
    .ZN(net572));
 AOI22_X1 _18769_ (.A1(_04944_),
    .A2(_05829_),
    .B1(_05802_),
    .B2(_06609_),
    .ZN(_04952_));
 OAI221_X1 _18770_ (.A(_04952_),
    .B1(_03393_),
    .B2(_04920_),
    .C1(_04905_),
    .C2(_03395_),
    .ZN(_04953_));
 AOI21_X1 _18771_ (.A(_04953_),
    .B1(_05902_),
    .B2(_04941_),
    .ZN(_04954_));
 NOR2_X1 _18772_ (.A1(_04948_),
    .A2(_04954_),
    .ZN(net573));
 AOI22_X1 _18773_ (.A1(_04944_),
    .A2(_05832_),
    .B1(_05792_),
    .B2(_06609_),
    .ZN(_04955_));
 OAI221_X1 _18774_ (.A(_04955_),
    .B1(_03399_),
    .B2(_04862_),
    .C1(_04905_),
    .C2(_03400_),
    .ZN(_04956_));
 AOI21_X1 _18775_ (.A(_04956_),
    .B1(_03403_),
    .B2(_04941_),
    .ZN(_04957_));
 NOR2_X1 _18776_ (.A1(_04948_),
    .A2(_04957_),
    .ZN(net574));
 AOI22_X1 _18777_ (.A1(_04944_),
    .A2(_05836_),
    .B1(_05809_),
    .B2(_06609_),
    .ZN(_04958_));
 BUF_X4 _18778_ (.A(_04859_),
    .Z(_04959_));
 OAI221_X1 _18779_ (.A(_04958_),
    .B1(_07196_),
    .B2(_04862_),
    .C1(_04959_),
    .C2(_07233_),
    .ZN(_04960_));
 AOI21_X1 _18780_ (.A(_04960_),
    .B1(_05972_),
    .B2(_04941_),
    .ZN(_04961_));
 NOR2_X1 _18781_ (.A1(_04948_),
    .A2(_04961_),
    .ZN(net575));
 AOI22_X1 _18782_ (.A1(_04944_),
    .A2(_05843_),
    .B1(_05806_),
    .B2(_06609_),
    .ZN(_04962_));
 OAI221_X1 _18783_ (.A(_04962_),
    .B1(_07192_),
    .B2(_04862_),
    .C1(_04959_),
    .C2(_07229_),
    .ZN(_04963_));
 AOI21_X1 _18784_ (.A(_04963_),
    .B1(_06008_),
    .B2(_04941_),
    .ZN(_04964_));
 NOR2_X1 _18785_ (.A1(_04948_),
    .A2(_04964_),
    .ZN(net576));
 AOI22_X1 _18786_ (.A1(_05469_),
    .A2(_05778_),
    .B1(_06071_),
    .B2(_04937_),
    .ZN(_04965_));
 OAI221_X1 _18787_ (.A(_04965_),
    .B1(_07105_),
    .B2(_04939_),
    .C1(_06691_),
    .C2(_03412_),
    .ZN(_04966_));
 AOI21_X1 _18788_ (.A(_04966_),
    .B1(_05993_),
    .B2(_04941_),
    .ZN(_04967_));
 NOR2_X1 _18789_ (.A1(_04948_),
    .A2(_04967_),
    .ZN(net577));
 BUF_X4 _18790_ (.A(_04861_),
    .Z(_04968_));
 OAI22_X2 _18791_ (.A1(_04876_),
    .A2(_03418_),
    .B1(_03428_),
    .B2(_04968_),
    .ZN(_04969_));
 OAI22_X2 _18792_ (.A1(_04865_),
    .A2(_03422_),
    .B1(_03432_),
    .B2(_04939_),
    .ZN(_04970_));
 NOR2_X1 _18793_ (.A1(_04871_),
    .A2(_03450_),
    .ZN(_04971_));
 NOR3_X2 _18794_ (.A1(_04971_),
    .A2(_04970_),
    .A3(_04969_),
    .ZN(_04972_));
 NOR2_X1 _18795_ (.A1(_04948_),
    .A2(_04972_),
    .ZN(net578));
 AOI22_X2 _18796_ (.A1(_04943_),
    .A2(_06524_),
    .B1(_05492_),
    .B2(_05469_),
    .ZN(_04973_));
 OAI221_X2 _18797_ (.A(_04973_),
    .B1(_06099_),
    .B2(_04862_),
    .C1(_06691_),
    .C2(_05274_),
    .ZN(_04974_));
 AOI21_X1 _18798_ (.A(_04974_),
    .B1(_06179_),
    .B2(_04941_),
    .ZN(_04975_));
 NOR2_X1 _18799_ (.A1(_04948_),
    .A2(_04975_),
    .ZN(net579));
 AOI22_X1 _18800_ (.A1(_07015_),
    .A2(_06514_),
    .B1(_06100_),
    .B2(_04937_),
    .ZN(_04976_));
 OAI221_X1 _18801_ (.A(_04976_),
    .B1(_05376_),
    .B2(_04939_),
    .C1(_04959_),
    .C2(_06789_),
    .ZN(_04977_));
 AOI21_X1 _18802_ (.A(_04977_),
    .B1(_06146_),
    .B2(_04941_),
    .ZN(_04978_));
 NOR2_X1 _18803_ (.A1(_04948_),
    .A2(_04978_),
    .ZN(net580));
 AOI22_X2 _18804_ (.A1(_04943_),
    .A2(_05370_),
    .B1(_05500_),
    .B2(_05469_),
    .ZN(_04979_));
 OAI221_X2 _18805_ (.A(_04979_),
    .B1(_06098_),
    .B2(_04862_),
    .C1(_06611_),
    .C2(_06513_),
    .ZN(_04980_));
 AOI21_X1 _18806_ (.A(_04980_),
    .B1(_06163_),
    .B2(_04882_),
    .ZN(_04981_));
 NOR2_X1 _18807_ (.A1(_04948_),
    .A2(_04981_),
    .ZN(net581));
 BUF_X4 _18808_ (.A(_04857_),
    .Z(_04982_));
 OAI22_X1 _18809_ (.A1(_04876_),
    .A2(_03465_),
    .B1(_03471_),
    .B2(_04968_),
    .ZN(_04983_));
 OAI22_X1 _18810_ (.A1(_04865_),
    .A2(_03476_),
    .B1(_03480_),
    .B2(_04939_),
    .ZN(_04984_));
 NOR2_X1 _18811_ (.A1(_04871_),
    .A2(_03498_),
    .ZN(_04985_));
 NOR3_X1 _18812_ (.A1(_04983_),
    .A2(_04984_),
    .A3(_04985_),
    .ZN(_04986_));
 NOR2_X1 _18813_ (.A1(_04982_),
    .A2(_04986_),
    .ZN(net582));
 AOI22_X1 _18814_ (.A1(_04937_),
    .A2(_10225_),
    .B1(_10348_),
    .B2(_05469_),
    .ZN(_04987_));
 OAI221_X1 _18815_ (.A(_04987_),
    .B1(_05327_),
    .B2(_04867_),
    .C1(_06611_),
    .C2(_03502_),
    .ZN(_04988_));
 AOI21_X1 _18816_ (.A(_04988_),
    .B1(_10417_),
    .B2(_04882_),
    .ZN(_04989_));
 NOR2_X2 _18817_ (.A1(_04982_),
    .A2(_04989_),
    .ZN(net583));
 BUF_X4 _18818_ (.A(_04857_),
    .Z(_04990_));
 OAI22_X2 _18819_ (.A1(_04859_),
    .A2(_10351_),
    .B1(_10255_),
    .B2(_06610_),
    .ZN(_04991_));
 AOI221_X2 _18820_ (.A(_04991_),
    .B1(_04450_),
    .B2(_04937_),
    .C1(_04944_),
    .C2(net694),
    .ZN(_04992_));
 NAND2_X1 _18821_ (.A1(_04883_),
    .A2(_07676_),
    .ZN(_04993_));
 AOI21_X2 _18822_ (.A(_04990_),
    .B1(_04992_),
    .B2(_04993_),
    .ZN(net584));
 OAI22_X2 _18823_ (.A1(_06610_),
    .A2(_10261_),
    .B1(_10315_),
    .B2(_04867_),
    .ZN(_04994_));
 AOI221_X2 _18824_ (.A(_04994_),
    .B1(_07434_),
    .B2(_04937_),
    .C1(_05469_),
    .C2(_03510_),
    .ZN(_04995_));
 NAND2_X1 _18825_ (.A1(_04883_),
    .A2(_07661_),
    .ZN(_04996_));
 AOI21_X2 _18826_ (.A(_04990_),
    .B1(_04995_),
    .B2(_04996_),
    .ZN(net585));
 OAI22_X2 _18827_ (.A1(_06610_),
    .A2(_10258_),
    .B1(_10354_),
    .B2(_04859_),
    .ZN(_04997_));
 AOI221_X2 _18828_ (.A(_04997_),
    .B1(_07267_),
    .B2(_04937_),
    .C1(_04944_),
    .C2(_04179_),
    .ZN(_04998_));
 NAND2_X1 _18829_ (.A1(_04883_),
    .A2(_07409_),
    .ZN(_04999_));
 AOI21_X2 _18830_ (.A(_04990_),
    .B1(_04998_),
    .B2(_04999_),
    .ZN(net586));
 AOI22_X2 _18831_ (.A1(_07015_),
    .A2(_07282_),
    .B1(net673),
    .B2(_04936_),
    .ZN(_05000_));
 OAI221_X2 _18832_ (.A(_05000_),
    .B1(net697),
    .B2(_04867_),
    .C1(_04959_),
    .C2(_10369_),
    .ZN(_05001_));
 AOI21_X1 _18833_ (.A(_05001_),
    .B1(_07646_),
    .B2(_04882_),
    .ZN(_05002_));
 NOR2_X2 _18834_ (.A1(_04982_),
    .A2(_05002_),
    .ZN(net587));
 AOI22_X2 _18835_ (.A1(_07015_),
    .A2(_07279_),
    .B1(net664),
    .B2(_04943_),
    .ZN(_05003_));
 OAI221_X2 _18836_ (.A(_05003_),
    .B1(_10209_),
    .B2(_04862_),
    .C1(_04959_),
    .C2(_10366_),
    .ZN(_05004_));
 AOI21_X1 _18837_ (.A(_05004_),
    .B1(_07631_),
    .B2(_04882_),
    .ZN(_05005_));
 NOR2_X1 _18838_ (.A1(_04982_),
    .A2(_05005_),
    .ZN(net588));
 OAI22_X1 _18839_ (.A1(_04875_),
    .A2(_03530_),
    .B1(_03534_),
    .B2(_06611_),
    .ZN(_05006_));
 OAI22_X1 _18840_ (.A1(_04905_),
    .A2(_03539_),
    .B1(_03543_),
    .B2(_04939_),
    .ZN(_05007_));
 CLKBUF_X3 _18841_ (.A(_04870_),
    .Z(_05008_));
 NOR2_X1 _18842_ (.A1(_05008_),
    .A2(_03562_),
    .ZN(_05009_));
 NOR3_X1 _18843_ (.A1(_05006_),
    .A2(_05007_),
    .A3(_05009_),
    .ZN(_05010_));
 NOR2_X2 _18844_ (.A1(_04982_),
    .A2(_05010_),
    .ZN(net589));
 AOI22_X1 _18845_ (.A1(_07015_),
    .A2(_07473_),
    .B1(_07506_),
    .B2(_04943_),
    .ZN(_05011_));
 OAI221_X1 _18846_ (.A(_05011_),
    .B1(_10206_),
    .B2(_04862_),
    .C1(_04959_),
    .C2(_10363_),
    .ZN(_05012_));
 AOI21_X1 _18847_ (.A(_05012_),
    .B1(_07616_),
    .B2(_04882_),
    .ZN(_05013_));
 NOR2_X2 _18848_ (.A1(_04982_),
    .A2(_05013_),
    .ZN(net590));
 OAI22_X1 _18849_ (.A1(_06699_),
    .A2(net640),
    .B1(net713),
    .B2(_04905_),
    .ZN(_05014_));
 OAI22_X2 _18850_ (.A1(_04875_),
    .A2(net650),
    .B1(net632),
    .B2(_04868_),
    .ZN(_05015_));
 NOR2_X1 _18851_ (.A1(_05014_),
    .A2(_05015_),
    .ZN(_05016_));
 NAND2_X1 _18852_ (.A1(_04883_),
    .A2(_07394_),
    .ZN(_05017_));
 AOI21_X2 _18853_ (.A(_04990_),
    .B1(_05016_),
    .B2(_05017_),
    .ZN(net591));
 AOI22_X1 _18854_ (.A1(_07015_),
    .A2(_10249_),
    .B1(_10276_),
    .B2(_04943_),
    .ZN(_05018_));
 OAI221_X1 _18855_ (.A(_05018_),
    .B1(net685),
    .B2(_04862_),
    .C1(_04959_),
    .C2(_03574_),
    .ZN(_05019_));
 AOI21_X1 _18856_ (.A(_05019_),
    .B1(_10372_),
    .B2(_04882_),
    .ZN(_05020_));
 NOR2_X2 _18857_ (.A1(_04982_),
    .A2(_05020_),
    .ZN(net592));
 OAI22_X2 _18858_ (.A1(_04861_),
    .A2(net642),
    .B1(_10246_),
    .B2(_06610_),
    .ZN(_05021_));
 AOI221_X2 _18859_ (.A(_05021_),
    .B1(_03578_),
    .B2(_04943_),
    .C1(_05469_),
    .C2(_03577_),
    .ZN(_05022_));
 CLKBUF_X3 _18860_ (.A(_04882_),
    .Z(_05023_));
 NAND2_X1 _18861_ (.A1(_05023_),
    .A2(_07556_),
    .ZN(_05024_));
 AOI21_X2 _18862_ (.A(_04990_),
    .B1(_05022_),
    .B2(_05024_),
    .ZN(net593));
 OAI22_X2 _18863_ (.A1(_04861_),
    .A2(net645),
    .B1(net723),
    .B2(_04859_),
    .ZN(_05025_));
 AOI221_X2 _18864_ (.A(_05025_),
    .B1(net689),
    .B2(_04943_),
    .C1(_07015_),
    .C2(_03583_),
    .ZN(_05026_));
 NAND2_X1 _18865_ (.A1(_05023_),
    .A2(_07571_),
    .ZN(_05027_));
 AOI21_X2 _18866_ (.A(_04990_),
    .B1(_05026_),
    .B2(_05027_),
    .ZN(net594));
 OAI22_X2 _18867_ (.A1(_06610_),
    .A2(_10240_),
    .B1(_10336_),
    .B2(_04859_),
    .ZN(_05028_));
 AOI221_X2 _18868_ (.A(_05028_),
    .B1(_04210_),
    .B2(_04937_),
    .C1(_04944_),
    .C2(_04211_),
    .ZN(_05029_));
 NAND2_X1 _18869_ (.A1(_05023_),
    .A2(_07342_),
    .ZN(_05030_));
 AOI21_X2 _18870_ (.A(_04990_),
    .B1(_05029_),
    .B2(_05030_),
    .ZN(net595));
 OAI22_X2 _18871_ (.A1(_04861_),
    .A2(net647),
    .B1(_10288_),
    .B2(_04867_),
    .ZN(_05031_));
 AOI221_X2 _18872_ (.A(_05031_),
    .B1(net651),
    .B2(_05469_),
    .C1(_07015_),
    .C2(_03590_),
    .ZN(_05032_));
 NAND2_X1 _18873_ (.A1(_05023_),
    .A2(_07376_),
    .ZN(_05033_));
 AOI21_X2 _18874_ (.A(_04990_),
    .B1(_05032_),
    .B2(_05033_),
    .ZN(net596));
 OAI22_X2 _18875_ (.A1(_04859_),
    .A2(net703),
    .B1(_10234_),
    .B2(_06610_),
    .ZN(_05034_));
 AOI221_X2 _18876_ (.A(_05034_),
    .B1(_04220_),
    .B2(_04937_),
    .C1(_04944_),
    .C2(_07489_),
    .ZN(_05035_));
 NAND2_X1 _18877_ (.A1(_05023_),
    .A2(_07361_),
    .ZN(_05036_));
 AOI21_X2 _18878_ (.A(_04990_),
    .B1(_05035_),
    .B2(_05036_),
    .ZN(net597));
 OAI22_X2 _18879_ (.A1(_06610_),
    .A2(net730),
    .B1(_10294_),
    .B2(_04866_),
    .ZN(_05037_));
 AOI221_X2 _18880_ (.A(_05037_),
    .B1(net753),
    .B2(_04937_),
    .C1(_05469_),
    .C2(_03599_),
    .ZN(_05038_));
 NAND2_X1 _18881_ (.A1(_05023_),
    .A2(_07601_),
    .ZN(_05039_));
 AOI21_X2 _18882_ (.A(_04990_),
    .B1(_05038_),
    .B2(_05039_),
    .ZN(net598));
 OAI22_X1 _18883_ (.A1(_06699_),
    .A2(net731),
    .B1(net670),
    .B2(_04905_),
    .ZN(_05040_));
 OAI22_X1 _18884_ (.A1(_04875_),
    .A2(_10191_),
    .B1(_10297_),
    .B2(_04868_),
    .ZN(_05041_));
 NOR2_X1 _18885_ (.A1(_05040_),
    .A2(_05041_),
    .ZN(_05042_));
 NAND2_X1 _18886_ (.A1(_05023_),
    .A2(_07586_),
    .ZN(_05043_));
 AOI21_X4 _18887_ (.A(_04857_),
    .B1(_05042_),
    .B2(_05043_),
    .ZN(net599));
 OAI22_X2 _18888_ (.A1(_04875_),
    .A2(_03610_),
    .B1(_03614_),
    .B2(_04865_),
    .ZN(_05044_));
 OAI22_X2 _18889_ (.A1(_04860_),
    .A2(_03619_),
    .B1(_03623_),
    .B2(_04868_),
    .ZN(_05045_));
 NOR2_X2 _18890_ (.A1(_05044_),
    .A2(_05045_),
    .ZN(_05046_));
 NAND2_X1 _18891_ (.A1(_05023_),
    .A2(_03640_),
    .ZN(_05047_));
 AOI21_X4 _18892_ (.A(_04857_),
    .B1(_05046_),
    .B2(_05047_),
    .ZN(net600));
 OAI22_X1 _18893_ (.A1(_06699_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(_04968_),
    .ZN(_05048_));
 CLKBUF_X3 _18894_ (.A(_04859_),
    .Z(_05049_));
 OAI22_X1 _18895_ (.A1(_04918_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_05049_),
    .ZN(_05050_));
 NOR2_X1 _18896_ (.A1(_05008_),
    .A2(_03655_),
    .ZN(_05051_));
 NOR3_X1 _18897_ (.A1(_05048_),
    .A2(_05050_),
    .A3(_05051_),
    .ZN(_05052_));
 NOR2_X2 _18898_ (.A1(_04982_),
    .A2(_05052_),
    .ZN(net601));
 AOI22_X2 _18899_ (.A1(_07015_),
    .A2(_05189_),
    .B1(_05649_),
    .B2(_04936_),
    .ZN(_05053_));
 OAI221_X2 _18900_ (.A(_05053_),
    .B1(_03660_),
    .B2(_04867_),
    .C1(_04959_),
    .C2(_03662_),
    .ZN(_05054_));
 AOI21_X1 _18901_ (.A(_05054_),
    .B1(_06249_),
    .B2(_04882_),
    .ZN(_05055_));
 NOR2_X2 _18902_ (.A1(_04982_),
    .A2(_05055_),
    .ZN(net602));
 OAI22_X1 _18903_ (.A1(_06699_),
    .A2(_03666_),
    .B1(_03669_),
    .B2(_04968_),
    .ZN(_05056_));
 OAI22_X1 _18904_ (.A1(_04918_),
    .A2(_03672_),
    .B1(_03674_),
    .B2(_05049_),
    .ZN(_05057_));
 NOR2_X1 _18905_ (.A1(_05008_),
    .A2(_03677_),
    .ZN(_05058_));
 NOR3_X1 _18906_ (.A1(_05056_),
    .A2(_05057_),
    .A3(_05058_),
    .ZN(_05059_));
 NOR2_X2 _18907_ (.A1(_04982_),
    .A2(_05059_),
    .ZN(net603));
 BUF_X4 _18908_ (.A(_04857_),
    .Z(_05060_));
 OAI22_X1 _18909_ (.A1(_06612_),
    .A2(_03681_),
    .B1(_03683_),
    .B2(_04959_),
    .ZN(_05061_));
 OAI22_X1 _18910_ (.A1(_04918_),
    .A2(_03686_),
    .B1(_03689_),
    .B2(_04920_),
    .ZN(_05062_));
 NOR2_X1 _18911_ (.A1(_05008_),
    .A2(_03692_),
    .ZN(_05063_));
 NOR3_X1 _18912_ (.A1(_05061_),
    .A2(_05062_),
    .A3(_05063_),
    .ZN(_05064_));
 NOR2_X2 _18913_ (.A1(_05060_),
    .A2(_05064_),
    .ZN(net604));
 OAI22_X1 _18914_ (.A1(_06612_),
    .A2(_03696_),
    .B1(_03699_),
    .B2(_04968_),
    .ZN(_05065_));
 OAI22_X1 _18915_ (.A1(_04878_),
    .A2(_03702_),
    .B1(_03704_),
    .B2(_05049_),
    .ZN(_05066_));
 NOR2_X1 _18916_ (.A1(_05008_),
    .A2(_03707_),
    .ZN(_05067_));
 NOR3_X1 _18917_ (.A1(_05065_),
    .A2(_05066_),
    .A3(_05067_),
    .ZN(_05068_));
 NOR2_X2 _18918_ (.A1(_05060_),
    .A2(_05068_),
    .ZN(net605));
 OAI22_X1 _18919_ (.A1(_06612_),
    .A2(_03717_),
    .B1(_03720_),
    .B2(_04968_),
    .ZN(_05069_));
 OAI22_X1 _18920_ (.A1(_04878_),
    .A2(_03712_),
    .B1(_03714_),
    .B2(_05049_),
    .ZN(_05070_));
 NOR2_X1 _18921_ (.A1(_05008_),
    .A2(_03723_),
    .ZN(_05071_));
 NOR3_X1 _18922_ (.A1(_05069_),
    .A2(_05070_),
    .A3(_05071_),
    .ZN(_05072_));
 NOR2_X2 _18923_ (.A1(_05060_),
    .A2(_05072_),
    .ZN(net606));
 OAI22_X1 _18924_ (.A1(_06699_),
    .A2(_03733_),
    .B1(_03735_),
    .B2(_04918_),
    .ZN(_05073_));
 OAI22_X1 _18925_ (.A1(_04860_),
    .A2(_03727_),
    .B1(_03730_),
    .B2(_04863_),
    .ZN(_05074_));
 NOR2_X1 _18926_ (.A1(_05073_),
    .A2(_05074_),
    .ZN(_05075_));
 NAND2_X1 _18927_ (.A1(_05023_),
    .A2(_03738_),
    .ZN(_05076_));
 AOI21_X4 _18928_ (.A(_04857_),
    .B1(_05075_),
    .B2(_05076_),
    .ZN(net607));
 OAI22_X1 _18929_ (.A1(_04918_),
    .A2(_03741_),
    .B1(_03743_),
    .B2(_05049_),
    .ZN(_05077_));
 OAI22_X1 _18930_ (.A1(_04865_),
    .A2(_03746_),
    .B1(_03749_),
    .B2(_04920_),
    .ZN(_05078_));
 NOR2_X1 _18931_ (.A1(_05008_),
    .A2(_03752_),
    .ZN(_05079_));
 NOR3_X1 _18932_ (.A1(_05077_),
    .A2(_05078_),
    .A3(_05079_),
    .ZN(_05080_));
 NOR2_X2 _18933_ (.A1(_05060_),
    .A2(_05080_),
    .ZN(net608));
 OAI22_X1 _18934_ (.A1(_06612_),
    .A2(_03756_),
    .B1(_03759_),
    .B2(_04968_),
    .ZN(_05081_));
 OAI22_X1 _18935_ (.A1(_04878_),
    .A2(_03762_),
    .B1(_03764_),
    .B2(_05049_),
    .ZN(_05082_));
 NOR2_X1 _18936_ (.A1(_05008_),
    .A2(_03767_),
    .ZN(_05083_));
 NOR3_X1 _18937_ (.A1(_05081_),
    .A2(_05082_),
    .A3(_05083_),
    .ZN(_05084_));
 NOR2_X2 _18938_ (.A1(_05060_),
    .A2(_05084_),
    .ZN(net609));
 OAI22_X1 _18939_ (.A1(_04918_),
    .A2(_03771_),
    .B1(_03773_),
    .B2(_05049_),
    .ZN(_05085_));
 OAI22_X1 _18940_ (.A1(_06691_),
    .A2(_03776_),
    .B1(_03779_),
    .B2(_04920_),
    .ZN(_05086_));
 NOR2_X1 _18941_ (.A1(_05008_),
    .A2(_03782_),
    .ZN(_05087_));
 NOR3_X1 _18942_ (.A1(_05085_),
    .A2(_05086_),
    .A3(_05087_),
    .ZN(_05088_));
 NOR2_X2 _18943_ (.A1(_05060_),
    .A2(_05088_),
    .ZN(net610));
 OAI22_X1 _18944_ (.A1(_04876_),
    .A2(_03788_),
    .B1(_03793_),
    .B2(_04968_),
    .ZN(_05089_));
 OAI22_X1 _18945_ (.A1(_06691_),
    .A2(_03798_),
    .B1(_03802_),
    .B2(_04939_),
    .ZN(_05090_));
 NOR2_X1 _18946_ (.A1(_05008_),
    .A2(_03820_),
    .ZN(_05091_));
 NOR3_X1 _18947_ (.A1(_05089_),
    .A2(_05090_),
    .A3(_05091_),
    .ZN(_05092_));
 NOR2_X2 _18948_ (.A1(_05060_),
    .A2(_05092_),
    .ZN(net611));
 AOI22_X2 _18949_ (.A1(_07015_),
    .A2(_05194_),
    .B1(_05639_),
    .B2(_04936_),
    .ZN(_05093_));
 OAI221_X2 _18950_ (.A(_05093_),
    .B1(_04282_),
    .B2(_04867_),
    .C1(_04959_),
    .C2(_04281_),
    .ZN(_05094_));
 AOI21_X1 _18951_ (.A(_05094_),
    .B1(_03827_),
    .B2(_04882_),
    .ZN(_05095_));
 NOR2_X2 _18952_ (.A1(_05060_),
    .A2(_05095_),
    .ZN(net612));
 OAI22_X1 _18953_ (.A1(_04918_),
    .A2(_03836_),
    .B1(_03833_),
    .B2(_05049_),
    .ZN(_05096_));
 OAI22_X1 _18954_ (.A1(_06691_),
    .A2(_03831_),
    .B1(_03839_),
    .B2(_04920_),
    .ZN(_05097_));
 NOR2_X1 _18955_ (.A1(_04870_),
    .A2(_03849_),
    .ZN(_05098_));
 NOR3_X1 _18956_ (.A1(_05096_),
    .A2(_05097_),
    .A3(_05098_),
    .ZN(_05099_));
 NOR2_X2 _18957_ (.A1(_05060_),
    .A2(_05099_),
    .ZN(net613));
 OAI22_X2 _18958_ (.A1(_06699_),
    .A2(_03853_),
    .B1(_03855_),
    .B2(_04918_),
    .ZN(_05100_));
 OAI22_X2 _18959_ (.A1(_04860_),
    .A2(_03858_),
    .B1(_03861_),
    .B2(_04863_),
    .ZN(_05101_));
 NOR2_X2 _18960_ (.A1(_05100_),
    .A2(_05101_),
    .ZN(_05102_));
 NAND2_X1 _18961_ (.A1(_05023_),
    .A2(_03864_),
    .ZN(_05103_));
 AOI21_X4 _18962_ (.A(_04857_),
    .B1(_05102_),
    .B2(_05103_),
    .ZN(net614));
 OAI22_X1 _18963_ (.A1(_06612_),
    .A2(_03867_),
    .B1(_03875_),
    .B2(_04968_),
    .ZN(_05104_));
 OAI22_X1 _18964_ (.A1(_04878_),
    .A2(_03872_),
    .B1(_03869_),
    .B2(_05049_),
    .ZN(_05105_));
 NOR2_X1 _18965_ (.A1(_04870_),
    .A2(_06229_),
    .ZN(_05106_));
 NOR3_X1 _18966_ (.A1(_05104_),
    .A2(_05105_),
    .A3(_05106_),
    .ZN(_05107_));
 NOR2_X2 _18967_ (.A1(_05060_),
    .A2(_05107_),
    .ZN(net615));
 OAI22_X1 _18968_ (.A1(_04876_),
    .A2(_03882_),
    .B1(_03887_),
    .B2(_04968_),
    .ZN(_05108_));
 OAI22_X1 _18969_ (.A1(_06691_),
    .A2(_03892_),
    .B1(_03896_),
    .B2(_04939_),
    .ZN(_05109_));
 NOR2_X1 _18970_ (.A1(_04870_),
    .A2(_03914_),
    .ZN(_05110_));
 NOR3_X1 _18971_ (.A1(_05108_),
    .A2(_05109_),
    .A3(_05110_),
    .ZN(_05111_));
 NOR2_X1 _18972_ (.A1(_04874_),
    .A2(_05111_),
    .ZN(net616));
 OAI22_X1 _18973_ (.A1(_04876_),
    .A2(_03920_),
    .B1(_03925_),
    .B2(_04920_),
    .ZN(_05112_));
 OAI22_X1 _18974_ (.A1(_06691_),
    .A2(_03930_),
    .B1(_03934_),
    .B2(_04939_),
    .ZN(_05113_));
 NOR2_X1 _18975_ (.A1(_04870_),
    .A2(_03952_),
    .ZN(_05114_));
 NOR3_X1 _18976_ (.A1(_05112_),
    .A2(_05113_),
    .A3(_05114_),
    .ZN(_05115_));
 NOR2_X1 _18977_ (.A1(_04874_),
    .A2(_05115_),
    .ZN(net617));
 OAI22_X1 _18978_ (.A1(_04918_),
    .A2(_03958_),
    .B1(_03967_),
    .B2(_05049_),
    .ZN(_05116_));
 OAI22_X1 _18979_ (.A1(_06691_),
    .A2(_03962_),
    .B1(_03972_),
    .B2(_04920_),
    .ZN(_05117_));
 NOR2_X1 _18980_ (.A1(_04870_),
    .A2(_03990_),
    .ZN(_05118_));
 NOR3_X1 _18981_ (.A1(_05116_),
    .A2(_05117_),
    .A3(_05118_),
    .ZN(_05119_));
 NOR2_X1 _18982_ (.A1(_04874_),
    .A2(_05119_),
    .ZN(net618));
 OAI22_X1 _18983_ (.A1(_04863_),
    .A2(_03997_),
    .B1(_04001_),
    .B2(_06611_),
    .ZN(_05120_));
 OAI22_X1 _18984_ (.A1(_04905_),
    .A2(_04006_),
    .B1(_04010_),
    .B2(_04939_),
    .ZN(_05121_));
 NOR2_X1 _18985_ (.A1(_04870_),
    .A2(_04028_),
    .ZN(_05122_));
 NOR3_X1 _18986_ (.A1(_05120_),
    .A2(_05121_),
    .A3(_05122_),
    .ZN(_05123_));
 NOR2_X1 _18987_ (.A1(_04874_),
    .A2(_05123_),
    .ZN(net619));
 FA_X1 _18988_ (.A(\dynamic_node_top.east_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.east_input.NIB.elements_in_array_f[1] ),
    .CI(_10162_),
    .CO(_10163_),
    .S(_10164_));
 FA_X1 _18989_ (.A(\dynamic_node_top.north_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.north_input.NIB.elements_in_array_f[1] ),
    .CI(_10165_),
    .CO(_10166_),
    .S(_10167_));
 FA_X1 _18990_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_next[0] ),
    .B(_10168_),
    .CI(_10169_),
    .CO(_10170_),
    .S(_10171_));
 FA_X1 _18991_ (.A(\dynamic_node_top.south_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.south_input.NIB.elements_in_array_f[1] ),
    .CI(_10172_),
    .CO(_10173_),
    .S(_10174_));
 FA_X1 _18992_ (.A(\dynamic_node_top.west_input.NIB.elements_in_array_f[0] ),
    .B(\dynamic_node_top.west_input.NIB.elements_in_array_f[1] ),
    .CI(_10175_),
    .CO(_10176_),
    .S(_10177_));
 HA_X1 _18993_ (.A(_10178_),
    .B(_10179_),
    .CO(_10180_),
    .S(_10181_));
 HA_X1 _18994_ (.A(_10182_),
    .B(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .CO(_10183_),
    .S(_10184_));
 HA_X1 _18995_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .B(_10185_),
    .CO(_10186_),
    .S(_10187_));
 HA_X1 _18996_ (.A(_10188_),
    .B(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .CO(_10189_),
    .S(_10190_));
 HA_X1 _18997_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .B(_10191_),
    .CO(_10192_),
    .S(_10193_));
 HA_X1 _18998_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .B(_10194_),
    .CO(_10195_),
    .S(_10196_));
 HA_X1 _18999_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .B(_10197_),
    .CO(_10198_),
    .S(_10199_));
 HA_X1 _19000_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .B(_10200_),
    .CO(_10201_),
    .S(_10202_));
 HA_X1 _19001_ (.A(_10203_),
    .B(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .CO(_10204_),
    .S(_10205_));
 HA_X1 _19002_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .B(_10206_),
    .CO(_10207_),
    .S(_10208_));
 HA_X1 _19003_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .B(_10209_),
    .CO(_10210_),
    .S(_10211_));
 HA_X1 _19004_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .B(_10212_),
    .CO(_10213_),
    .S(_10214_));
 HA_X1 _19005_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .B(_10215_),
    .CO(_10216_),
    .S(_10217_));
 HA_X1 _19006_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .B(_10218_),
    .CO(_10219_),
    .S(_10220_));
 HA_X1 _19007_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .B(_10221_),
    .CO(_10222_),
    .S(_10223_));
 HA_X1 _19008_ (.A(_10224_),
    .B(_10225_),
    .CO(_10226_),
    .S(_10227_));
 HA_X1 _19009_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .B(_10228_),
    .CO(_10229_),
    .S(_10230_));
 HA_X1 _19010_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .B(_10231_),
    .CO(_10232_),
    .S(_10233_));
 HA_X1 _19011_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .B(_10234_),
    .CO(_10235_),
    .S(_10236_));
 HA_X1 _19012_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .B(_10237_),
    .CO(_10238_),
    .S(_10239_));
 HA_X1 _19013_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .B(_10240_),
    .CO(_10241_),
    .S(_10242_));
 HA_X1 _19014_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .B(_10243_),
    .CO(_10244_),
    .S(_10245_));
 HA_X1 _19015_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .B(_10246_),
    .CO(_10247_),
    .S(_10248_));
 HA_X1 _19016_ (.A(_10178_),
    .B(_10249_),
    .CO(_10250_),
    .S(_10251_));
 HA_X1 _19017_ (.A(_10224_),
    .B(_10252_),
    .CO(_10253_),
    .S(_10254_));
 HA_X1 _19018_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .B(_10255_),
    .CO(_10256_),
    .S(_10257_));
 HA_X1 _19019_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .B(_10258_),
    .CO(_10259_),
    .S(_10260_));
 HA_X1 _19020_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .B(_10261_),
    .CO(_10262_),
    .S(_10263_));
 HA_X1 _19021_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .B(_10264_),
    .CO(_10265_),
    .S(_10266_));
 HA_X1 _19022_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .B(_10267_),
    .CO(_10268_),
    .S(_10269_));
 HA_X1 _19023_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .B(_10270_),
    .CO(_10271_),
    .S(_10272_));
 HA_X1 _19024_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .B(_10273_),
    .CO(_10274_),
    .S(_10275_));
 HA_X1 _19025_ (.A(_10178_),
    .B(_10276_),
    .CO(_10277_),
    .S(_10278_));
 HA_X1 _19026_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .B(_10279_),
    .CO(_10280_),
    .S(_10281_));
 HA_X1 _19027_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .B(_10282_),
    .CO(_10283_),
    .S(_10284_));
 HA_X1 _19028_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .B(_10285_),
    .CO(_10286_),
    .S(_10287_));
 HA_X1 _19029_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .B(_10288_),
    .CO(_10289_),
    .S(_10290_));
 HA_X1 _19030_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .B(_10291_),
    .CO(_10292_),
    .S(_10293_));
 HA_X1 _19031_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .B(_10294_),
    .CO(_10295_),
    .S(_10296_));
 HA_X1 _19032_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .B(_10297_),
    .CO(_10298_),
    .S(_10299_));
 HA_X1 _19033_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .B(_10300_),
    .CO(_10301_),
    .S(_10302_));
 HA_X1 _19034_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .B(_10303_),
    .CO(_10304_),
    .S(_10305_));
 HA_X1 _19035_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .B(_10306_),
    .CO(_10307_),
    .S(_10308_));
 HA_X1 _19036_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .B(_10309_),
    .CO(_10310_),
    .S(_10311_));
 HA_X1 _19037_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .B(_10312_),
    .CO(_10313_),
    .S(_10314_));
 HA_X1 _19038_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .B(_10315_),
    .CO(_10316_),
    .S(_10317_));
 HA_X1 _19039_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .B(_10318_),
    .CO(_10319_),
    .S(_10320_));
 HA_X1 _19040_ (.A(_10224_),
    .B(_10321_),
    .CO(_10322_),
    .S(_10323_));
 HA_X1 _19041_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .B(_10324_),
    .CO(_10325_),
    .S(_10326_));
 HA_X1 _19042_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .B(_10327_),
    .CO(_10328_),
    .S(_10329_));
 HA_X1 _19043_ (.A(_10330_),
    .B(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .CO(_10331_),
    .S(_10332_));
 HA_X1 _19044_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .B(_10333_),
    .CO(_10334_),
    .S(_10335_));
 HA_X1 _19045_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .B(_10336_),
    .CO(_10337_),
    .S(_10338_));
 HA_X1 _19046_ (.A(_10339_),
    .B(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .CO(_10340_),
    .S(_10341_));
 HA_X1 _19047_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .B(_10342_),
    .CO(_10343_),
    .S(_10344_));
 HA_X1 _19048_ (.A(_10178_),
    .B(_10345_),
    .CO(_10346_),
    .S(_10347_));
 HA_X1 _19049_ (.A(_10224_),
    .B(_10348_),
    .CO(_10349_),
    .S(_10350_));
 HA_X1 _19050_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .B(_10351_),
    .CO(_10352_),
    .S(_10353_));
 HA_X1 _19051_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .B(_10354_),
    .CO(_10355_),
    .S(_10356_));
 HA_X1 _19052_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .B(_10357_),
    .CO(_10358_),
    .S(_10359_));
 HA_X1 _19053_ (.A(_10360_),
    .B(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .CO(_10361_),
    .S(_10362_));
 HA_X1 _19054_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .B(_10363_),
    .CO(_10364_),
    .S(_10365_));
 HA_X1 _19055_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .B(_10366_),
    .CO(_10367_),
    .S(_10368_));
 HA_X1 _19056_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .B(_10369_),
    .CO(_10370_),
    .S(_10371_));
 HA_X1 _19057_ (.A(_10178_),
    .B(_10372_),
    .CO(_10373_),
    .S(_10374_));
 HA_X1 _19058_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .B(_10375_),
    .CO(_10376_),
    .S(_10377_));
 HA_X1 _19059_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .B(_10378_),
    .CO(_10379_),
    .S(_10380_));
 HA_X1 _19060_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .B(_10381_),
    .CO(_10382_),
    .S(_10383_));
 HA_X1 _19061_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .B(_10384_),
    .CO(_10385_),
    .S(_10386_));
 HA_X1 _19062_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .B(_10387_),
    .CO(_10388_),
    .S(_10389_));
 HA_X1 _19063_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .B(_10390_),
    .CO(_10391_),
    .S(_10392_));
 HA_X1 _19064_ (.A(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .B(_10393_),
    .CO(_10394_),
    .S(_10395_));
 HA_X1 _19065_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .B(_10396_),
    .CO(_10397_),
    .S(_10398_));
 HA_X1 _19066_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .B(_10399_),
    .CO(_10400_),
    .S(_10401_));
 HA_X1 _19067_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .B(_10402_),
    .CO(_10403_),
    .S(_10404_));
 HA_X1 _19068_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .B(_10405_),
    .CO(_10406_),
    .S(_10407_));
 HA_X1 _19069_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .B(_10408_),
    .CO(_10409_),
    .S(_10410_));
 HA_X1 _19070_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .B(_10411_),
    .CO(_10412_),
    .S(_10413_));
 HA_X1 _19071_ (.A(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .B(_10414_),
    .CO(_10415_),
    .S(_10416_));
 HA_X1 _19072_ (.A(_10224_),
    .B(_10417_),
    .CO(_10418_),
    .S(_10419_));
 HA_X1 _19073_ (.A(_10420_),
    .B(_10421_),
    .CO(_10422_),
    .S(_10423_));
 HA_X1 _19074_ (.A(_10424_),
    .B(\dynamic_node_top.east_output.space.valid_f ),
    .CO(_10425_),
    .S(_10426_));
 HA_X1 _19075_ (.A(\dynamic_node_top.east_output.space.yummy_f ),
    .B(_10427_),
    .CO(_10428_),
    .S(_10429_));
 HA_X1 _19076_ (.A(_10430_),
    .B(_10431_),
    .CO(_10432_),
    .S(_10433_));
 HA_X1 _19077_ (.A(_10430_),
    .B(_10431_),
    .CO(_10434_),
    .S(_10435_));
 HA_X1 _19078_ (.A(\dynamic_node_top.east_output.space.count_f[0] ),
    .B(\dynamic_node_top.east_output.space.count_f[1] ),
    .CO(_10436_),
    .S(_10437_));
 HA_X1 _19079_ (.A(_10438_),
    .B(_10439_),
    .CO(_10440_),
    .S(_10441_));
 HA_X1 _19080_ (.A(_10442_),
    .B(\dynamic_node_top.west_output.space.valid_f ),
    .CO(_10443_),
    .S(_10444_));
 HA_X1 _19081_ (.A(\dynamic_node_top.west_output.space.yummy_f ),
    .B(_10445_),
    .CO(_10446_),
    .S(_10447_));
 HA_X1 _19082_ (.A(_10448_),
    .B(_10449_),
    .CO(_10450_),
    .S(_10451_));
 HA_X1 _19083_ (.A(_10448_),
    .B(_10449_),
    .CO(_10452_),
    .S(_10453_));
 HA_X1 _19084_ (.A(\dynamic_node_top.west_output.space.count_f[0] ),
    .B(\dynamic_node_top.west_output.space.count_f[1] ),
    .CO(_10454_),
    .S(_10455_));
 HA_X1 _19085_ (.A(_10456_),
    .B(_10457_),
    .CO(_10458_),
    .S(_10459_));
 HA_X1 _19086_ (.A(_10456_),
    .B(net292),
    .CO(_10169_),
    .S(_10460_));
 HA_X1 _19087_ (.A(net620),
    .B(_10457_),
    .CO(_10461_),
    .S(_10462_));
 HA_X1 _19088_ (.A(_10463_),
    .B(_10464_),
    .CO(_10465_),
    .S(_10466_));
 HA_X1 _19089_ (.A(_10463_),
    .B(\dynamic_node_top.south_input.NIB.thanks_in ),
    .CO(_10467_),
    .S(_10468_));
 HA_X1 _19090_ (.A(net293),
    .B(_10464_),
    .CO(_10469_),
    .S(_10470_));
 HA_X1 _19091_ (.A(_10471_),
    .B(_10472_),
    .CO(_10473_),
    .S(_10474_));
 HA_X1 _19092_ (.A(_10471_),
    .B(\dynamic_node_top.north_input.NIB.thanks_in ),
    .CO(_10475_),
    .S(_10476_));
 HA_X1 _19093_ (.A(net291),
    .B(_10472_),
    .CO(_10477_),
    .S(_10478_));
 HA_X1 _19094_ (.A(_10479_),
    .B(_10480_),
    .CO(_10481_),
    .S(_10482_));
 HA_X1 _19095_ (.A(_10483_),
    .B(\dynamic_node_top.south_output.space.valid_f ),
    .CO(_10484_),
    .S(_10485_));
 HA_X1 _19096_ (.A(\dynamic_node_top.south_output.space.yummy_f ),
    .B(_10486_),
    .CO(_10487_),
    .S(_10488_));
 HA_X1 _19097_ (.A(_10489_),
    .B(_10490_),
    .CO(_10491_),
    .S(_10492_));
 HA_X1 _19098_ (.A(_10489_),
    .B(_10490_),
    .CO(_10493_),
    .S(_10494_));
 HA_X1 _19099_ (.A(\dynamic_node_top.south_output.space.count_f[0] ),
    .B(\dynamic_node_top.south_output.space.count_f[1] ),
    .CO(_10495_),
    .S(_10496_));
 HA_X1 _19100_ (.A(_10497_),
    .B(_10498_),
    .CO(_10499_),
    .S(_10500_));
 HA_X1 _19101_ (.A(_10497_),
    .B(\dynamic_node_top.west_input.NIB.thanks_in ),
    .CO(_10501_),
    .S(_10502_));
 HA_X1 _19102_ (.A(net294),
    .B(_10498_),
    .CO(_10503_),
    .S(_10504_));
 HA_X1 _19103_ (.A(_10505_),
    .B(_10506_),
    .CO(_10507_),
    .S(_10508_));
 HA_X1 _19104_ (.A(_10505_),
    .B(\dynamic_node_top.east_input.NIB.thanks_in ),
    .CO(_10509_),
    .S(_10510_));
 HA_X1 _19105_ (.A(net290),
    .B(_10506_),
    .CO(_10511_),
    .S(_10512_));
 HA_X1 _19106_ (.A(_10513_),
    .B(_10514_),
    .CO(_10515_),
    .S(_10516_));
 HA_X1 _19107_ (.A(_10517_),
    .B(\dynamic_node_top.proc_output.space.valid_f ),
    .CO(_10518_),
    .S(_10519_));
 HA_X1 _19108_ (.A(\dynamic_node_top.proc_output.space.yummy_f ),
    .B(_10520_),
    .CO(_10521_),
    .S(_10522_));
 HA_X1 _19109_ (.A(_10523_),
    .B(_10524_),
    .CO(_10525_),
    .S(_10526_));
 HA_X1 _19110_ (.A(_10523_),
    .B(_10524_),
    .CO(_10527_),
    .S(_10528_));
 HA_X1 _19111_ (.A(\dynamic_node_top.proc_output.space.count_f[0] ),
    .B(\dynamic_node_top.proc_output.space.count_f[1] ),
    .CO(_10529_),
    .S(_10530_));
 HA_X1 _19112_ (.A(_10531_),
    .B(_10532_),
    .CO(_10533_),
    .S(_10534_));
 HA_X1 _19113_ (.A(_10535_),
    .B(\dynamic_node_top.north_output.space.valid_f ),
    .CO(_10536_),
    .S(_10537_));
 HA_X1 _19114_ (.A(\dynamic_node_top.north_output.space.yummy_f ),
    .B(_10538_),
    .CO(_10539_),
    .S(_10540_));
 HA_X1 _19115_ (.A(_10541_),
    .B(_10542_),
    .CO(_10543_),
    .S(_10544_));
 HA_X1 _19116_ (.A(_10541_),
    .B(_10542_),
    .CO(_10545_),
    .S(_10546_));
 HA_X1 _19117_ (.A(\dynamic_node_top.north_output.space.count_f[0] ),
    .B(\dynamic_node_top.north_output.space.count_f[1] ),
    .CO(_10547_),
    .S(_10548_));
 HA_X1 _19118_ (.A(_10448_),
    .B(_10443_),
    .CO(_10549_),
    .S(_10550_));
 HA_X1 _19119_ (.A(_10448_),
    .B(_10446_),
    .CO(_10551_),
    .S(_10552_));
 HA_X1 _19120_ (.A(_10523_),
    .B(_10518_),
    .CO(_10553_),
    .S(_10554_));
 HA_X1 _19121_ (.A(_10523_),
    .B(_10521_),
    .CO(_10555_),
    .S(_10556_));
 HA_X1 _19122_ (.A(_10489_),
    .B(_10484_),
    .CO(_10557_),
    .S(_10558_));
 HA_X1 _19123_ (.A(_10489_),
    .B(_10487_),
    .CO(_10559_),
    .S(_10560_));
 HA_X1 _19124_ (.A(_10541_),
    .B(_10536_),
    .CO(_10561_),
    .S(_10562_));
 HA_X1 _19125_ (.A(_10541_),
    .B(_10539_),
    .CO(_10563_),
    .S(_10564_));
 HA_X1 _19126_ (.A(_10430_),
    .B(_10425_),
    .CO(_10565_),
    .S(_10566_));
 HA_X1 _19127_ (.A(_10430_),
    .B(_10428_),
    .CO(_10567_),
    .S(_10568_));
 HA_X1 _19128_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[1] ),
    .B(_10569_),
    .CO(_10570_),
    .S(_10571_));
 HA_X1 _19129_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[2] ),
    .B(_10569_),
    .CO(_10572_),
    .S(_10573_));
 HA_X1 _19130_ (.A(\dynamic_node_top.proc_input.NIB.elements_in_array_f[3] ),
    .B(_10569_),
    .CO(_10574_),
    .S(_10575_));
 HA_X1 _19131_ (.A(\dynamic_node_top.east_input.NIB.tail_ptr_next[0] ),
    .B(_10576_),
    .CO(_10577_),
    .S(\dynamic_node_top.east_input.NIB.tail_ptr_next[1] ));
 HA_X1 _19132_ (.A(\dynamic_node_top.east_input.NIB.tail_ptr_next[0] ),
    .B(\dynamic_node_top.east_input.NIB.tail_ptr_f[1] ),
    .CO(_10578_),
    .S(_10579_));
 HA_X1 _19133_ (.A(\dynamic_node_top.east_input.NIB.tail_ptr_f[0] ),
    .B(_10576_),
    .CO(_10580_),
    .S(_10581_));
 HA_X1 _19134_ (.A(\dynamic_node_top.east_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.east_input.NIB.tail_ptr_f[1] ),
    .CO(_10582_),
    .S(_10583_));
 HA_X1 _19135_ (.A(\dynamic_node_top.north_input.NIB.tail_ptr_next[0] ),
    .B(_10584_),
    .CO(_10585_),
    .S(\dynamic_node_top.north_input.NIB.tail_ptr_next[1] ));
 HA_X1 _19136_ (.A(\dynamic_node_top.north_input.NIB.tail_ptr_next[0] ),
    .B(\dynamic_node_top.north_input.NIB.tail_ptr_f[1] ),
    .CO(_10586_),
    .S(_10587_));
 HA_X1 _19137_ (.A(\dynamic_node_top.north_input.NIB.tail_ptr_f[0] ),
    .B(_10584_),
    .CO(_10588_),
    .S(_10589_));
 HA_X1 _19138_ (.A(\dynamic_node_top.north_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.north_input.NIB.tail_ptr_f[1] ),
    .CO(_10590_),
    .S(_10591_));
 HA_X1 _19139_ (.A(\dynamic_node_top.proc_input.NIB.head_ptr_f[0] ),
    .B(\dynamic_node_top.proc_input.NIB.head_ptr_f[1] ),
    .CO(_10592_),
    .S(\dynamic_node_top.proc_input.NIB.head_ptr_next[1] ));
 HA_X1 _19140_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_next[0] ),
    .B(_10593_),
    .CO(_10594_),
    .S(\dynamic_node_top.proc_input.NIB.tail_ptr_next[1] ));
 HA_X1 _19141_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_next[0] ),
    .B(\dynamic_node_top.proc_input.NIB.tail_ptr_f[1] ),
    .CO(_10595_),
    .S(_10596_));
 HA_X1 _19142_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_f[0] ),
    .B(_10593_),
    .CO(_10597_),
    .S(_10598_));
 HA_X1 _19143_ (.A(\dynamic_node_top.proc_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.proc_input.NIB.tail_ptr_f[1] ),
    .CO(_10599_),
    .S(_10600_));
 HA_X1 _19144_ (.A(\dynamic_node_top.south_input.NIB.tail_ptr_next[0] ),
    .B(_10601_),
    .CO(_10602_),
    .S(\dynamic_node_top.south_input.NIB.tail_ptr_next[1] ));
 HA_X1 _19145_ (.A(\dynamic_node_top.south_input.NIB.tail_ptr_next[0] ),
    .B(\dynamic_node_top.south_input.NIB.tail_ptr_f[1] ),
    .CO(_10603_),
    .S(_10604_));
 HA_X1 _19146_ (.A(\dynamic_node_top.south_input.NIB.tail_ptr_f[0] ),
    .B(_10601_),
    .CO(_10605_),
    .S(_10606_));
 HA_X1 _19147_ (.A(\dynamic_node_top.south_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.south_input.NIB.tail_ptr_f[1] ),
    .CO(_10607_),
    .S(_10608_));
 HA_X1 _19148_ (.A(\dynamic_node_top.west_input.NIB.tail_ptr_next[0] ),
    .B(_10609_),
    .CO(_10610_),
    .S(\dynamic_node_top.west_input.NIB.tail_ptr_next[1] ));
 HA_X1 _19149_ (.A(\dynamic_node_top.west_input.NIB.tail_ptr_next[0] ),
    .B(\dynamic_node_top.west_input.NIB.tail_ptr_f[1] ),
    .CO(_10611_),
    .S(_10612_));
 HA_X1 _19150_ (.A(\dynamic_node_top.west_input.NIB.tail_ptr_f[0] ),
    .B(_10609_),
    .CO(_10613_),
    .S(_10614_));
 HA_X1 _19151_ (.A(\dynamic_node_top.west_input.NIB.tail_ptr_f[0] ),
    .B(\dynamic_node_top.west_input.NIB.tail_ptr_f[1] ),
    .CO(_10615_),
    .S(_10616_));
 DFF_X1 _19152_ (.D(_00077_),
    .CK(clknet_leaf_175_clk),
    .Q(_00015_),
    .QN(_10149_));
 DFF_X1 _19153_ (.D(_00078_),
    .CK(clknet_leaf_193_clk),
    .Q(_00016_),
    .QN(_10148_));
 DFF_X1 _19154_ (.D(_00079_),
    .CK(clknet_leaf_287_clk),
    .Q(_00013_),
    .QN(_10147_));
 DFF_X2 _19155_ (.D(_00080_),
    .CK(clknet_leaf_293_clk),
    .Q(_00014_),
    .QN(_10146_));
 DFF_X1 _19156_ (.D(_00081_),
    .CK(clknet_leaf_291_clk),
    .Q(_00005_),
    .QN(_10145_));
 DFF_X1 _19157_ (.D(_00082_),
    .CK(clknet_leaf_291_clk),
    .Q(_00006_),
    .QN(_10144_));
 DFF_X1 _19158_ (.D(_00083_),
    .CK(clknet_leaf_128_clk),
    .Q(_00009_),
    .QN(_10143_));
 DFF_X1 _19159_ (.D(_00084_),
    .CK(clknet_leaf_125_clk),
    .Q(_00010_),
    .QN(_10142_));
 DFF_X1 _19160_ (.D(_00085_),
    .CK(clknet_leaf_128_clk),
    .Q(_00011_),
    .QN(_10141_));
 DFF_X1 _19161_ (.D(_00086_),
    .CK(clknet_leaf_128_clk),
    .Q(_00012_),
    .QN(_10140_));
 DFF_X1 _19162_ (.D(_00087_),
    .CK(clknet_leaf_144_clk),
    .Q(_00007_),
    .QN(_10139_));
 DFF_X1 _19163_ (.D(_00088_),
    .CK(clknet_leaf_198_clk),
    .Q(_00008_),
    .QN(_10150_));
 DFF_X1 \dynamic_node_top.REG_reset_fin.q$_DFF_P_  (.D(net289),
    .CK(clknet_leaf_108_clk),
    .Q(\dynamic_node_top.REG_reset_fin.q ),
    .QN(_00056_));
 DFF_X1 \dynamic_node_top.east_input.NIB.elements_in_array_f[0]$_SDFFE_PP0N_  (.D(_00089_),
    .CK(clknet_leaf_175_clk),
    .Q(\dynamic_node_top.east_input.NIB.elements_in_array_f[0] ),
    .QN(\dynamic_node_top.east_input.NIB.elements_in_array_next[0] ));
 DFF_X1 \dynamic_node_top.east_input.NIB.elements_in_array_f[1]$_SDFFE_PP0N_  (.D(_00090_),
    .CK(clknet_leaf_175_clk),
    .Q(\dynamic_node_top.east_input.NIB.elements_in_array_f[1] ),
    .QN(_10138_));
 DFF_X1 \dynamic_node_top.east_input.NIB.elements_in_array_f[2]$_SDFFE_PP0N_  (.D(_00091_),
    .CK(clknet_leaf_167_clk),
    .Q(\dynamic_node_top.east_input.NIB.elements_in_array_f[2] ),
    .QN(_10137_));
 DFF_X1 \dynamic_node_top.east_input.NIB.head_ptr_f[0]$_SDFFE_PP0N_  (.D(_00092_),
    .CK(clknet_leaf_291_clk),
    .Q(\dynamic_node_top.east_input.NIB.head_ptr_f[0] ),
    .QN(\dynamic_node_top.east_input.NIB.head_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.east_input.NIB.head_ptr_f[1]$_SDFFE_PP0N_  (.D(_00082_),
    .CK(clknet_leaf_291_clk),
    .Q(\dynamic_node_top.east_input.NIB.head_ptr_f[1] ),
    .QN(_10136_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][0]$_DFFE_PP_  (.D(_00093_),
    .CK(clknet_leaf_246_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][0] ),
    .QN(_10135_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][10]$_DFFE_PP_  (.D(_00094_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][10] ),
    .QN(_10134_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][11]$_DFFE_PP_  (.D(_00095_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][11] ),
    .QN(_10133_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][12]$_DFFE_PP_  (.D(_00096_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][12] ),
    .QN(_10132_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][13]$_DFFE_PP_  (.D(_00097_),
    .CK(clknet_leaf_237_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][13] ),
    .QN(_10131_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][14]$_DFFE_PP_  (.D(_00098_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][14] ),
    .QN(_10130_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][15]$_DFFE_PP_  (.D(_00099_),
    .CK(clknet_leaf_246_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][15] ),
    .QN(_10129_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][16]$_DFFE_PP_  (.D(_00100_),
    .CK(clknet_leaf_237_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][16] ),
    .QN(_10128_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][17]$_DFFE_PP_  (.D(_00101_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][17] ),
    .QN(_10127_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][18]$_DFFE_PP_  (.D(_00102_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][18] ),
    .QN(_10126_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][19]$_DFFE_PP_  (.D(_00103_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][19] ),
    .QN(_10125_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][1]$_DFFE_PP_  (.D(_00104_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][1] ),
    .QN(_10124_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][20]$_DFFE_PP_  (.D(_00105_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][20] ),
    .QN(_10123_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][21]$_DFFE_PP_  (.D(_00106_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][21] ),
    .QN(_10122_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][22]$_DFFE_PP_  (.D(_00107_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][22] ),
    .QN(_10121_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][23]$_DFFE_PP_  (.D(_00108_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][23] ),
    .QN(_10120_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][24]$_DFFE_PP_  (.D(_00109_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][24] ),
    .QN(_10119_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][25]$_DFFE_PP_  (.D(_00110_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][25] ),
    .QN(_10118_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][26]$_DFFE_PP_  (.D(_00111_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][26] ),
    .QN(_10117_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][27]$_DFFE_PP_  (.D(_00112_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][27] ),
    .QN(_10116_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][28]$_DFFE_PP_  (.D(_00113_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][28] ),
    .QN(_10115_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][29]$_DFFE_PP_  (.D(_00114_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][29] ),
    .QN(_10114_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][2]$_DFFE_PP_  (.D(_00115_),
    .CK(clknet_leaf_228_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][2] ),
    .QN(_10113_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][30]$_DFFE_PP_  (.D(_00116_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][30] ),
    .QN(_10112_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][31]$_DFFE_PP_  (.D(_00117_),
    .CK(clknet_leaf_221_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][31] ),
    .QN(_10111_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][32]$_DFFE_PP_  (.D(_00118_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][32] ),
    .QN(_10110_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][33]$_DFFE_PP_  (.D(_00119_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][33] ),
    .QN(_10109_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][34]$_DFFE_PP_  (.D(_00120_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][34] ),
    .QN(_10108_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][35]$_DFFE_PP_  (.D(_00121_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][35] ),
    .QN(_10107_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][36]$_DFFE_PP_  (.D(_00122_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][36] ),
    .QN(_10106_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][37]$_DFFE_PP_  (.D(_00123_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][37] ),
    .QN(_10105_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][38]$_DFFE_PP_  (.D(_00124_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][38] ),
    .QN(_10104_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][39]$_DFFE_PP_  (.D(_00125_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][39] ),
    .QN(_10103_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][3]$_DFFE_PP_  (.D(_00126_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][3] ),
    .QN(_10102_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][40]$_DFFE_PP_  (.D(_00127_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][40] ),
    .QN(_10101_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][41]$_DFFE_PP_  (.D(_00128_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][41] ),
    .QN(_10100_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][42]$_DFFE_PP_  (.D(_00129_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][42] ),
    .QN(_10099_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][43]$_DFFE_PP_  (.D(_00130_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][43] ),
    .QN(_10098_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][44]$_DFFE_PP_  (.D(_00131_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][44] ),
    .QN(_10097_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][45]$_DFFE_PP_  (.D(_00132_),
    .CK(clknet_leaf_210_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][45] ),
    .QN(_10096_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][46]$_DFFE_PP_  (.D(_00133_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][46] ),
    .QN(_10095_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][47]$_DFFE_PP_  (.D(_00134_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][47] ),
    .QN(_10094_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][48]$_DFFE_PP_  (.D(_00135_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][48] ),
    .QN(_10093_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][49]$_DFFE_PP_  (.D(_00136_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][49] ),
    .QN(_10092_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][4]$_DFFE_PP_  (.D(_00137_),
    .CK(clknet_leaf_235_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][4] ),
    .QN(_10091_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][50]$_DFFE_PP_  (.D(_00138_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][50] ),
    .QN(_10090_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][51]$_DFFE_PP_  (.D(_00139_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][51] ),
    .QN(_10089_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][52]$_DFFE_PP_  (.D(_00140_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][52] ),
    .QN(_10088_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][53]$_DFFE_PP_  (.D(_00141_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][53] ),
    .QN(_10087_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][54]$_DFFE_PP_  (.D(_00142_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][54] ),
    .QN(_10086_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][55]$_DFFE_PP_  (.D(_00143_),
    .CK(clknet_leaf_287_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][55] ),
    .QN(_10085_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][56]$_DFFE_PP_  (.D(_00144_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][56] ),
    .QN(_10084_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][57]$_DFFE_PP_  (.D(_00145_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][57] ),
    .QN(_10083_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][58]$_DFFE_PP_  (.D(_00146_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][58] ),
    .QN(_10082_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][59]$_DFFE_PP_  (.D(_00147_),
    .CK(clknet_leaf_286_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][59] ),
    .QN(_10081_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][5]$_DFFE_PP_  (.D(_00148_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][5] ),
    .QN(_10080_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][60]$_DFFE_PP_  (.D(_00149_),
    .CK(clknet_leaf_287_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][60] ),
    .QN(_10079_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][61]$_DFFE_PP_  (.D(_00150_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][61] ),
    .QN(_10078_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][62]$_DFFE_PP_  (.D(_00151_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][62] ),
    .QN(_10077_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][63]$_DFFE_PP_  (.D(_00152_),
    .CK(clknet_leaf_290_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][63] ),
    .QN(_10076_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][6]$_DFFE_PP_  (.D(_00153_),
    .CK(clknet_leaf_237_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][6] ),
    .QN(_10075_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][7]$_DFFE_PP_  (.D(_00154_),
    .CK(clknet_leaf_237_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][7] ),
    .QN(_10074_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][8]$_DFFE_PP_  (.D(_00155_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][8] ),
    .QN(_10073_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[0][9]$_DFFE_PP_  (.D(_00156_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[0][9] ),
    .QN(_10072_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][0]$_DFFE_PP_  (.D(_00157_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][0] ),
    .QN(_10071_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][10]$_DFFE_PP_  (.D(_00158_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][10] ),
    .QN(_10070_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][11]$_DFFE_PP_  (.D(_00159_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][11] ),
    .QN(_10069_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][12]$_DFFE_PP_  (.D(_00160_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][12] ),
    .QN(_10068_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][13]$_DFFE_PP_  (.D(_00161_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][13] ),
    .QN(_10067_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][14]$_DFFE_PP_  (.D(_00162_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][14] ),
    .QN(_10066_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][15]$_DFFE_PP_  (.D(_00163_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][15] ),
    .QN(_10065_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][16]$_DFFE_PP_  (.D(_00164_),
    .CK(clknet_leaf_237_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][16] ),
    .QN(_10064_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][17]$_DFFE_PP_  (.D(_00165_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][17] ),
    .QN(_10063_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][18]$_DFFE_PP_  (.D(_00166_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][18] ),
    .QN(_10062_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][19]$_DFFE_PP_  (.D(_00167_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][19] ),
    .QN(_10061_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][1]$_DFFE_PP_  (.D(_00168_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][1] ),
    .QN(_10060_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][20]$_DFFE_PP_  (.D(_00169_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][20] ),
    .QN(_10059_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][21]$_DFFE_PP_  (.D(_00170_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][21] ),
    .QN(_10058_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][22]$_DFFE_PP_  (.D(_00171_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][22] ),
    .QN(_10057_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][23]$_DFFE_PP_  (.D(_00172_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][23] ),
    .QN(_10056_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][24]$_DFFE_PP_  (.D(_00173_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][24] ),
    .QN(_10055_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][25]$_DFFE_PP_  (.D(_00174_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][25] ),
    .QN(_10054_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][26]$_DFFE_PP_  (.D(_00175_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][26] ),
    .QN(_10053_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][27]$_DFFE_PP_  (.D(_00176_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][27] ),
    .QN(_10052_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][28]$_DFFE_PP_  (.D(_00177_),
    .CK(clknet_leaf_229_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][28] ),
    .QN(_10051_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][29]$_DFFE_PP_  (.D(_00178_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][29] ),
    .QN(_10050_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][2]$_DFFE_PP_  (.D(_00179_),
    .CK(clknet_leaf_229_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][2] ),
    .QN(_10049_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][30]$_DFFE_PP_  (.D(_00180_),
    .CK(clknet_leaf_229_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][30] ),
    .QN(_10048_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][31]$_DFFE_PP_  (.D(_00181_),
    .CK(clknet_leaf_221_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][31] ),
    .QN(_10047_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][32]$_DFFE_PP_  (.D(_00182_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][32] ),
    .QN(_10046_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][33]$_DFFE_PP_  (.D(_00183_),
    .CK(clknet_leaf_228_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][33] ),
    .QN(_10045_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][34]$_DFFE_PP_  (.D(_00184_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][34] ),
    .QN(_10044_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][35]$_DFFE_PP_  (.D(_00185_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][35] ),
    .QN(_10043_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][36]$_DFFE_PP_  (.D(_00186_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][36] ),
    .QN(_10042_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][37]$_DFFE_PP_  (.D(_00187_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][37] ),
    .QN(_10041_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][38]$_DFFE_PP_  (.D(_00188_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][38] ),
    .QN(_10040_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][39]$_DFFE_PP_  (.D(_00189_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][39] ),
    .QN(_10039_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][3]$_DFFE_PP_  (.D(_00190_),
    .CK(clknet_leaf_229_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][3] ),
    .QN(_10038_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][40]$_DFFE_PP_  (.D(_00191_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][40] ),
    .QN(_10037_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][41]$_DFFE_PP_  (.D(_00192_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][41] ),
    .QN(_10036_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][42]$_DFFE_PP_  (.D(_00193_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][42] ),
    .QN(_10035_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][43]$_DFFE_PP_  (.D(_00194_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][43] ),
    .QN(_10034_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][44]$_DFFE_PP_  (.D(_00195_),
    .CK(clknet_leaf_210_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][44] ),
    .QN(_10033_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][45]$_DFFE_PP_  (.D(_00196_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][45] ),
    .QN(_10032_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][46]$_DFFE_PP_  (.D(_00197_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][46] ),
    .QN(_10031_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][47]$_DFFE_PP_  (.D(_00198_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][47] ),
    .QN(_10030_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][48]$_DFFE_PP_  (.D(_00199_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][48] ),
    .QN(_10029_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][49]$_DFFE_PP_  (.D(_00200_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][49] ),
    .QN(_10028_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][4]$_DFFE_PP_  (.D(_00201_),
    .CK(clknet_leaf_235_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][4] ),
    .QN(_10027_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][50]$_DFFE_PP_  (.D(_00202_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][50] ),
    .QN(_10026_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][51]$_DFFE_PP_  (.D(_00203_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][51] ),
    .QN(_10025_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][52]$_DFFE_PP_  (.D(_00204_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][52] ),
    .QN(_10024_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][53]$_DFFE_PP_  (.D(_00205_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][53] ),
    .QN(_10023_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][54]$_DFFE_PP_  (.D(_00206_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][54] ),
    .QN(_10022_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][55]$_DFFE_PP_  (.D(_00207_),
    .CK(clknet_leaf_290_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][55] ),
    .QN(_10021_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][56]$_DFFE_PP_  (.D(_00208_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][56] ),
    .QN(_10020_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][57]$_DFFE_PP_  (.D(_00209_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][57] ),
    .QN(_10019_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][58]$_DFFE_PP_  (.D(_00210_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][58] ),
    .QN(_10018_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][59]$_DFFE_PP_  (.D(_00211_),
    .CK(clknet_leaf_286_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][59] ),
    .QN(_10017_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][5]$_DFFE_PP_  (.D(_00212_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][5] ),
    .QN(_10016_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][60]$_DFFE_PP_  (.D(_00213_),
    .CK(clknet_leaf_287_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][60] ),
    .QN(_10015_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][61]$_DFFE_PP_  (.D(_00214_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][61] ),
    .QN(_10014_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][62]$_DFFE_PP_  (.D(_00215_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][62] ),
    .QN(_10013_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][63]$_DFFE_PP_  (.D(_00216_),
    .CK(clknet_leaf_290_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][63] ),
    .QN(_10012_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][6]$_DFFE_PP_  (.D(_00217_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][6] ),
    .QN(_10011_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][7]$_DFFE_PP_  (.D(_00218_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][7] ),
    .QN(_10010_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][8]$_DFFE_PP_  (.D(_00219_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][8] ),
    .QN(_10009_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[1][9]$_DFFE_PP_  (.D(_00220_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[1][9] ),
    .QN(_10008_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][0]$_DFFE_PP_  (.D(_00221_),
    .CK(clknet_leaf_246_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][0] ),
    .QN(_10007_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][10]$_DFFE_PP_  (.D(_00222_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][10] ),
    .QN(_10006_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][11]$_DFFE_PP_  (.D(_00223_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][11] ),
    .QN(_10005_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][12]$_DFFE_PP_  (.D(_00224_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][12] ),
    .QN(_10004_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][13]$_DFFE_PP_  (.D(_00225_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][13] ),
    .QN(_10003_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][14]$_DFFE_PP_  (.D(_00226_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][14] ),
    .QN(_10002_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][15]$_DFFE_PP_  (.D(_00227_),
    .CK(clknet_leaf_246_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][15] ),
    .QN(_10001_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][16]$_DFFE_PP_  (.D(_00228_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][16] ),
    .QN(_10000_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][17]$_DFFE_PP_  (.D(_00229_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][17] ),
    .QN(_09999_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][18]$_DFFE_PP_  (.D(_00230_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][18] ),
    .QN(_09998_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][19]$_DFFE_PP_  (.D(_00231_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][19] ),
    .QN(_09997_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][1]$_DFFE_PP_  (.D(_00232_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][1] ),
    .QN(_09996_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][20]$_DFFE_PP_  (.D(_00233_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][20] ),
    .QN(_09995_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][21]$_DFFE_PP_  (.D(_00234_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][21] ),
    .QN(_09994_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][22]$_DFFE_PP_  (.D(_00235_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][22] ),
    .QN(_09993_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][23]$_DFFE_PP_  (.D(_00236_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][23] ),
    .QN(_09992_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][24]$_DFFE_PP_  (.D(_00237_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][24] ),
    .QN(_09991_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][25]$_DFFE_PP_  (.D(_00238_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][25] ),
    .QN(_09990_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][26]$_DFFE_PP_  (.D(_00239_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][26] ),
    .QN(_09989_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][27]$_DFFE_PP_  (.D(_00240_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][27] ),
    .QN(_09988_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][28]$_DFFE_PP_  (.D(_00241_),
    .CK(clknet_leaf_229_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][28] ),
    .QN(_09987_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][29]$_DFFE_PP_  (.D(_00242_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][29] ),
    .QN(_09986_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][2]$_DFFE_PP_  (.D(_00243_),
    .CK(clknet_leaf_228_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][2] ),
    .QN(_09985_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][30]$_DFFE_PP_  (.D(_00244_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][30] ),
    .QN(_09984_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][31]$_DFFE_PP_  (.D(_00245_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][31] ),
    .QN(_09983_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][32]$_DFFE_PP_  (.D(_00246_),
    .CK(clknet_leaf_221_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][32] ),
    .QN(_09982_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][33]$_DFFE_PP_  (.D(_00247_),
    .CK(clknet_leaf_228_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][33] ),
    .QN(_09981_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][34]$_DFFE_PP_  (.D(_00248_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][34] ),
    .QN(_09980_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][35]$_DFFE_PP_  (.D(_00249_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][35] ),
    .QN(_09979_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][36]$_DFFE_PP_  (.D(_00250_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][36] ),
    .QN(_09978_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][37]$_DFFE_PP_  (.D(_00251_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][37] ),
    .QN(_09977_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][38]$_DFFE_PP_  (.D(_00252_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][38] ),
    .QN(_09976_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][39]$_DFFE_PP_  (.D(_00253_),
    .CK(clknet_leaf_230_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][39] ),
    .QN(_09975_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][3]$_DFFE_PP_  (.D(_00254_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][3] ),
    .QN(_09974_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][40]$_DFFE_PP_  (.D(_00255_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][40] ),
    .QN(_09973_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][41]$_DFFE_PP_  (.D(_00256_),
    .CK(clknet_leaf_235_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][41] ),
    .QN(_09972_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][42]$_DFFE_PP_  (.D(_00257_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][42] ),
    .QN(_09971_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][43]$_DFFE_PP_  (.D(_00258_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][43] ),
    .QN(_09970_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][44]$_DFFE_PP_  (.D(_00259_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][44] ),
    .QN(_09969_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][45]$_DFFE_PP_  (.D(_00260_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][45] ),
    .QN(_09968_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][46]$_DFFE_PP_  (.D(_00261_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][46] ),
    .QN(_09967_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][47]$_DFFE_PP_  (.D(_00262_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][47] ),
    .QN(_09966_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][48]$_DFFE_PP_  (.D(_00263_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][48] ),
    .QN(_09965_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][49]$_DFFE_PP_  (.D(_00264_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][49] ),
    .QN(_09964_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][4]$_DFFE_PP_  (.D(_00265_),
    .CK(clknet_leaf_235_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][4] ),
    .QN(_09963_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][50]$_DFFE_PP_  (.D(_00266_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][50] ),
    .QN(_09962_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][51]$_DFFE_PP_  (.D(_00267_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][51] ),
    .QN(_09961_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][52]$_DFFE_PP_  (.D(_00268_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][52] ),
    .QN(_09960_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][53]$_DFFE_PP_  (.D(_00269_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][53] ),
    .QN(_09959_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][54]$_DFFE_PP_  (.D(_00270_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][54] ),
    .QN(_09958_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][55]$_DFFE_PP_  (.D(_00271_),
    .CK(clknet_leaf_287_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][55] ),
    .QN(_09957_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][56]$_DFFE_PP_  (.D(_00272_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][56] ),
    .QN(_09956_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][57]$_DFFE_PP_  (.D(_00273_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][57] ),
    .QN(_09955_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][58]$_DFFE_PP_  (.D(_00274_),
    .CK(clknet_leaf_235_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][58] ),
    .QN(_09954_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][59]$_DFFE_PP_  (.D(_00275_),
    .CK(clknet_leaf_286_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][59] ),
    .QN(_09953_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][5]$_DFFE_PP_  (.D(_00276_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][5] ),
    .QN(_09952_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][60]$_DFFE_PP_  (.D(_00277_),
    .CK(clknet_leaf_287_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][60] ),
    .QN(_09951_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][61]$_DFFE_PP_  (.D(_00278_),
    .CK(clknet_leaf_286_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][61] ),
    .QN(_09950_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][62]$_DFFE_PP_  (.D(_00279_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][62] ),
    .QN(_09949_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][63]$_DFFE_PP_  (.D(_00280_),
    .CK(clknet_leaf_290_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][63] ),
    .QN(_09948_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][6]$_DFFE_PP_  (.D(_00281_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][6] ),
    .QN(_09947_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][7]$_DFFE_PP_  (.D(_00282_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][7] ),
    .QN(_09946_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][8]$_DFFE_PP_  (.D(_00283_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][8] ),
    .QN(_09945_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[2][9]$_DFFE_PP_  (.D(_00284_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[2][9] ),
    .QN(_09944_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][0]$_DFFE_PP_  (.D(_00285_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][0] ),
    .QN(_09943_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][10]$_DFFE_PP_  (.D(_00286_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][10] ),
    .QN(_09942_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][11]$_DFFE_PP_  (.D(_00287_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][11] ),
    .QN(_09941_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][12]$_DFFE_PP_  (.D(_00288_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][12] ),
    .QN(_09940_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][13]$_DFFE_PP_  (.D(_00289_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][13] ),
    .QN(_09939_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][14]$_DFFE_PP_  (.D(_00290_),
    .CK(clknet_leaf_245_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][14] ),
    .QN(_09938_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][15]$_DFFE_PP_  (.D(_00291_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][15] ),
    .QN(_09937_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][16]$_DFFE_PP_  (.D(_00292_),
    .CK(clknet_leaf_237_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][16] ),
    .QN(_09936_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][17]$_DFFE_PP_  (.D(_00293_),
    .CK(clknet_leaf_244_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][17] ),
    .QN(_09935_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][18]$_DFFE_PP_  (.D(_00294_),
    .CK(clknet_leaf_243_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][18] ),
    .QN(_09934_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][19]$_DFFE_PP_  (.D(_00295_),
    .CK(clknet_leaf_238_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][19] ),
    .QN(_09933_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][1]$_DFFE_PP_  (.D(_00296_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][1] ),
    .QN(_09932_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][20]$_DFFE_PP_  (.D(_00297_),
    .CK(clknet_leaf_242_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][20] ),
    .QN(_09931_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][21]$_DFFE_PP_  (.D(_00298_),
    .CK(clknet_leaf_239_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][21] ),
    .QN(_09930_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][22]$_DFFE_PP_  (.D(_00299_),
    .CK(clknet_leaf_240_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][22] ),
    .QN(_09929_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][23]$_DFFE_PP_  (.D(_00300_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][23] ),
    .QN(_09928_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][24]$_DFFE_PP_  (.D(_00301_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][24] ),
    .QN(_09927_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][25]$_DFFE_PP_  (.D(_00302_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][25] ),
    .QN(_09926_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][26]$_DFFE_PP_  (.D(_00303_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][26] ),
    .QN(_09925_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][27]$_DFFE_PP_  (.D(_00304_),
    .CK(clknet_leaf_241_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][27] ),
    .QN(_09924_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][28]$_DFFE_PP_  (.D(_00305_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][28] ),
    .QN(_09923_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][29]$_DFFE_PP_  (.D(_00306_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][29] ),
    .QN(_09922_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][2]$_DFFE_PP_  (.D(_00307_),
    .CK(clknet_leaf_227_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][2] ),
    .QN(_09921_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][30]$_DFFE_PP_  (.D(_00308_),
    .CK(clknet_leaf_229_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][30] ),
    .QN(_09920_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][31]$_DFFE_PP_  (.D(_00309_),
    .CK(clknet_leaf_221_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][31] ),
    .QN(_09919_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][32]$_DFFE_PP_  (.D(_00310_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][32] ),
    .QN(_09918_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][33]$_DFFE_PP_  (.D(_00311_),
    .CK(clknet_leaf_228_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][33] ),
    .QN(_09917_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][34]$_DFFE_PP_  (.D(_00312_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][34] ),
    .QN(_09916_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][35]$_DFFE_PP_  (.D(_00313_),
    .CK(clknet_leaf_222_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][35] ),
    .QN(_09915_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][36]$_DFFE_PP_  (.D(_00314_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][36] ),
    .QN(_09914_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][37]$_DFFE_PP_  (.D(_00315_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][37] ),
    .QN(_09913_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][38]$_DFFE_PP_  (.D(_00316_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][38] ),
    .QN(_09912_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][39]$_DFFE_PP_  (.D(_00317_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][39] ),
    .QN(_09911_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][3]$_DFFE_PP_  (.D(_00318_),
    .CK(clknet_leaf_228_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][3] ),
    .QN(_09910_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][40]$_DFFE_PP_  (.D(_00319_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][40] ),
    .QN(_09909_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][41]$_DFFE_PP_  (.D(_00320_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][41] ),
    .QN(_09908_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][42]$_DFFE_PP_  (.D(_00321_),
    .CK(clknet_leaf_231_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][42] ),
    .QN(_09907_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][43]$_DFFE_PP_  (.D(_00322_),
    .CK(clknet_leaf_208_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][43] ),
    .QN(_09906_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][44]$_DFFE_PP_  (.D(_00323_),
    .CK(clknet_leaf_209_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][44] ),
    .QN(_09905_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][45]$_DFFE_PP_  (.D(_00324_),
    .CK(clknet_leaf_210_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][45] ),
    .QN(_09904_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][46]$_DFFE_PP_  (.D(_00325_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][46] ),
    .QN(_09903_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][47]$_DFFE_PP_  (.D(_00326_),
    .CK(clknet_leaf_207_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][47] ),
    .QN(_09902_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][48]$_DFFE_PP_  (.D(_00327_),
    .CK(clknet_leaf_232_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][48] ),
    .QN(_09901_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][49]$_DFFE_PP_  (.D(_00328_),
    .CK(clknet_leaf_233_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][49] ),
    .QN(_09900_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][4]$_DFFE_PP_  (.D(_00329_),
    .CK(clknet_leaf_235_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][4] ),
    .QN(_09899_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][50]$_DFFE_PP_  (.D(_00330_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][50] ),
    .QN(_09898_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][51]$_DFFE_PP_  (.D(_00331_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][51] ),
    .QN(_09897_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][52]$_DFFE_PP_  (.D(_00332_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][52] ),
    .QN(_09896_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][53]$_DFFE_PP_  (.D(_00333_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][53] ),
    .QN(_09895_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][54]$_DFFE_PP_  (.D(_00334_),
    .CK(clknet_leaf_289_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][54] ),
    .QN(_09894_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][55]$_DFFE_PP_  (.D(_00335_),
    .CK(clknet_leaf_290_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][55] ),
    .QN(_09893_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][56]$_DFFE_PP_  (.D(_00336_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][56] ),
    .QN(_09892_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][57]$_DFFE_PP_  (.D(_00337_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][57] ),
    .QN(_09891_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][58]$_DFFE_PP_  (.D(_00338_),
    .CK(clknet_leaf_234_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][58] ),
    .QN(_09890_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][59]$_DFFE_PP_  (.D(_00339_),
    .CK(clknet_leaf_286_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][59] ),
    .QN(_09889_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][5]$_DFFE_PP_  (.D(_00340_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][5] ),
    .QN(_09888_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][60]$_DFFE_PP_  (.D(_00341_),
    .CK(clknet_leaf_287_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][60] ),
    .QN(_09887_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][61]$_DFFE_PP_  (.D(_00342_),
    .CK(clknet_leaf_288_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][61] ),
    .QN(_09886_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][62]$_DFFE_PP_  (.D(_00343_),
    .CK(clknet_leaf_261_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][62] ),
    .QN(_09885_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][63]$_DFFE_PP_  (.D(_00344_),
    .CK(clknet_leaf_290_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][63] ),
    .QN(_09884_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][6]$_DFFE_PP_  (.D(_00345_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][6] ),
    .QN(_09883_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][7]$_DFFE_PP_  (.D(_00346_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][7] ),
    .QN(_09882_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][8]$_DFFE_PP_  (.D(_00347_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][8] ),
    .QN(_09881_));
 DFF_X1 \dynamic_node_top.east_input.NIB.storage_data_f[3][9]$_DFFE_PP_  (.D(_00348_),
    .CK(clknet_leaf_260_clk),
    .Q(\dynamic_node_top.east_input.NIB.storage_data_f[3][9] ),
    .QN(_09880_));
 DFF_X1 \dynamic_node_top.east_input.NIB.tail_ptr_f[0]$_SDFFE_PP0N_  (.D(_00349_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.tail_ptr_f[0] ),
    .QN(\dynamic_node_top.east_input.NIB.tail_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.east_input.NIB.tail_ptr_f[1]$_SDFFE_PP0N_  (.D(_00350_),
    .CK(clknet_leaf_236_clk),
    .Q(\dynamic_node_top.east_input.NIB.tail_ptr_f[1] ),
    .QN(_10576_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[0]$_SDFF_PP0_  (.D(_00351_),
    .CK(clknet_leaf_177_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[0] ),
    .QN(_10438_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[1]$_SDFF_PP0_  (.D(_00352_),
    .CK(clknet_leaf_177_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[1] ),
    .QN(_10439_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[2]$_SDFF_PP0_  (.D(_00353_),
    .CK(clknet_leaf_174_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[2] ),
    .QN(_09879_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[3]$_SDFF_PP0_  (.D(_00354_),
    .CK(clknet_leaf_174_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[3] ),
    .QN(_09878_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[4]$_SDFF_PP0_  (.D(_00355_),
    .CK(clknet_leaf_174_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[4] ),
    .QN(_09877_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[5]$_SDFF_PP0_  (.D(_00356_),
    .CK(clknet_leaf_174_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[5] ),
    .QN(_09876_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[6]$_SDFF_PP0_  (.D(_00357_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[6] ),
    .QN(_09875_));
 DFF_X1 \dynamic_node_top.east_input.control.count_f[7]$_SDFF_PP0_  (.D(_00358_),
    .CK(clknet_leaf_174_clk),
    .Q(\dynamic_node_top.east_input.control.count_f[7] ),
    .QN(_09874_));
 DFF_X1 \dynamic_node_top.east_input.control.count_one_f$_SDFF_PP0_  (.D(_00359_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.east_input.control.count_one_f ),
    .QN(_10151_));
 DFF_X1 \dynamic_node_top.east_input.control.header_temp$_DFF_P_  (.D(_00000_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.east_input.control.header_last_temp ),
    .QN(_09873_));
 DFF_X1 \dynamic_node_top.east_input.control.tail_last_f$_SDFF_PP0_  (.D(_00360_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.east_input.control.tail_last_f ),
    .QN(_09872_));
 DFF_X1 \dynamic_node_top.east_input.control.thanks_all_f$_SDFF_PP0_  (.D(_00361_),
    .CK(clknet_leaf_175_clk),
    .Q(net626),
    .QN(_10152_));
 DFF_X1 \dynamic_node_top.east_output.control.current_route_f[0]$_DFF_P_  (.D(_00037_),
    .CK(clknet_leaf_159_clk),
    .Q(\dynamic_node_top.east_output.control.current_route_f[0] ),
    .QN(_00045_));
 DFF_X1 \dynamic_node_top.east_output.control.current_route_f[1]$_DFF_P_  (.D(_00038_),
    .CK(clknet_leaf_160_clk),
    .Q(\dynamic_node_top.east_output.control.current_route_f[1] ),
    .QN(_00044_));
 DFF_X1 \dynamic_node_top.east_output.control.current_route_f[2]$_DFF_P_  (.D(_00039_),
    .CK(clknet_leaf_159_clk),
    .Q(\dynamic_node_top.east_output.control.current_route_f[2] ),
    .QN(_00075_));
 DFF_X1 \dynamic_node_top.east_output.control.current_route_f[3]$_DFF_P_  (.D(_00040_),
    .CK(clknet_leaf_159_clk),
    .Q(\dynamic_node_top.east_output.control.current_route_f[3] ),
    .QN(_00076_));
 DFF_X1 \dynamic_node_top.east_output.control.current_route_f[4]$_DFF_P_  (.D(_00041_),
    .CK(clknet_leaf_159_clk),
    .Q(\dynamic_node_top.east_output.control.current_route_f[4] ),
    .QN(_00074_));
 DFF_X2 \dynamic_node_top.east_output.control.planned_f$_SDFF_PP0_  (.D(_00362_),
    .CK(clknet_leaf_160_clk),
    .Q(\dynamic_node_top.east_output.control.planned_f ),
    .QN(_00046_));
 DFF_X2 \dynamic_node_top.east_output.space.count_f[0]$_SDFF_PP0_  (.D(_00363_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.east_output.space.count_f[0] ),
    .QN(_10430_));
 DFF_X2 \dynamic_node_top.east_output.space.count_f[1]$_SDFF_PP0_  (.D(_00364_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.east_output.space.count_f[1] ),
    .QN(_10431_));
 DFF_X1 \dynamic_node_top.east_output.space.count_f[2]$_SDFF_PP1_  (.D(_00365_),
    .CK(clknet_leaf_163_clk),
    .Q(\dynamic_node_top.east_output.space.count_f[2] ),
    .QN(_00057_));
 DFF_X1 \dynamic_node_top.east_output.space.is_one_f$_SDFF_PP0_  (.D(_00366_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.east_output.space.is_one_f ),
    .QN(_09871_));
 DFF_X1 \dynamic_node_top.east_output.space.is_two_or_more_f$_SDFF_PP1_  (.D(_00367_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.east_output.space.is_two_or_more_f ),
    .QN(_09870_));
 DFF_X1 \dynamic_node_top.east_output.space.valid_f$_SDFF_PP0_  (.D(_00368_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.east_output.space.valid_f ),
    .QN(_10427_));
 DFF_X1 \dynamic_node_top.east_output.space.yummy_f$_SDFF_PP0_  (.D(_00369_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.east_output.space.yummy_f ),
    .QN(_10424_));
 DFF_X2 \dynamic_node_top.myChipID_f[0]$_SDFF_PP0_  (.D(_00370_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[0] ),
    .QN(_09869_));
 DFF_X2 \dynamic_node_top.myChipID_f[10]$_SDFF_PP0_  (.D(_00371_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[10] ),
    .QN(_09868_));
 DFF_X1 \dynamic_node_top.myChipID_f[11]$_SDFF_PP0_  (.D(_00372_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[11] ),
    .QN(_09867_));
 DFF_X2 \dynamic_node_top.myChipID_f[12]$_SDFF_PP0_  (.D(_00373_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[12] ),
    .QN(_09866_));
 DFF_X1 \dynamic_node_top.myChipID_f[13]$_SDFF_PP0_  (.D(_00374_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[13] ),
    .QN(_09865_));
 DFF_X1 \dynamic_node_top.myChipID_f[1]$_SDFF_PP0_  (.D(_00375_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[1] ),
    .QN(_09864_));
 DFF_X1 \dynamic_node_top.myChipID_f[2]$_SDFF_PP0_  (.D(_00376_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[2] ),
    .QN(_09863_));
 DFF_X1 \dynamic_node_top.myChipID_f[3]$_SDFF_PP0_  (.D(_00377_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[3] ),
    .QN(_09862_));
 DFF_X2 \dynamic_node_top.myChipID_f[4]$_SDFF_PP0_  (.D(_00378_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[4] ),
    .QN(_09861_));
 DFF_X1 \dynamic_node_top.myChipID_f[5]$_SDFF_PP0_  (.D(_00379_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[5] ),
    .QN(_09860_));
 DFF_X1 \dynamic_node_top.myChipID_f[6]$_SDFF_PP0_  (.D(_00380_),
    .CK(clknet_leaf_48_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[6] ),
    .QN(_09859_));
 DFF_X1 \dynamic_node_top.myChipID_f[7]$_SDFF_PP0_  (.D(_00381_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[7] ),
    .QN(_09858_));
 DFF_X1 \dynamic_node_top.myChipID_f[8]$_SDFF_PP0_  (.D(_00382_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[8] ),
    .QN(_09857_));
 DFF_X1 \dynamic_node_top.myChipID_f[9]$_SDFF_PP0_  (.D(_00383_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.east_input.control.my_chip_id_in[9] ),
    .QN(_09856_));
 DFF_X2 \dynamic_node_top.myLocX_f[0]$_SDFF_PP0_  (.D(_00384_),
    .CK(clknet_leaf_139_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[0] ),
    .QN(_10178_));
 DFF_X2 \dynamic_node_top.myLocX_f[1]$_SDFF_PP0_  (.D(_00385_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[1] ),
    .QN(_09855_));
 DFF_X2 \dynamic_node_top.myLocX_f[2]$_SDFF_PP0_  (.D(_00386_),
    .CK(clknet_leaf_145_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[2] ),
    .QN(_09854_));
 DFF_X2 \dynamic_node_top.myLocX_f[3]$_SDFF_PP0_  (.D(_00387_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[3] ),
    .QN(_09853_));
 DFF_X2 \dynamic_node_top.myLocX_f[4]$_SDFF_PP0_  (.D(_00388_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[4] ),
    .QN(_09852_));
 DFF_X2 \dynamic_node_top.myLocX_f[5]$_SDFF_PP0_  (.D(_00389_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[5] ),
    .QN(_09851_));
 DFF_X2 \dynamic_node_top.myLocX_f[6]$_SDFF_PP0_  (.D(_00390_),
    .CK(clknet_leaf_164_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[6] ),
    .QN(_09850_));
 DFF_X2 \dynamic_node_top.myLocX_f[7]$_SDFF_PP0_  (.D(_00391_),
    .CK(clknet_leaf_164_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_x_in[7] ),
    .QN(_09849_));
 DFF_X2 \dynamic_node_top.myLocY_f[0]$_SDFF_PP0_  (.D(_00392_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[0] ),
    .QN(_10224_));
 DFF_X2 \dynamic_node_top.myLocY_f[1]$_SDFF_PP0_  (.D(_00393_),
    .CK(clknet_leaf_164_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[1] ),
    .QN(_09848_));
 DFF_X2 \dynamic_node_top.myLocY_f[2]$_SDFF_PP0_  (.D(_00394_),
    .CK(clknet_leaf_162_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[2] ),
    .QN(_09847_));
 DFF_X2 \dynamic_node_top.myLocY_f[3]$_SDFF_PP0_  (.D(_00395_),
    .CK(clknet_leaf_162_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[3] ),
    .QN(_09846_));
 DFF_X2 \dynamic_node_top.myLocY_f[4]$_SDFF_PP0_  (.D(_00396_),
    .CK(clknet_leaf_162_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[4] ),
    .QN(_09845_));
 DFF_X2 \dynamic_node_top.myLocY_f[5]$_SDFF_PP0_  (.D(_00397_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[5] ),
    .QN(_09844_));
 DFF_X2 \dynamic_node_top.myLocY_f[6]$_SDFF_PP0_  (.D(_00398_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[6] ),
    .QN(_09843_));
 DFF_X2 \dynamic_node_top.myLocY_f[7]$_SDFF_PP0_  (.D(_00399_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.east_input.control.my_loc_y_in[7] ),
    .QN(_09842_));
 DFF_X1 \dynamic_node_top.north_input.NIB.elements_in_array_f[0]$_SDFFE_PP0N_  (.D(_00400_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.NIB.elements_in_array_f[0] ),
    .QN(\dynamic_node_top.north_input.NIB.elements_in_array_next[0] ));
 DFF_X2 \dynamic_node_top.north_input.NIB.elements_in_array_f[1]$_SDFFE_PP0N_  (.D(_00401_),
    .CK(clknet_leaf_152_clk),
    .Q(\dynamic_node_top.north_input.NIB.elements_in_array_f[1] ),
    .QN(_09841_));
 DFF_X1 \dynamic_node_top.north_input.NIB.elements_in_array_f[2]$_SDFFE_PP0N_  (.D(_00402_),
    .CK(clknet_leaf_152_clk),
    .Q(\dynamic_node_top.north_input.NIB.elements_in_array_f[2] ),
    .QN(_09840_));
 DFF_X1 \dynamic_node_top.north_input.NIB.head_ptr_f[0]$_SDFFE_PP0N_  (.D(_00403_),
    .CK(clknet_leaf_143_clk),
    .Q(\dynamic_node_top.north_input.NIB.head_ptr_f[0] ),
    .QN(\dynamic_node_top.north_input.NIB.head_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.north_input.NIB.head_ptr_f[1]$_SDFFE_PP0N_  (.D(_00088_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.north_input.NIB.head_ptr_f[1] ),
    .QN(_09839_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][0]$_DFFE_PP_  (.D(_00404_),
    .CK(clknet_leaf_293_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][0] ),
    .QN(_09838_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][10]$_DFFE_PP_  (.D(_00405_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][10] ),
    .QN(_09837_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][11]$_DFFE_PP_  (.D(_00406_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][11] ),
    .QN(_09836_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][12]$_DFFE_PP_  (.D(_00407_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][12] ),
    .QN(_09835_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][13]$_DFFE_PP_  (.D(_00408_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][13] ),
    .QN(_09834_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][14]$_DFFE_PP_  (.D(_00409_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][14] ),
    .QN(_09833_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][15]$_DFFE_PP_  (.D(_00410_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][15] ),
    .QN(_09832_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][16]$_DFFE_PP_  (.D(_00411_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][16] ),
    .QN(_09831_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][17]$_DFFE_PP_  (.D(_00412_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][17] ),
    .QN(_09830_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][18]$_DFFE_PP_  (.D(_00413_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][18] ),
    .QN(_09829_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][19]$_DFFE_PP_  (.D(_00414_),
    .CK(clknet_leaf_198_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][19] ),
    .QN(_09828_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][1]$_DFFE_PP_  (.D(_00415_),
    .CK(clknet_leaf_139_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][1] ),
    .QN(_09827_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][20]$_DFFE_PP_  (.D(_00416_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][20] ),
    .QN(_09826_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][21]$_DFFE_PP_  (.D(_00417_),
    .CK(clknet_leaf_139_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][21] ),
    .QN(_09825_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][22]$_DFFE_PP_  (.D(_00418_),
    .CK(clknet_leaf_152_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][22] ),
    .QN(_09824_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][23]$_DFFE_PP_  (.D(_00419_),
    .CK(clknet_leaf_151_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][23] ),
    .QN(_09823_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][24]$_DFFE_PP_  (.D(_00420_),
    .CK(clknet_leaf_151_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][24] ),
    .QN(_09822_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][25]$_DFFE_PP_  (.D(_00421_),
    .CK(clknet_leaf_152_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][25] ),
    .QN(_09821_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][26]$_DFFE_PP_  (.D(_00422_),
    .CK(clknet_leaf_150_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][26] ),
    .QN(_09820_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][27]$_DFFE_PP_  (.D(_00423_),
    .CK(clknet_leaf_150_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][27] ),
    .QN(_09819_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][28]$_DFFE_PP_  (.D(_00424_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][28] ),
    .QN(_09818_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][29]$_DFFE_PP_  (.D(_00425_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][29] ),
    .QN(_09817_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][2]$_DFFE_PP_  (.D(_00426_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][2] ),
    .QN(_09816_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][30]$_DFFE_PP_  (.D(_00427_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][30] ),
    .QN(_09815_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][31]$_DFFE_PP_  (.D(_00428_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][31] ),
    .QN(_09814_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][32]$_DFFE_PP_  (.D(_00429_),
    .CK(clknet_leaf_145_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][32] ),
    .QN(_09813_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][33]$_DFFE_PP_  (.D(_00430_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][33] ),
    .QN(_09812_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][34]$_DFFE_PP_  (.D(_00431_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][34] ),
    .QN(_09811_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][35]$_DFFE_PP_  (.D(_00432_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][35] ),
    .QN(_09810_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][36]$_DFFE_PP_  (.D(_00433_),
    .CK(clknet_leaf_145_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][36] ),
    .QN(_09809_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][37]$_DFFE_PP_  (.D(_00434_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][37] ),
    .QN(_09808_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][38]$_DFFE_PP_  (.D(_00435_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][38] ),
    .QN(_09807_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][39]$_DFFE_PP_  (.D(_00436_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][39] ),
    .QN(_09806_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][3]$_DFFE_PP_  (.D(_00437_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][3] ),
    .QN(_09805_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][40]$_DFFE_PP_  (.D(_00438_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][40] ),
    .QN(_09804_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][41]$_DFFE_PP_  (.D(_00439_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][41] ),
    .QN(_09803_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][42]$_DFFE_PP_  (.D(_00440_),
    .CK(clknet_leaf_124_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][42] ),
    .QN(_09802_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][43]$_DFFE_PP_  (.D(_00441_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][43] ),
    .QN(_09801_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][44]$_DFFE_PP_  (.D(_00442_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][44] ),
    .QN(_09800_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][45]$_DFFE_PP_  (.D(_00443_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][45] ),
    .QN(_09799_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][46]$_DFFE_PP_  (.D(_00444_),
    .CK(clknet_leaf_129_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][46] ),
    .QN(_09798_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][47]$_DFFE_PP_  (.D(_00445_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][47] ),
    .QN(_09797_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][48]$_DFFE_PP_  (.D(_00446_),
    .CK(clknet_leaf_129_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][48] ),
    .QN(_09796_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][49]$_DFFE_PP_  (.D(_00447_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][49] ),
    .QN(_09795_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][4]$_DFFE_PP_  (.D(_00448_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][4] ),
    .QN(_09794_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][50]$_DFFE_PP_  (.D(_00449_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][50] ),
    .QN(_09793_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][51]$_DFFE_PP_  (.D(_00450_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][51] ),
    .QN(_09792_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][52]$_DFFE_PP_  (.D(_00451_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][52] ),
    .QN(_09791_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][53]$_DFFE_PP_  (.D(_00452_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][53] ),
    .QN(_09790_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][54]$_DFFE_PP_  (.D(_00453_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][54] ),
    .QN(_09789_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][55]$_DFFE_PP_  (.D(_00454_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][55] ),
    .QN(_09788_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][56]$_DFFE_PP_  (.D(_00455_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][56] ),
    .QN(_09787_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][57]$_DFFE_PP_  (.D(_00456_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][57] ),
    .QN(_09786_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][58]$_DFFE_PP_  (.D(_00457_),
    .CK(clknet_leaf_204_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][58] ),
    .QN(_09785_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][59]$_DFFE_PP_  (.D(_00458_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][59] ),
    .QN(_09784_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][5]$_DFFE_PP_  (.D(_00459_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][5] ),
    .QN(_09783_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][60]$_DFFE_PP_  (.D(_00460_),
    .CK(clknet_leaf_199_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][60] ),
    .QN(_09782_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][61]$_DFFE_PP_  (.D(_00461_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][61] ),
    .QN(_09781_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][62]$_DFFE_PP_  (.D(_00462_),
    .CK(clknet_leaf_196_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][62] ),
    .QN(_09780_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][63]$_DFFE_PP_  (.D(_00463_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][63] ),
    .QN(_09779_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][6]$_DFFE_PP_  (.D(_00464_),
    .CK(clknet_leaf_301_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][6] ),
    .QN(_09778_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][7]$_DFFE_PP_  (.D(_00465_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][7] ),
    .QN(_09777_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][8]$_DFFE_PP_  (.D(_00466_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][8] ),
    .QN(_09776_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[0][9]$_DFFE_PP_  (.D(_00467_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[0][9] ),
    .QN(_09775_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][0]$_DFFE_PP_  (.D(_00468_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][0] ),
    .QN(_09774_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][10]$_DFFE_PP_  (.D(_00469_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][10] ),
    .QN(_09773_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][11]$_DFFE_PP_  (.D(_00470_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][11] ),
    .QN(_09772_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][12]$_DFFE_PP_  (.D(_00471_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][12] ),
    .QN(_09771_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][13]$_DFFE_PP_  (.D(_00472_),
    .CK(clknet_leaf_291_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][13] ),
    .QN(_09770_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][14]$_DFFE_PP_  (.D(_00473_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][14] ),
    .QN(_09769_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][15]$_DFFE_PP_  (.D(_00474_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][15] ),
    .QN(_09768_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][16]$_DFFE_PP_  (.D(_00475_),
    .CK(clknet_leaf_291_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][16] ),
    .QN(_09767_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][17]$_DFFE_PP_  (.D(_00476_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][17] ),
    .QN(_09766_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][18]$_DFFE_PP_  (.D(_00477_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][18] ),
    .QN(_09765_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][19]$_DFFE_PP_  (.D(_00478_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][19] ),
    .QN(_09764_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][1]$_DFFE_PP_  (.D(_00479_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][1] ),
    .QN(_09763_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][20]$_DFFE_PP_  (.D(_00480_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][20] ),
    .QN(_09762_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][21]$_DFFE_PP_  (.D(_00481_),
    .CK(clknet_leaf_139_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][21] ),
    .QN(_09761_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][22]$_DFFE_PP_  (.D(_00482_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][22] ),
    .QN(_09760_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][23]$_DFFE_PP_  (.D(_00483_),
    .CK(clknet_leaf_151_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][23] ),
    .QN(_09759_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][24]$_DFFE_PP_  (.D(_00484_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][24] ),
    .QN(_09758_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][25]$_DFFE_PP_  (.D(_00485_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][25] ),
    .QN(_09757_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][26]$_DFFE_PP_  (.D(_00486_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][26] ),
    .QN(_09756_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][27]$_DFFE_PP_  (.D(_00487_),
    .CK(clknet_leaf_150_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][27] ),
    .QN(_09755_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][28]$_DFFE_PP_  (.D(_00488_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][28] ),
    .QN(_09754_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][29]$_DFFE_PP_  (.D(_00489_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][29] ),
    .QN(_09753_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][2]$_DFFE_PP_  (.D(_00490_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][2] ),
    .QN(_09752_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][30]$_DFFE_PP_  (.D(_00491_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][30] ),
    .QN(_09751_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][31]$_DFFE_PP_  (.D(_00492_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][31] ),
    .QN(_09750_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][32]$_DFFE_PP_  (.D(_00493_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][32] ),
    .QN(_09749_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][33]$_DFFE_PP_  (.D(_00494_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][33] ),
    .QN(_09748_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][34]$_DFFE_PP_  (.D(_00495_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][34] ),
    .QN(_09747_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][35]$_DFFE_PP_  (.D(_00496_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][35] ),
    .QN(_09746_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][36]$_DFFE_PP_  (.D(_00497_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][36] ),
    .QN(_09745_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][37]$_DFFE_PP_  (.D(_00498_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][37] ),
    .QN(_09744_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][38]$_DFFE_PP_  (.D(_00499_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][38] ),
    .QN(_09743_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][39]$_DFFE_PP_  (.D(_00500_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][39] ),
    .QN(_09742_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][3]$_DFFE_PP_  (.D(_00501_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][3] ),
    .QN(_09741_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][40]$_DFFE_PP_  (.D(_00502_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][40] ),
    .QN(_09740_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][41]$_DFFE_PP_  (.D(_00503_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][41] ),
    .QN(_09739_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][42]$_DFFE_PP_  (.D(_00504_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][42] ),
    .QN(_09738_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][43]$_DFFE_PP_  (.D(_00505_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][43] ),
    .QN(_09737_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][44]$_DFFE_PP_  (.D(_00506_),
    .CK(clknet_leaf_124_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][44] ),
    .QN(_09736_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][45]$_DFFE_PP_  (.D(_00507_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][45] ),
    .QN(_09735_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][46]$_DFFE_PP_  (.D(_00508_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][46] ),
    .QN(_09734_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][47]$_DFFE_PP_  (.D(_00509_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][47] ),
    .QN(_09733_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][48]$_DFFE_PP_  (.D(_00510_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][48] ),
    .QN(_09732_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][49]$_DFFE_PP_  (.D(_00511_),
    .CK(clknet_leaf_198_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][49] ),
    .QN(_09731_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][4]$_DFFE_PP_  (.D(_00512_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][4] ),
    .QN(_09730_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][50]$_DFFE_PP_  (.D(_00513_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][50] ),
    .QN(_09729_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][51]$_DFFE_PP_  (.D(_00514_),
    .CK(clknet_leaf_198_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][51] ),
    .QN(_09728_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][52]$_DFFE_PP_  (.D(_00515_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][52] ),
    .QN(_09727_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][53]$_DFFE_PP_  (.D(_00516_),
    .CK(clknet_leaf_199_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][53] ),
    .QN(_09726_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][54]$_DFFE_PP_  (.D(_00517_),
    .CK(clknet_leaf_199_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][54] ),
    .QN(_09725_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][55]$_DFFE_PP_  (.D(_00518_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][55] ),
    .QN(_09724_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][56]$_DFFE_PP_  (.D(_00519_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][56] ),
    .QN(_09723_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][57]$_DFFE_PP_  (.D(_00520_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][57] ),
    .QN(_09722_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][58]$_DFFE_PP_  (.D(_00521_),
    .CK(clknet_leaf_204_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][58] ),
    .QN(_09721_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][59]$_DFFE_PP_  (.D(_00522_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][59] ),
    .QN(_09720_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][5]$_DFFE_PP_  (.D(_00523_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][5] ),
    .QN(_09719_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][60]$_DFFE_PP_  (.D(_00524_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][60] ),
    .QN(_09718_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][61]$_DFFE_PP_  (.D(_00525_),
    .CK(clknet_leaf_206_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][61] ),
    .QN(_09717_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][62]$_DFFE_PP_  (.D(_00526_),
    .CK(clknet_leaf_206_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][62] ),
    .QN(_09716_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][63]$_DFFE_PP_  (.D(_00527_),
    .CK(clknet_leaf_204_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][63] ),
    .QN(_09715_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][6]$_DFFE_PP_  (.D(_00528_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][6] ),
    .QN(_09714_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][7]$_DFFE_PP_  (.D(_00529_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][7] ),
    .QN(_09713_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][8]$_DFFE_PP_  (.D(_00530_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][8] ),
    .QN(_09712_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[1][9]$_DFFE_PP_  (.D(_00531_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[1][9] ),
    .QN(_09711_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][0]$_DFFE_PP_  (.D(_00532_),
    .CK(clknet_leaf_293_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][0] ),
    .QN(_09710_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][10]$_DFFE_PP_  (.D(_00533_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][10] ),
    .QN(_09709_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][11]$_DFFE_PP_  (.D(_00534_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][11] ),
    .QN(_09708_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][12]$_DFFE_PP_  (.D(_00535_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][12] ),
    .QN(_09707_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][13]$_DFFE_PP_  (.D(_00536_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][13] ),
    .QN(_09706_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][14]$_DFFE_PP_  (.D(_00537_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][14] ),
    .QN(_09705_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][15]$_DFFE_PP_  (.D(_00538_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][15] ),
    .QN(_09704_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][16]$_DFFE_PP_  (.D(_00539_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][16] ),
    .QN(_09703_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][17]$_DFFE_PP_  (.D(_00540_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][17] ),
    .QN(_09702_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][18]$_DFFE_PP_  (.D(_00541_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][18] ),
    .QN(_09701_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][19]$_DFFE_PP_  (.D(_00542_),
    .CK(clknet_leaf_198_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][19] ),
    .QN(_09700_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][1]$_DFFE_PP_  (.D(_00543_),
    .CK(clknet_leaf_140_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][1] ),
    .QN(_09699_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][20]$_DFFE_PP_  (.D(_00544_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][20] ),
    .QN(_09698_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][21]$_DFFE_PP_  (.D(_00545_),
    .CK(clknet_leaf_139_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][21] ),
    .QN(_09697_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][22]$_DFFE_PP_  (.D(_00546_),
    .CK(clknet_leaf_151_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][22] ),
    .QN(_09696_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][23]$_DFFE_PP_  (.D(_00547_),
    .CK(clknet_leaf_151_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][23] ),
    .QN(_09695_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][24]$_DFFE_PP_  (.D(_00548_),
    .CK(clknet_leaf_151_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][24] ),
    .QN(_09694_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][25]$_DFFE_PP_  (.D(_00549_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][25] ),
    .QN(_09693_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][26]$_DFFE_PP_  (.D(_00550_),
    .CK(clknet_leaf_150_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][26] ),
    .QN(_09692_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][27]$_DFFE_PP_  (.D(_00551_),
    .CK(clknet_leaf_150_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][27] ),
    .QN(_09691_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][28]$_DFFE_PP_  (.D(_00552_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][28] ),
    .QN(_09690_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][29]$_DFFE_PP_  (.D(_00553_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][29] ),
    .QN(_09689_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][2]$_DFFE_PP_  (.D(_00554_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][2] ),
    .QN(_09688_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][30]$_DFFE_PP_  (.D(_00555_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][30] ),
    .QN(_09687_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][31]$_DFFE_PP_  (.D(_00556_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][31] ),
    .QN(_09686_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][32]$_DFFE_PP_  (.D(_00557_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][32] ),
    .QN(_09685_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][33]$_DFFE_PP_  (.D(_00558_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][33] ),
    .QN(_09684_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][34]$_DFFE_PP_  (.D(_00559_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][34] ),
    .QN(_09683_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][35]$_DFFE_PP_  (.D(_00560_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][35] ),
    .QN(_09682_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][36]$_DFFE_PP_  (.D(_00561_),
    .CK(clknet_leaf_145_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][36] ),
    .QN(_09681_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][37]$_DFFE_PP_  (.D(_00562_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][37] ),
    .QN(_09680_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][38]$_DFFE_PP_  (.D(_00563_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][38] ),
    .QN(_09679_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][39]$_DFFE_PP_  (.D(_00564_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][39] ),
    .QN(_09678_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][3]$_DFFE_PP_  (.D(_00565_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][3] ),
    .QN(_09677_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][40]$_DFFE_PP_  (.D(_00566_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][40] ),
    .QN(_09676_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][41]$_DFFE_PP_  (.D(_00567_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][41] ),
    .QN(_09675_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][42]$_DFFE_PP_  (.D(_00568_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][42] ),
    .QN(_09674_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][43]$_DFFE_PP_  (.D(_00569_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][43] ),
    .QN(_09673_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][44]$_DFFE_PP_  (.D(_00570_),
    .CK(clknet_leaf_124_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][44] ),
    .QN(_09672_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][45]$_DFFE_PP_  (.D(_00571_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][45] ),
    .QN(_09671_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][46]$_DFFE_PP_  (.D(_00572_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][46] ),
    .QN(_09670_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][47]$_DFFE_PP_  (.D(_00573_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][47] ),
    .QN(_09669_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][48]$_DFFE_PP_  (.D(_00574_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][48] ),
    .QN(_09668_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][49]$_DFFE_PP_  (.D(_00575_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][49] ),
    .QN(_09667_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][4]$_DFFE_PP_  (.D(_00576_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][4] ),
    .QN(_09666_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][50]$_DFFE_PP_  (.D(_00577_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][50] ),
    .QN(_09665_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][51]$_DFFE_PP_  (.D(_00578_),
    .CK(clknet_leaf_199_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][51] ),
    .QN(_09664_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][52]$_DFFE_PP_  (.D(_00579_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][52] ),
    .QN(_09663_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][53]$_DFFE_PP_  (.D(_00580_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][53] ),
    .QN(_09662_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][54]$_DFFE_PP_  (.D(_00581_),
    .CK(clknet_leaf_196_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][54] ),
    .QN(_09661_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][55]$_DFFE_PP_  (.D(_00582_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][55] ),
    .QN(_09660_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][56]$_DFFE_PP_  (.D(_00583_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][56] ),
    .QN(_09659_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][57]$_DFFE_PP_  (.D(_00584_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][57] ),
    .QN(_09658_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][58]$_DFFE_PP_  (.D(_00585_),
    .CK(clknet_leaf_204_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][58] ),
    .QN(_09657_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][59]$_DFFE_PP_  (.D(_00586_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][59] ),
    .QN(_09656_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][5]$_DFFE_PP_  (.D(_00587_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][5] ),
    .QN(_09655_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][60]$_DFFE_PP_  (.D(_00588_),
    .CK(clknet_leaf_199_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][60] ),
    .QN(_09654_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][61]$_DFFE_PP_  (.D(_00589_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][61] ),
    .QN(_09653_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][62]$_DFFE_PP_  (.D(_00590_),
    .CK(clknet_leaf_196_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][62] ),
    .QN(_09652_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][63]$_DFFE_PP_  (.D(_00591_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][63] ),
    .QN(_09651_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][6]$_DFFE_PP_  (.D(_00592_),
    .CK(clknet_leaf_301_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][6] ),
    .QN(_09650_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][7]$_DFFE_PP_  (.D(_00593_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][7] ),
    .QN(_09649_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][8]$_DFFE_PP_  (.D(_00594_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][8] ),
    .QN(_09648_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[2][9]$_DFFE_PP_  (.D(_00595_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[2][9] ),
    .QN(_09647_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][0]$_DFFE_PP_  (.D(_00596_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][0] ),
    .QN(_09646_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][10]$_DFFE_PP_  (.D(_00597_),
    .CK(clknet_leaf_298_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][10] ),
    .QN(_09645_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][11]$_DFFE_PP_  (.D(_00598_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][11] ),
    .QN(_09644_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][12]$_DFFE_PP_  (.D(_00599_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][12] ),
    .QN(_09643_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][13]$_DFFE_PP_  (.D(_00600_),
    .CK(clknet_leaf_291_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][13] ),
    .QN(_09642_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][14]$_DFFE_PP_  (.D(_00601_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][14] ),
    .QN(_09641_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][15]$_DFFE_PP_  (.D(_00602_),
    .CK(clknet_leaf_295_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][15] ),
    .QN(_09640_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][16]$_DFFE_PP_  (.D(_00603_),
    .CK(clknet_leaf_291_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][16] ),
    .QN(_09639_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][17]$_DFFE_PP_  (.D(_00604_),
    .CK(clknet_leaf_297_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][17] ),
    .QN(_09638_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][18]$_DFFE_PP_  (.D(_00605_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][18] ),
    .QN(_09637_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][19]$_DFFE_PP_  (.D(_00606_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][19] ),
    .QN(_09636_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][1]$_DFFE_PP_  (.D(_00607_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][1] ),
    .QN(_09635_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][20]$_DFFE_PP_  (.D(_00608_),
    .CK(clknet_leaf_134_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][20] ),
    .QN(_09634_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][21]$_DFFE_PP_  (.D(_00609_),
    .CK(clknet_leaf_139_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][21] ),
    .QN(_09633_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][22]$_DFFE_PP_  (.D(_00610_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][22] ),
    .QN(_09632_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][23]$_DFFE_PP_  (.D(_00611_),
    .CK(clknet_leaf_150_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][23] ),
    .QN(_09631_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][24]$_DFFE_PP_  (.D(_00612_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][24] ),
    .QN(_09630_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][25]$_DFFE_PP_  (.D(_00613_),
    .CK(clknet_leaf_149_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][25] ),
    .QN(_09629_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][26]$_DFFE_PP_  (.D(_00614_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][26] ),
    .QN(_09628_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][27]$_DFFE_PP_  (.D(_00615_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][27] ),
    .QN(_09627_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][28]$_DFFE_PP_  (.D(_00616_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][28] ),
    .QN(_09626_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][29]$_DFFE_PP_  (.D(_00617_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][29] ),
    .QN(_09625_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][2]$_DFFE_PP_  (.D(_00618_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][2] ),
    .QN(_09624_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][30]$_DFFE_PP_  (.D(_00619_),
    .CK(clknet_leaf_147_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][30] ),
    .QN(_09623_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][31]$_DFFE_PP_  (.D(_00620_),
    .CK(clknet_leaf_144_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][31] ),
    .QN(_09622_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][32]$_DFFE_PP_  (.D(_00621_),
    .CK(clknet_leaf_146_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][32] ),
    .QN(_09621_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][33]$_DFFE_PP_  (.D(_00622_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][33] ),
    .QN(_09620_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][34]$_DFFE_PP_  (.D(_00623_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][34] ),
    .QN(_09619_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][35]$_DFFE_PP_  (.D(_00624_),
    .CK(clknet_leaf_137_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][35] ),
    .QN(_09618_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][36]$_DFFE_PP_  (.D(_00625_),
    .CK(clknet_leaf_138_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][36] ),
    .QN(_09617_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][37]$_DFFE_PP_  (.D(_00626_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][37] ),
    .QN(_09616_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][38]$_DFFE_PP_  (.D(_00627_),
    .CK(clknet_leaf_123_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][38] ),
    .QN(_09615_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][39]$_DFFE_PP_  (.D(_00628_),
    .CK(clknet_leaf_122_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][39] ),
    .QN(_09614_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][3]$_DFFE_PP_  (.D(_00629_),
    .CK(clknet_leaf_136_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][3] ),
    .QN(_09613_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][40]$_DFFE_PP_  (.D(_00630_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][40] ),
    .QN(_09612_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][41]$_DFFE_PP_  (.D(_00631_),
    .CK(clknet_leaf_135_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][41] ),
    .QN(_09611_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][42]$_DFFE_PP_  (.D(_00632_),
    .CK(clknet_leaf_124_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][42] ),
    .QN(_09610_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][43]$_DFFE_PP_  (.D(_00633_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][43] ),
    .QN(_09609_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][44]$_DFFE_PP_  (.D(_00634_),
    .CK(clknet_leaf_124_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][44] ),
    .QN(_09608_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][45]$_DFFE_PP_  (.D(_00635_),
    .CK(clknet_leaf_124_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][45] ),
    .QN(_09607_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][46]$_DFFE_PP_  (.D(_00636_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][46] ),
    .QN(_09606_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][47]$_DFFE_PP_  (.D(_00637_),
    .CK(clknet_leaf_133_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][47] ),
    .QN(_09605_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][48]$_DFFE_PP_  (.D(_00638_),
    .CK(clknet_leaf_132_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][48] ),
    .QN(_09604_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][49]$_DFFE_PP_  (.D(_00639_),
    .CK(clknet_leaf_198_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][49] ),
    .QN(_09603_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][4]$_DFFE_PP_  (.D(_00640_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][4] ),
    .QN(_09602_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][50]$_DFFE_PP_  (.D(_00641_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][50] ),
    .QN(_09601_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][51]$_DFFE_PP_  (.D(_00642_),
    .CK(clknet_leaf_198_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][51] ),
    .QN(_09600_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][52]$_DFFE_PP_  (.D(_00643_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][52] ),
    .QN(_09599_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][53]$_DFFE_PP_  (.D(_00644_),
    .CK(clknet_leaf_199_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][53] ),
    .QN(_09598_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][54]$_DFFE_PP_  (.D(_00645_),
    .CK(clknet_leaf_197_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][54] ),
    .QN(_09597_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][55]$_DFFE_PP_  (.D(_00646_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][55] ),
    .QN(_09596_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][56]$_DFFE_PP_  (.D(_00647_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][56] ),
    .QN(_09595_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][57]$_DFFE_PP_  (.D(_00648_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][57] ),
    .QN(_09594_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][58]$_DFFE_PP_  (.D(_00649_),
    .CK(clknet_leaf_204_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][58] ),
    .QN(_09593_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][59]$_DFFE_PP_  (.D(_00650_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][59] ),
    .QN(_09592_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][5]$_DFFE_PP_  (.D(_00651_),
    .CK(clknet_leaf_205_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][5] ),
    .QN(_09591_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][60]$_DFFE_PP_  (.D(_00652_),
    .CK(clknet_leaf_203_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][60] ),
    .QN(_09590_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][61]$_DFFE_PP_  (.D(_00653_),
    .CK(clknet_leaf_206_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][61] ),
    .QN(_09589_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][62]$_DFFE_PP_  (.D(_00654_),
    .CK(clknet_leaf_206_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][62] ),
    .QN(_09588_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][63]$_DFFE_PP_  (.D(_00655_),
    .CK(clknet_leaf_204_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][63] ),
    .QN(_09587_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][6]$_DFFE_PP_  (.D(_00656_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][6] ),
    .QN(_09586_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][7]$_DFFE_PP_  (.D(_00657_),
    .CK(clknet_leaf_202_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][7] ),
    .QN(_09585_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][8]$_DFFE_PP_  (.D(_00658_),
    .CK(clknet_leaf_299_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][8] ),
    .QN(_09584_));
 DFF_X1 \dynamic_node_top.north_input.NIB.storage_data_f[3][9]$_DFFE_PP_  (.D(_00659_),
    .CK(clknet_leaf_200_clk),
    .Q(\dynamic_node_top.north_input.NIB.storage_data_f[3][9] ),
    .QN(_09583_));
 DFF_X1 \dynamic_node_top.north_input.NIB.tail_ptr_f[0]$_SDFFE_PP0N_  (.D(_00660_),
    .CK(clknet_leaf_145_clk),
    .Q(\dynamic_node_top.north_input.NIB.tail_ptr_f[0] ),
    .QN(\dynamic_node_top.north_input.NIB.tail_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.north_input.NIB.tail_ptr_f[1]$_SDFFE_PP0N_  (.D(_00661_),
    .CK(clknet_leaf_145_clk),
    .Q(\dynamic_node_top.north_input.NIB.tail_ptr_f[1] ),
    .QN(_10584_));
 DFF_X1 \dynamic_node_top.north_input.NIB.yummy_out_f$_SDFF_PP0_  (.D(_00662_),
    .CK(clknet_leaf_152_clk),
    .Q(net627),
    .QN(_09582_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[0]$_SDFF_PP0_  (.D(_00663_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[0] ),
    .QN(_10420_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[1]$_SDFF_PP0_  (.D(_00664_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[1] ),
    .QN(_10421_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[2]$_SDFF_PP0_  (.D(_00665_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[2] ),
    .QN(_09581_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[3]$_SDFF_PP0_  (.D(_00666_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[3] ),
    .QN(_09580_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[4]$_SDFF_PP0_  (.D(_00667_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[4] ),
    .QN(_09579_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[5]$_SDFF_PP0_  (.D(_00668_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[5] ),
    .QN(_09578_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[6]$_SDFF_PP0_  (.D(_00669_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[6] ),
    .QN(_09577_));
 DFF_X1 \dynamic_node_top.north_input.control.count_f[7]$_SDFF_PP0_  (.D(_00670_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.north_input.control.count_f[7] ),
    .QN(_09576_));
 DFF_X1 \dynamic_node_top.north_input.control.count_one_f$_SDFF_PP0_  (.D(_00671_),
    .CK(clknet_leaf_158_clk),
    .Q(\dynamic_node_top.north_input.control.count_one_f ),
    .QN(_10153_));
 DFF_X1 \dynamic_node_top.north_input.control.header_temp$_DFF_P_  (.D(_00001_),
    .CK(clknet_leaf_143_clk),
    .Q(\dynamic_node_top.north_input.control.header_last_temp ),
    .QN(_09575_));
 DFF_X1 \dynamic_node_top.north_input.control.tail_last_f$_SDFF_PP0_  (.D(_00672_),
    .CK(clknet_leaf_153_clk),
    .Q(\dynamic_node_top.north_input.control.tail_last_f ),
    .QN(_10154_));
 DFF_X1 \dynamic_node_top.north_output.control.current_route_f[0]$_DFF_P_  (.D(_00017_),
    .CK(clknet_leaf_158_clk),
    .Q(\dynamic_node_top.north_output.control.current_route_f[0] ),
    .QN(_00042_));
 DFF_X1 \dynamic_node_top.north_output.control.current_route_f[1]$_DFF_P_  (.D(_00018_),
    .CK(clknet_leaf_157_clk),
    .Q(\dynamic_node_top.north_output.control.current_route_f[1] ),
    .QN(_10155_));
 DFF_X1 \dynamic_node_top.north_output.control.current_route_f[2]$_DFF_P_  (.D(_00019_),
    .CK(clknet_leaf_154_clk),
    .Q(\dynamic_node_top.north_output.control.current_route_f[2] ),
    .QN(_00072_));
 DFF_X1 \dynamic_node_top.north_output.control.current_route_f[3]$_DFF_P_  (.D(_00020_),
    .CK(clknet_leaf_157_clk),
    .Q(\dynamic_node_top.north_output.control.current_route_f[3] ),
    .QN(_00073_));
 DFF_X1 \dynamic_node_top.north_output.control.current_route_f[4]$_DFF_P_  (.D(_00021_),
    .CK(clknet_leaf_157_clk),
    .Q(\dynamic_node_top.north_output.control.current_route_f[4] ),
    .QN(_00071_));
 DFF_X1 \dynamic_node_top.north_output.control.planned_f$_SDFF_PP0_  (.D(_00673_),
    .CK(clknet_leaf_154_clk),
    .Q(\dynamic_node_top.north_output.control.planned_f ),
    .QN(_00043_));
 DFF_X2 \dynamic_node_top.north_output.space.count_f[0]$_SDFF_PP0_  (.D(_00674_),
    .CK(clknet_leaf_152_clk),
    .Q(\dynamic_node_top.north_output.space.count_f[0] ),
    .QN(_10541_));
 DFF_X2 \dynamic_node_top.north_output.space.count_f[1]$_SDFF_PP0_  (.D(_00675_),
    .CK(clknet_leaf_152_clk),
    .Q(\dynamic_node_top.north_output.space.count_f[1] ),
    .QN(_10542_));
 DFF_X1 \dynamic_node_top.north_output.space.count_f[2]$_SDFF_PP1_  (.D(_00676_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.north_output.space.count_f[2] ),
    .QN(_00061_));
 DFF_X1 \dynamic_node_top.north_output.space.is_one_f$_SDFF_PP0_  (.D(_00677_),
    .CK(clknet_leaf_154_clk),
    .Q(\dynamic_node_top.north_output.space.is_one_f ),
    .QN(_09574_));
 DFF_X1 \dynamic_node_top.north_output.space.is_two_or_more_f$_SDFF_PP1_  (.D(_00678_),
    .CK(clknet_leaf_154_clk),
    .Q(\dynamic_node_top.north_output.space.is_two_or_more_f ),
    .QN(_09573_));
 DFF_X1 \dynamic_node_top.north_output.space.valid_f$_SDFF_PP0_  (.D(_00679_),
    .CK(clknet_leaf_154_clk),
    .Q(\dynamic_node_top.north_output.space.valid_f ),
    .QN(_10538_));
 DFF_X1 \dynamic_node_top.north_output.space.yummy_f$_SDFF_PP0_  (.D(_00680_),
    .CK(clknet_leaf_154_clk),
    .Q(\dynamic_node_top.north_output.space.yummy_f ),
    .QN(_10535_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.elements_in_array_f[0]$_SDFFE_PP0N_  (.D(_00681_),
    .CK(clknet_leaf_108_clk),
    .Q(\dynamic_node_top.proc_input.NIB.elements_in_array_f[0] ),
    .QN(\dynamic_node_top.proc_input.NIB.elements_in_array_next[0] ));
 DFF_X2 \dynamic_node_top.proc_input.NIB.elements_in_array_f[1]$_SDFFE_PP0N_  (.D(_00682_),
    .CK(clknet_leaf_108_clk),
    .Q(\dynamic_node_top.proc_input.NIB.elements_in_array_f[1] ),
    .QN(_10168_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.elements_in_array_f[2]$_SDFFE_PP0N_  (.D(_00683_),
    .CK(clknet_leaf_108_clk),
    .Q(\dynamic_node_top.proc_input.NIB.elements_in_array_f[2] ),
    .QN(_09572_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.elements_in_array_f[3]$_SDFFE_PP0N_  (.D(_00684_),
    .CK(clknet_leaf_108_clk),
    .Q(\dynamic_node_top.proc_input.NIB.elements_in_array_f[3] ),
    .QN(_09571_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.elements_in_array_f[4]$_SDFFE_PP0N_  (.D(_00685_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.proc_input.NIB.elements_in_array_f[4] ),
    .QN(_09570_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.head_ptr_f[0]$_SDFFE_PP0N_  (.D(_00686_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.proc_input.NIB.head_ptr_f[0] ),
    .QN(\dynamic_node_top.proc_input.NIB.head_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.proc_input.NIB.head_ptr_f[1]$_SDFFE_PP0N_  (.D(_00084_),
    .CK(clknet_leaf_125_clk),
    .Q(\dynamic_node_top.proc_input.NIB.head_ptr_f[1] ),
    .QN(_09569_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.head_ptr_f[2]$_SDFFE_PP0N_  (.D(_00085_),
    .CK(clknet_leaf_128_clk),
    .Q(\dynamic_node_top.proc_input.NIB.head_ptr_f[2] ),
    .QN(_09568_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.head_ptr_f[3]$_SDFFE_PP0N_  (.D(_00086_),
    .CK(clknet_leaf_128_clk),
    .Q(\dynamic_node_top.proc_input.NIB.head_ptr_f[3] ),
    .QN(_09567_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][0]$_DFFE_PP_  (.D(_00687_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][0] ),
    .QN(_09566_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][10]$_DFFE_PP_  (.D(_00688_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][10] ),
    .QN(_09565_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][11]$_DFFE_PP_  (.D(_00689_),
    .CK(clknet_leaf_324_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][11] ),
    .QN(_09564_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][12]$_DFFE_PP_  (.D(_00690_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][12] ),
    .QN(_09563_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][13]$_DFFE_PP_  (.D(_00691_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][13] ),
    .QN(_09562_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][14]$_DFFE_PP_  (.D(_00692_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][14] ),
    .QN(_09561_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][15]$_DFFE_PP_  (.D(_00693_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][15] ),
    .QN(_09560_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][16]$_DFFE_PP_  (.D(_00694_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][16] ),
    .QN(_09559_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][17]$_DFFE_PP_  (.D(_00695_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][17] ),
    .QN(_09558_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][18]$_DFFE_PP_  (.D(_00696_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][18] ),
    .QN(_09557_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][19]$_DFFE_PP_  (.D(_00697_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][19] ),
    .QN(_09556_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][1]$_DFFE_PP_  (.D(_00698_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][1] ),
    .QN(_09555_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][20]$_DFFE_PP_  (.D(_00699_),
    .CK(clknet_leaf_322_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][20] ),
    .QN(_09554_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][21]$_DFFE_PP_  (.D(_00700_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][21] ),
    .QN(_09553_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][22]$_DFFE_PP_  (.D(_00701_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][22] ),
    .QN(_09552_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][23]$_DFFE_PP_  (.D(_00702_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][23] ),
    .QN(_09551_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][24]$_DFFE_PP_  (.D(_00703_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][24] ),
    .QN(_09550_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][25]$_DFFE_PP_  (.D(_00704_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][25] ),
    .QN(_09549_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][26]$_DFFE_PP_  (.D(_00705_),
    .CK(clknet_leaf_37_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][26] ),
    .QN(_09548_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][27]$_DFFE_PP_  (.D(_00706_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][27] ),
    .QN(_09547_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][28]$_DFFE_PP_  (.D(_00707_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][28] ),
    .QN(_09546_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][29]$_DFFE_PP_  (.D(_00708_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][29] ),
    .QN(_09545_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][2]$_DFFE_PP_  (.D(_00709_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][2] ),
    .QN(_09544_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][30]$_DFFE_PP_  (.D(_00710_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][30] ),
    .QN(_09543_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][31]$_DFFE_PP_  (.D(_00711_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][31] ),
    .QN(_09542_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][32]$_DFFE_PP_  (.D(_00712_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][32] ),
    .QN(_09541_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][33]$_DFFE_PP_  (.D(_00713_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][33] ),
    .QN(_09540_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][34]$_DFFE_PP_  (.D(_00714_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][34] ),
    .QN(_09539_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][35]$_DFFE_PP_  (.D(_00715_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][35] ),
    .QN(_09538_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][36]$_DFFE_PP_  (.D(_00716_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][36] ),
    .QN(_09537_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][37]$_DFFE_PP_  (.D(_00717_),
    .CK(clknet_leaf_103_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][37] ),
    .QN(_09536_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][38]$_DFFE_PP_  (.D(_00718_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][38] ),
    .QN(_09535_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][39]$_DFFE_PP_  (.D(_00719_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][39] ),
    .QN(_09534_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][3]$_DFFE_PP_  (.D(_00720_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][3] ),
    .QN(_09533_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][40]$_DFFE_PP_  (.D(_00721_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][40] ),
    .QN(_09532_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][41]$_DFFE_PP_  (.D(_00722_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][41] ),
    .QN(_09531_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][42]$_DFFE_PP_  (.D(_00723_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][42] ),
    .QN(_09530_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][43]$_DFFE_PP_  (.D(_00724_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][43] ),
    .QN(_09529_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][44]$_DFFE_PP_  (.D(_00725_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][44] ),
    .QN(_09528_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][45]$_DFFE_PP_  (.D(_00726_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][45] ),
    .QN(_09527_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][46]$_DFFE_PP_  (.D(_00727_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][46] ),
    .QN(_09526_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][47]$_DFFE_PP_  (.D(_00728_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][47] ),
    .QN(_09525_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][48]$_DFFE_PP_  (.D(_00729_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][48] ),
    .QN(_09524_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][49]$_DFFE_PP_  (.D(_00730_),
    .CK(clknet_leaf_112_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][49] ),
    .QN(_09523_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][4]$_DFFE_PP_  (.D(_00731_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][4] ),
    .QN(_09522_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][50]$_DFFE_PP_  (.D(_00732_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][50] ),
    .QN(_09521_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][51]$_DFFE_PP_  (.D(_00733_),
    .CK(clknet_leaf_55_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][51] ),
    .QN(_09520_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][52]$_DFFE_PP_  (.D(_00734_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][52] ),
    .QN(_09519_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][53]$_DFFE_PP_  (.D(_00735_),
    .CK(clknet_leaf_111_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][53] ),
    .QN(_09518_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][54]$_DFFE_PP_  (.D(_00736_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][54] ),
    .QN(_09517_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][55]$_DFFE_PP_  (.D(_00737_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][55] ),
    .QN(_09516_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][56]$_DFFE_PP_  (.D(_00738_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][56] ),
    .QN(_09515_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][57]$_DFFE_PP_  (.D(_00739_),
    .CK(clknet_leaf_51_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][57] ),
    .QN(_09514_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][58]$_DFFE_PP_  (.D(_00740_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][58] ),
    .QN(_09513_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][59]$_DFFE_PP_  (.D(_00741_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][59] ),
    .QN(_09512_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][5]$_DFFE_PP_  (.D(_00742_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][5] ),
    .QN(_09511_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][60]$_DFFE_PP_  (.D(_00743_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][60] ),
    .QN(_09510_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][61]$_DFFE_PP_  (.D(_00744_),
    .CK(clknet_leaf_46_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][61] ),
    .QN(_09509_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][62]$_DFFE_PP_  (.D(_00745_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][62] ),
    .QN(_09508_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][63]$_DFFE_PP_  (.D(_00746_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][63] ),
    .QN(_09507_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][6]$_DFFE_PP_  (.D(_00747_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][6] ),
    .QN(_09506_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][7]$_DFFE_PP_  (.D(_00748_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][7] ),
    .QN(_09505_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][8]$_DFFE_PP_  (.D(_00749_),
    .CK(clknet_leaf_17_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][8] ),
    .QN(_09504_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[0][9]$_DFFE_PP_  (.D(_00750_),
    .CK(clknet_leaf_17_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[0][9] ),
    .QN(_09503_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][0]$_DFFE_PP_  (.D(_00751_),
    .CK(clknet_leaf_30_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][0] ),
    .QN(_09502_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][10]$_DFFE_PP_  (.D(_00752_),
    .CK(clknet_leaf_6_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][10] ),
    .QN(_09501_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][11]$_DFFE_PP_  (.D(_00753_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][11] ),
    .QN(_09500_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][12]$_DFFE_PP_  (.D(_00754_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][12] ),
    .QN(_09499_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][13]$_DFFE_PP_  (.D(_00755_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][13] ),
    .QN(_09498_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][14]$_DFFE_PP_  (.D(_00756_),
    .CK(clknet_leaf_6_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][14] ),
    .QN(_09497_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][15]$_DFFE_PP_  (.D(_00757_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][15] ),
    .QN(_09496_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][16]$_DFFE_PP_  (.D(_00758_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][16] ),
    .QN(_09495_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][17]$_DFFE_PP_  (.D(_00759_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][17] ),
    .QN(_09494_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][18]$_DFFE_PP_  (.D(_00760_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][18] ),
    .QN(_09493_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][19]$_DFFE_PP_  (.D(_00761_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][19] ),
    .QN(_09492_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][1]$_DFFE_PP_  (.D(_00762_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][1] ),
    .QN(_09491_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][20]$_DFFE_PP_  (.D(_00763_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][20] ),
    .QN(_09490_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][21]$_DFFE_PP_  (.D(_00764_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][21] ),
    .QN(_09489_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][22]$_DFFE_PP_  (.D(_00765_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][22] ),
    .QN(_09488_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][23]$_DFFE_PP_  (.D(_00766_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][23] ),
    .QN(_09487_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][24]$_DFFE_PP_  (.D(_00767_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][24] ),
    .QN(_09486_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][25]$_DFFE_PP_  (.D(_00768_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][25] ),
    .QN(_09485_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][26]$_DFFE_PP_  (.D(_00769_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][26] ),
    .QN(_09484_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][27]$_DFFE_PP_  (.D(_00770_),
    .CK(clknet_leaf_320_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][27] ),
    .QN(_09483_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][28]$_DFFE_PP_  (.D(_00771_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][28] ),
    .QN(_09482_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][29]$_DFFE_PP_  (.D(_00772_),
    .CK(clknet_leaf_56_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][29] ),
    .QN(_09481_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][2]$_DFFE_PP_  (.D(_00773_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][2] ),
    .QN(_09480_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][30]$_DFFE_PP_  (.D(_00774_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][30] ),
    .QN(_09479_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][31]$_DFFE_PP_  (.D(_00775_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][31] ),
    .QN(_09478_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][32]$_DFFE_PP_  (.D(_00776_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][32] ),
    .QN(_09477_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][33]$_DFFE_PP_  (.D(_00777_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][33] ),
    .QN(_09476_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][34]$_DFFE_PP_  (.D(_00778_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][34] ),
    .QN(_09475_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][35]$_DFFE_PP_  (.D(_00779_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][35] ),
    .QN(_09474_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][36]$_DFFE_PP_  (.D(_00780_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][36] ),
    .QN(_09473_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][37]$_DFFE_PP_  (.D(_00781_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][37] ),
    .QN(_09472_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][38]$_DFFE_PP_  (.D(_00782_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][38] ),
    .QN(_09471_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][39]$_DFFE_PP_  (.D(_00783_),
    .CK(clknet_leaf_86_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][39] ),
    .QN(_09470_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][3]$_DFFE_PP_  (.D(_00784_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][3] ),
    .QN(_09469_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][40]$_DFFE_PP_  (.D(_00785_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][40] ),
    .QN(_09468_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][41]$_DFFE_PP_  (.D(_00786_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][41] ),
    .QN(_09467_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][42]$_DFFE_PP_  (.D(_00787_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][42] ),
    .QN(_09466_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][43]$_DFFE_PP_  (.D(_00788_),
    .CK(clknet_leaf_98_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][43] ),
    .QN(_09465_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][44]$_DFFE_PP_  (.D(_00789_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][44] ),
    .QN(_09464_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][45]$_DFFE_PP_  (.D(_00790_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][45] ),
    .QN(_09463_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][46]$_DFFE_PP_  (.D(_00791_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][46] ),
    .QN(_09462_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][47]$_DFFE_PP_  (.D(_00792_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][47] ),
    .QN(_09461_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][48]$_DFFE_PP_  (.D(_00793_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][48] ),
    .QN(_09460_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][49]$_DFFE_PP_  (.D(_00794_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][49] ),
    .QN(_09459_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][4]$_DFFE_PP_  (.D(_00795_),
    .CK(clknet_leaf_56_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][4] ),
    .QN(_09458_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][50]$_DFFE_PP_  (.D(_00796_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][50] ),
    .QN(_09457_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][51]$_DFFE_PP_  (.D(_00797_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][51] ),
    .QN(_09456_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][52]$_DFFE_PP_  (.D(_00798_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][52] ),
    .QN(_09455_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][53]$_DFFE_PP_  (.D(_00799_),
    .CK(clknet_leaf_111_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][53] ),
    .QN(_09454_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][54]$_DFFE_PP_  (.D(_00800_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][54] ),
    .QN(_09453_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][55]$_DFFE_PP_  (.D(_00801_),
    .CK(clknet_leaf_51_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][55] ),
    .QN(_09452_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][56]$_DFFE_PP_  (.D(_00802_),
    .CK(clknet_leaf_296_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][56] ),
    .QN(_09451_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][57]$_DFFE_PP_  (.D(_00803_),
    .CK(clknet_leaf_51_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][57] ),
    .QN(_09450_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][58]$_DFFE_PP_  (.D(_00804_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][58] ),
    .QN(_09449_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][59]$_DFFE_PP_  (.D(_00805_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][59] ),
    .QN(_09448_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][5]$_DFFE_PP_  (.D(_00806_),
    .CK(clknet_leaf_40_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][5] ),
    .QN(_09447_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][60]$_DFFE_PP_  (.D(_00807_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][60] ),
    .QN(_09446_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][61]$_DFFE_PP_  (.D(_00808_),
    .CK(clknet_leaf_45_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][61] ),
    .QN(_09445_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][62]$_DFFE_PP_  (.D(_00809_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][62] ),
    .QN(_09444_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][63]$_DFFE_PP_  (.D(_00810_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][63] ),
    .QN(_09443_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][6]$_DFFE_PP_  (.D(_00811_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][6] ),
    .QN(_09442_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][7]$_DFFE_PP_  (.D(_00812_),
    .CK(clknet_leaf_25_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][7] ),
    .QN(_09441_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][8]$_DFFE_PP_  (.D(_00813_),
    .CK(clknet_leaf_30_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][8] ),
    .QN(_09440_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[10][9]$_DFFE_PP_  (.D(_00814_),
    .CK(clknet_leaf_23_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[10][9] ),
    .QN(_09439_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][0]$_DFFE_PP_  (.D(_00815_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][0] ),
    .QN(_09438_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][10]$_DFFE_PP_  (.D(_00816_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][10] ),
    .QN(_09437_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][11]$_DFFE_PP_  (.D(_00817_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][11] ),
    .QN(_09436_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][12]$_DFFE_PP_  (.D(_00818_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][12] ),
    .QN(_09435_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][13]$_DFFE_PP_  (.D(_00819_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][13] ),
    .QN(_09434_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][14]$_DFFE_PP_  (.D(_00820_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][14] ),
    .QN(_09433_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][15]$_DFFE_PP_  (.D(_00821_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][15] ),
    .QN(_09432_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][16]$_DFFE_PP_  (.D(_00822_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][16] ),
    .QN(_09431_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][17]$_DFFE_PP_  (.D(_00823_),
    .CK(clknet_leaf_6_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][17] ),
    .QN(_09430_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][18]$_DFFE_PP_  (.D(_00824_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][18] ),
    .QN(_09429_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][19]$_DFFE_PP_  (.D(_00825_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][19] ),
    .QN(_09428_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][1]$_DFFE_PP_  (.D(_00826_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][1] ),
    .QN(_09427_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][20]$_DFFE_PP_  (.D(_00827_),
    .CK(clknet_leaf_322_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][20] ),
    .QN(_09426_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][21]$_DFFE_PP_  (.D(_00828_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][21] ),
    .QN(_09425_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][22]$_DFFE_PP_  (.D(_00829_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][22] ),
    .QN(_09424_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][23]$_DFFE_PP_  (.D(_00830_),
    .CK(clknet_leaf_320_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][23] ),
    .QN(_09423_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][24]$_DFFE_PP_  (.D(_00831_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][24] ),
    .QN(_09422_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][25]$_DFFE_PP_  (.D(_00832_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][25] ),
    .QN(_09421_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][26]$_DFFE_PP_  (.D(_00833_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][26] ),
    .QN(_09420_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][27]$_DFFE_PP_  (.D(_00834_),
    .CK(clknet_leaf_320_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][27] ),
    .QN(_09419_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][28]$_DFFE_PP_  (.D(_00835_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][28] ),
    .QN(_09418_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][29]$_DFFE_PP_  (.D(_00836_),
    .CK(clknet_leaf_55_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][29] ),
    .QN(_09417_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][2]$_DFFE_PP_  (.D(_00837_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][2] ),
    .QN(_09416_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][30]$_DFFE_PP_  (.D(_00838_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][30] ),
    .QN(_09415_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][31]$_DFFE_PP_  (.D(_00839_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][31] ),
    .QN(_09414_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][32]$_DFFE_PP_  (.D(_00840_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][32] ),
    .QN(_09413_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][33]$_DFFE_PP_  (.D(_00841_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][33] ),
    .QN(_09412_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][34]$_DFFE_PP_  (.D(_00842_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][34] ),
    .QN(_09411_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][35]$_DFFE_PP_  (.D(_00843_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][35] ),
    .QN(_09410_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][36]$_DFFE_PP_  (.D(_00844_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][36] ),
    .QN(_09409_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][37]$_DFFE_PP_  (.D(_00845_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][37] ),
    .QN(_09408_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][38]$_DFFE_PP_  (.D(_00846_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][38] ),
    .QN(_09407_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][39]$_DFFE_PP_  (.D(_00847_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][39] ),
    .QN(_09406_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][3]$_DFFE_PP_  (.D(_00848_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][3] ),
    .QN(_09405_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][40]$_DFFE_PP_  (.D(_00849_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][40] ),
    .QN(_09404_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][41]$_DFFE_PP_  (.D(_00850_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][41] ),
    .QN(_09403_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][42]$_DFFE_PP_  (.D(_00851_),
    .CK(clknet_leaf_82_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][42] ),
    .QN(_09402_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][43]$_DFFE_PP_  (.D(_00852_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][43] ),
    .QN(_09401_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][44]$_DFFE_PP_  (.D(_00853_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][44] ),
    .QN(_09400_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][45]$_DFFE_PP_  (.D(_00854_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][45] ),
    .QN(_09399_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][46]$_DFFE_PP_  (.D(_00855_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][46] ),
    .QN(_09398_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][47]$_DFFE_PP_  (.D(_00856_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][47] ),
    .QN(_09397_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][48]$_DFFE_PP_  (.D(_00857_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][48] ),
    .QN(_09396_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][49]$_DFFE_PP_  (.D(_00858_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][49] ),
    .QN(_09395_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][4]$_DFFE_PP_  (.D(_00859_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][4] ),
    .QN(_09394_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][50]$_DFFE_PP_  (.D(_00860_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][50] ),
    .QN(_09393_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][51]$_DFFE_PP_  (.D(_00861_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][51] ),
    .QN(_09392_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][52]$_DFFE_PP_  (.D(_00862_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][52] ),
    .QN(_09391_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][53]$_DFFE_PP_  (.D(_00863_),
    .CK(clknet_leaf_121_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][53] ),
    .QN(_09390_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][54]$_DFFE_PP_  (.D(_00864_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][54] ),
    .QN(_09389_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][55]$_DFFE_PP_  (.D(_00865_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][55] ),
    .QN(_09388_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][56]$_DFFE_PP_  (.D(_00866_),
    .CK(clknet_leaf_304_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][56] ),
    .QN(_09387_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][57]$_DFFE_PP_  (.D(_00867_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][57] ),
    .QN(_09386_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][58]$_DFFE_PP_  (.D(_00868_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][58] ),
    .QN(_09385_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][59]$_DFFE_PP_  (.D(_00869_),
    .CK(clknet_leaf_51_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][59] ),
    .QN(_09384_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][5]$_DFFE_PP_  (.D(_00870_),
    .CK(clknet_leaf_40_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][5] ),
    .QN(_09383_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][60]$_DFFE_PP_  (.D(_00871_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][60] ),
    .QN(_09382_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][61]$_DFFE_PP_  (.D(_00872_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][61] ),
    .QN(_09381_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][62]$_DFFE_PP_  (.D(_00873_),
    .CK(clknet_leaf_302_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][62] ),
    .QN(_09380_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][63]$_DFFE_PP_  (.D(_00874_),
    .CK(clknet_leaf_305_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][63] ),
    .QN(_09379_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][6]$_DFFE_PP_  (.D(_00875_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][6] ),
    .QN(_09378_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][7]$_DFFE_PP_  (.D(_00876_),
    .CK(clknet_leaf_25_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][7] ),
    .QN(_09377_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][8]$_DFFE_PP_  (.D(_00877_),
    .CK(clknet_leaf_23_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][8] ),
    .QN(_09376_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[11][9]$_DFFE_PP_  (.D(_00878_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[11][9] ),
    .QN(_09375_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][0]$_DFFE_PP_  (.D(_00879_),
    .CK(clknet_leaf_30_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][0] ),
    .QN(_09374_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][10]$_DFFE_PP_  (.D(_00880_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][10] ),
    .QN(_09373_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][11]$_DFFE_PP_  (.D(_00881_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][11] ),
    .QN(_09372_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][12]$_DFFE_PP_  (.D(_00882_),
    .CK(clknet_leaf_31_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][12] ),
    .QN(_09371_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][13]$_DFFE_PP_  (.D(_00883_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][13] ),
    .QN(_09370_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][14]$_DFFE_PP_  (.D(_00884_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][14] ),
    .QN(_09369_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][15]$_DFFE_PP_  (.D(_00885_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][15] ),
    .QN(_09368_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][16]$_DFFE_PP_  (.D(_00886_),
    .CK(clknet_leaf_3_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][16] ),
    .QN(_09367_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][17]$_DFFE_PP_  (.D(_00887_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][17] ),
    .QN(_09366_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][18]$_DFFE_PP_  (.D(_00888_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][18] ),
    .QN(_09365_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][19]$_DFFE_PP_  (.D(_00889_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][19] ),
    .QN(_09364_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][1]$_DFFE_PP_  (.D(_00890_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][1] ),
    .QN(_09363_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][20]$_DFFE_PP_  (.D(_00891_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][20] ),
    .QN(_09362_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][21]$_DFFE_PP_  (.D(_00892_),
    .CK(clknet_leaf_36_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][21] ),
    .QN(_09361_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][22]$_DFFE_PP_  (.D(_00893_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][22] ),
    .QN(_09360_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][23]$_DFFE_PP_  (.D(_00894_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][23] ),
    .QN(_09359_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][24]$_DFFE_PP_  (.D(_00895_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][24] ),
    .QN(_09358_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][25]$_DFFE_PP_  (.D(_00896_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][25] ),
    .QN(_09357_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][26]$_DFFE_PP_  (.D(_00897_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][26] ),
    .QN(_09356_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][27]$_DFFE_PP_  (.D(_00898_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][27] ),
    .QN(_09355_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][28]$_DFFE_PP_  (.D(_00899_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][28] ),
    .QN(_09354_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][29]$_DFFE_PP_  (.D(_00900_),
    .CK(clknet_leaf_56_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][29] ),
    .QN(_09353_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][2]$_DFFE_PP_  (.D(_00901_),
    .CK(clknet_leaf_25_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][2] ),
    .QN(_09352_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][30]$_DFFE_PP_  (.D(_00902_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][30] ),
    .QN(_09351_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][31]$_DFFE_PP_  (.D(_00903_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][31] ),
    .QN(_09350_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][32]$_DFFE_PP_  (.D(_00904_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][32] ),
    .QN(_09349_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][33]$_DFFE_PP_  (.D(_00905_),
    .CK(clknet_leaf_72_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][33] ),
    .QN(_09348_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][34]$_DFFE_PP_  (.D(_00906_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][34] ),
    .QN(_09347_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][35]$_DFFE_PP_  (.D(_00907_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][35] ),
    .QN(_09346_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][36]$_DFFE_PP_  (.D(_00908_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][36] ),
    .QN(_09345_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][37]$_DFFE_PP_  (.D(_00909_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][37] ),
    .QN(_09344_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][38]$_DFFE_PP_  (.D(_00910_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][38] ),
    .QN(_09343_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][39]$_DFFE_PP_  (.D(_00911_),
    .CK(clknet_leaf_86_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][39] ),
    .QN(_09342_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][3]$_DFFE_PP_  (.D(_00912_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][3] ),
    .QN(_09341_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][40]$_DFFE_PP_  (.D(_00913_),
    .CK(clknet_leaf_98_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][40] ),
    .QN(_09340_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][41]$_DFFE_PP_  (.D(_00914_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][41] ),
    .QN(_09339_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][42]$_DFFE_PP_  (.D(_00915_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][42] ),
    .QN(_09338_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][43]$_DFFE_PP_  (.D(_00916_),
    .CK(clknet_leaf_98_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][43] ),
    .QN(_09337_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][44]$_DFFE_PP_  (.D(_00917_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][44] ),
    .QN(_09336_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][45]$_DFFE_PP_  (.D(_00918_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][45] ),
    .QN(_09335_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][46]$_DFFE_PP_  (.D(_00919_),
    .CK(clknet_leaf_116_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][46] ),
    .QN(_09334_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][47]$_DFFE_PP_  (.D(_00920_),
    .CK(clknet_leaf_114_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][47] ),
    .QN(_09333_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][48]$_DFFE_PP_  (.D(_00921_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][48] ),
    .QN(_09332_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][49]$_DFFE_PP_  (.D(_00922_),
    .CK(clknet_leaf_111_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][49] ),
    .QN(_09331_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][4]$_DFFE_PP_  (.D(_00923_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][4] ),
    .QN(_09330_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][50]$_DFFE_PP_  (.D(_00924_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][50] ),
    .QN(_09329_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][51]$_DFFE_PP_  (.D(_00925_),
    .CK(clknet_leaf_60_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][51] ),
    .QN(_09328_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][52]$_DFFE_PP_  (.D(_00926_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][52] ),
    .QN(_09327_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][53]$_DFFE_PP_  (.D(_00927_),
    .CK(clknet_leaf_121_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][53] ),
    .QN(_09326_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][54]$_DFFE_PP_  (.D(_00928_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][54] ),
    .QN(_09325_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][55]$_DFFE_PP_  (.D(_00929_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][55] ),
    .QN(_09324_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][56]$_DFFE_PP_  (.D(_00930_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][56] ),
    .QN(_09323_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][57]$_DFFE_PP_  (.D(_00931_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][57] ),
    .QN(_09322_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][58]$_DFFE_PP_  (.D(_00932_),
    .CK(clknet_leaf_302_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][58] ),
    .QN(_09321_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][59]$_DFFE_PP_  (.D(_00933_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][59] ),
    .QN(_09320_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][5]$_DFFE_PP_  (.D(_00934_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][5] ),
    .QN(_09319_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][60]$_DFFE_PP_  (.D(_00935_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][60] ),
    .QN(_09318_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][61]$_DFFE_PP_  (.D(_00936_),
    .CK(clknet_leaf_45_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][61] ),
    .QN(_09317_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][62]$_DFFE_PP_  (.D(_00937_),
    .CK(clknet_leaf_301_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][62] ),
    .QN(_09316_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][63]$_DFFE_PP_  (.D(_00938_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][63] ),
    .QN(_09315_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][6]$_DFFE_PP_  (.D(_00939_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][6] ),
    .QN(_09314_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][7]$_DFFE_PP_  (.D(_00940_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][7] ),
    .QN(_09313_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][8]$_DFFE_PP_  (.D(_00941_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][8] ),
    .QN(_09312_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[12][9]$_DFFE_PP_  (.D(_00942_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[12][9] ),
    .QN(_09311_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][0]$_DFFE_PP_  (.D(_00943_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][0] ),
    .QN(_09310_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][10]$_DFFE_PP_  (.D(_00944_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][10] ),
    .QN(_09309_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][11]$_DFFE_PP_  (.D(_00945_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][11] ),
    .QN(_09308_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][12]$_DFFE_PP_  (.D(_00946_),
    .CK(clknet_leaf_31_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][12] ),
    .QN(_09307_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][13]$_DFFE_PP_  (.D(_00947_),
    .CK(clknet_leaf_3_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][13] ),
    .QN(_09306_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][14]$_DFFE_PP_  (.D(_00948_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][14] ),
    .QN(_09305_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][15]$_DFFE_PP_  (.D(_00949_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][15] ),
    .QN(_09304_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][16]$_DFFE_PP_  (.D(_00950_),
    .CK(clknet_leaf_3_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][16] ),
    .QN(_09303_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][17]$_DFFE_PP_  (.D(_00951_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][17] ),
    .QN(_09302_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][18]$_DFFE_PP_  (.D(_00952_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][18] ),
    .QN(_09301_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][19]$_DFFE_PP_  (.D(_00953_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][19] ),
    .QN(_09300_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][1]$_DFFE_PP_  (.D(_00954_),
    .CK(clknet_leaf_37_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][1] ),
    .QN(_09299_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][20]$_DFFE_PP_  (.D(_00955_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][20] ),
    .QN(_09298_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][21]$_DFFE_PP_  (.D(_00956_),
    .CK(clknet_leaf_36_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][21] ),
    .QN(_09297_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][22]$_DFFE_PP_  (.D(_00957_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][22] ),
    .QN(_09296_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][23]$_DFFE_PP_  (.D(_00958_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][23] ),
    .QN(_09295_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][24]$_DFFE_PP_  (.D(_00959_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][24] ),
    .QN(_09294_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][25]$_DFFE_PP_  (.D(_00960_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][25] ),
    .QN(_09293_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][26]$_DFFE_PP_  (.D(_00961_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][26] ),
    .QN(_09292_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][27]$_DFFE_PP_  (.D(_00962_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][27] ),
    .QN(_09291_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][28]$_DFFE_PP_  (.D(_00963_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][28] ),
    .QN(_09290_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][29]$_DFFE_PP_  (.D(_00964_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][29] ),
    .QN(_09289_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][2]$_DFFE_PP_  (.D(_00965_),
    .CK(clknet_leaf_25_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][2] ),
    .QN(_09288_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][30]$_DFFE_PP_  (.D(_00966_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][30] ),
    .QN(_09287_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][31]$_DFFE_PP_  (.D(_00967_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][31] ),
    .QN(_09286_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][32]$_DFFE_PP_  (.D(_00968_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][32] ),
    .QN(_09285_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][33]$_DFFE_PP_  (.D(_00969_),
    .CK(clknet_leaf_72_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][33] ),
    .QN(_09284_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][34]$_DFFE_PP_  (.D(_00970_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][34] ),
    .QN(_09283_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][35]$_DFFE_PP_  (.D(_00971_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][35] ),
    .QN(_09282_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][36]$_DFFE_PP_  (.D(_00972_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][36] ),
    .QN(_09281_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][37]$_DFFE_PP_  (.D(_00973_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][37] ),
    .QN(_09280_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][38]$_DFFE_PP_  (.D(_00974_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][38] ),
    .QN(_09279_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][39]$_DFFE_PP_  (.D(_00975_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][39] ),
    .QN(_09278_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][3]$_DFFE_PP_  (.D(_00976_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][3] ),
    .QN(_09277_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][40]$_DFFE_PP_  (.D(_00977_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][40] ),
    .QN(_09276_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][41]$_DFFE_PP_  (.D(_00978_),
    .CK(clknet_leaf_92_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][41] ),
    .QN(_09275_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][42]$_DFFE_PP_  (.D(_00979_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][42] ),
    .QN(_09274_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][43]$_DFFE_PP_  (.D(_00980_),
    .CK(clknet_leaf_98_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][43] ),
    .QN(_09273_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][44]$_DFFE_PP_  (.D(_00981_),
    .CK(clknet_leaf_86_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][44] ),
    .QN(_09272_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][45]$_DFFE_PP_  (.D(_00982_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][45] ),
    .QN(_09271_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][46]$_DFFE_PP_  (.D(_00983_),
    .CK(clknet_leaf_116_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][46] ),
    .QN(_09270_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][47]$_DFFE_PP_  (.D(_00984_),
    .CK(clknet_leaf_114_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][47] ),
    .QN(_09269_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][48]$_DFFE_PP_  (.D(_00985_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][48] ),
    .QN(_09268_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][49]$_DFFE_PP_  (.D(_00986_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][49] ),
    .QN(_09267_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][4]$_DFFE_PP_  (.D(_00987_),
    .CK(clknet_leaf_56_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][4] ),
    .QN(_09266_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][50]$_DFFE_PP_  (.D(_00988_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][50] ),
    .QN(_09265_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][51]$_DFFE_PP_  (.D(_00989_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][51] ),
    .QN(_09264_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][52]$_DFFE_PP_  (.D(_00990_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][52] ),
    .QN(_09263_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][53]$_DFFE_PP_  (.D(_00991_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][53] ),
    .QN(_09262_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][54]$_DFFE_PP_  (.D(_00992_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][54] ),
    .QN(_09261_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][55]$_DFFE_PP_  (.D(_00993_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][55] ),
    .QN(_09260_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][56]$_DFFE_PP_  (.D(_00994_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][56] ),
    .QN(_09259_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][57]$_DFFE_PP_  (.D(_00995_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][57] ),
    .QN(_09258_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][58]$_DFFE_PP_  (.D(_00996_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][58] ),
    .QN(_09257_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][59]$_DFFE_PP_  (.D(_00997_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][59] ),
    .QN(_09256_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][5]$_DFFE_PP_  (.D(_00998_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][5] ),
    .QN(_09255_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][60]$_DFFE_PP_  (.D(_00999_),
    .CK(clknet_leaf_304_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][60] ),
    .QN(_09254_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][61]$_DFFE_PP_  (.D(_01000_),
    .CK(clknet_leaf_45_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][61] ),
    .QN(_09253_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][62]$_DFFE_PP_  (.D(_01001_),
    .CK(clknet_leaf_301_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][62] ),
    .QN(_09252_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][63]$_DFFE_PP_  (.D(_01002_),
    .CK(clknet_leaf_305_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][63] ),
    .QN(_09251_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][6]$_DFFE_PP_  (.D(_01003_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][6] ),
    .QN(_09250_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][7]$_DFFE_PP_  (.D(_01004_),
    .CK(clknet_leaf_25_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][7] ),
    .QN(_09249_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][8]$_DFFE_PP_  (.D(_01005_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][8] ),
    .QN(_09248_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[13][9]$_DFFE_PP_  (.D(_01006_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[13][9] ),
    .QN(_09247_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][0]$_DFFE_PP_  (.D(_01007_),
    .CK(clknet_leaf_30_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][0] ),
    .QN(_09246_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][10]$_DFFE_PP_  (.D(_01008_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][10] ),
    .QN(_09245_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][11]$_DFFE_PP_  (.D(_01009_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][11] ),
    .QN(_09244_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][12]$_DFFE_PP_  (.D(_01010_),
    .CK(clknet_leaf_31_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][12] ),
    .QN(_09243_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][13]$_DFFE_PP_  (.D(_01011_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][13] ),
    .QN(_09242_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][14]$_DFFE_PP_  (.D(_01012_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][14] ),
    .QN(_09241_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][15]$_DFFE_PP_  (.D(_01013_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][15] ),
    .QN(_09240_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][16]$_DFFE_PP_  (.D(_01014_),
    .CK(clknet_leaf_3_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][16] ),
    .QN(_09239_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][17]$_DFFE_PP_  (.D(_01015_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][17] ),
    .QN(_09238_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][18]$_DFFE_PP_  (.D(_01016_),
    .CK(clknet_leaf_31_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][18] ),
    .QN(_09237_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][19]$_DFFE_PP_  (.D(_01017_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][19] ),
    .QN(_09236_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][1]$_DFFE_PP_  (.D(_01018_),
    .CK(clknet_leaf_36_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][1] ),
    .QN(_09235_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][20]$_DFFE_PP_  (.D(_01019_),
    .CK(clknet_leaf_322_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][20] ),
    .QN(_09234_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][21]$_DFFE_PP_  (.D(_01020_),
    .CK(clknet_leaf_36_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][21] ),
    .QN(_09233_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][22]$_DFFE_PP_  (.D(_01021_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][22] ),
    .QN(_09232_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][23]$_DFFE_PP_  (.D(_01022_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][23] ),
    .QN(_09231_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][24]$_DFFE_PP_  (.D(_01023_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][24] ),
    .QN(_09230_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][25]$_DFFE_PP_  (.D(_01024_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][25] ),
    .QN(_09229_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][26]$_DFFE_PP_  (.D(_01025_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][26] ),
    .QN(_09228_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][27]$_DFFE_PP_  (.D(_01026_),
    .CK(clknet_leaf_320_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][27] ),
    .QN(_09227_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][28]$_DFFE_PP_  (.D(_01027_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][28] ),
    .QN(_09226_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][29]$_DFFE_PP_  (.D(_01028_),
    .CK(clknet_leaf_55_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][29] ),
    .QN(_09225_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][2]$_DFFE_PP_  (.D(_01029_),
    .CK(clknet_leaf_25_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][2] ),
    .QN(_09224_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][30]$_DFFE_PP_  (.D(_01030_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][30] ),
    .QN(_09223_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][31]$_DFFE_PP_  (.D(_01031_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][31] ),
    .QN(_09222_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][32]$_DFFE_PP_  (.D(_01032_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][32] ),
    .QN(_09221_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][33]$_DFFE_PP_  (.D(_01033_),
    .CK(clknet_leaf_72_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][33] ),
    .QN(_09220_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][34]$_DFFE_PP_  (.D(_01034_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][34] ),
    .QN(_09219_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][35]$_DFFE_PP_  (.D(_01035_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][35] ),
    .QN(_09218_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][36]$_DFFE_PP_  (.D(_01036_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][36] ),
    .QN(_09217_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][37]$_DFFE_PP_  (.D(_01037_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][37] ),
    .QN(_09216_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][38]$_DFFE_PP_  (.D(_01038_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][38] ),
    .QN(_09215_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][39]$_DFFE_PP_  (.D(_01039_),
    .CK(clknet_leaf_86_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][39] ),
    .QN(_09214_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][3]$_DFFE_PP_  (.D(_01040_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][3] ),
    .QN(_09213_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][40]$_DFFE_PP_  (.D(_01041_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][40] ),
    .QN(_09212_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][41]$_DFFE_PP_  (.D(_01042_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][41] ),
    .QN(_09211_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][42]$_DFFE_PP_  (.D(_01043_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][42] ),
    .QN(_09210_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][43]$_DFFE_PP_  (.D(_01044_),
    .CK(clknet_leaf_98_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][43] ),
    .QN(_09209_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][44]$_DFFE_PP_  (.D(_01045_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][44] ),
    .QN(_09208_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][45]$_DFFE_PP_  (.D(_01046_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][45] ),
    .QN(_09207_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][46]$_DFFE_PP_  (.D(_01047_),
    .CK(clknet_leaf_116_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][46] ),
    .QN(_09206_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][47]$_DFFE_PP_  (.D(_01048_),
    .CK(clknet_leaf_114_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][47] ),
    .QN(_09205_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][48]$_DFFE_PP_  (.D(_01049_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][48] ),
    .QN(_09204_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][49]$_DFFE_PP_  (.D(_01050_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][49] ),
    .QN(_09203_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][4]$_DFFE_PP_  (.D(_01051_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][4] ),
    .QN(_09202_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][50]$_DFFE_PP_  (.D(_01052_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][50] ),
    .QN(_09201_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][51]$_DFFE_PP_  (.D(_01053_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][51] ),
    .QN(_09200_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][52]$_DFFE_PP_  (.D(_01054_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][52] ),
    .QN(_09199_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][53]$_DFFE_PP_  (.D(_01055_),
    .CK(clknet_leaf_121_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][53] ),
    .QN(_09198_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][54]$_DFFE_PP_  (.D(_01056_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][54] ),
    .QN(_09197_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][55]$_DFFE_PP_  (.D(_01057_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][55] ),
    .QN(_09196_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][56]$_DFFE_PP_  (.D(_01058_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][56] ),
    .QN(_09195_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][57]$_DFFE_PP_  (.D(_01059_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][57] ),
    .QN(_09194_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][58]$_DFFE_PP_  (.D(_01060_),
    .CK(clknet_leaf_50_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][58] ),
    .QN(_09193_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][59]$_DFFE_PP_  (.D(_01061_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][59] ),
    .QN(_09192_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][5]$_DFFE_PP_  (.D(_01062_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][5] ),
    .QN(_09191_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][60]$_DFFE_PP_  (.D(_01063_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][60] ),
    .QN(_09190_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][61]$_DFFE_PP_  (.D(_01064_),
    .CK(clknet_leaf_45_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][61] ),
    .QN(_09189_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][62]$_DFFE_PP_  (.D(_01065_),
    .CK(clknet_leaf_302_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][62] ),
    .QN(_09188_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][63]$_DFFE_PP_  (.D(_01066_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][63] ),
    .QN(_09187_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][6]$_DFFE_PP_  (.D(_01067_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][6] ),
    .QN(_09186_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][7]$_DFFE_PP_  (.D(_01068_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][7] ),
    .QN(_09185_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][8]$_DFFE_PP_  (.D(_01069_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][8] ),
    .QN(_09184_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[14][9]$_DFFE_PP_  (.D(_01070_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[14][9] ),
    .QN(_09183_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][0]$_DFFE_PP_  (.D(_01071_),
    .CK(clknet_leaf_30_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][0] ),
    .QN(_09182_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][10]$_DFFE_PP_  (.D(_01072_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][10] ),
    .QN(_09181_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][11]$_DFFE_PP_  (.D(_01073_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][11] ),
    .QN(_09180_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][12]$_DFFE_PP_  (.D(_01074_),
    .CK(clknet_leaf_31_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][12] ),
    .QN(_09179_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][13]$_DFFE_PP_  (.D(_01075_),
    .CK(clknet_leaf_3_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][13] ),
    .QN(_09178_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][14]$_DFFE_PP_  (.D(_01076_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][14] ),
    .QN(_09177_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][15]$_DFFE_PP_  (.D(_01077_),
    .CK(clknet_leaf_5_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][15] ),
    .QN(_09176_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][16]$_DFFE_PP_  (.D(_01078_),
    .CK(clknet_leaf_3_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][16] ),
    .QN(_09175_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][17]$_DFFE_PP_  (.D(_01079_),
    .CK(clknet_leaf_6_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][17] ),
    .QN(_09174_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][18]$_DFFE_PP_  (.D(_01080_),
    .CK(clknet_leaf_31_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][18] ),
    .QN(_09173_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][19]$_DFFE_PP_  (.D(_01081_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][19] ),
    .QN(_09172_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][1]$_DFFE_PP_  (.D(_01082_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][1] ),
    .QN(_09171_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][20]$_DFFE_PP_  (.D(_01083_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][20] ),
    .QN(_09170_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][21]$_DFFE_PP_  (.D(_01084_),
    .CK(clknet_leaf_40_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][21] ),
    .QN(_09169_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][22]$_DFFE_PP_  (.D(_01085_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][22] ),
    .QN(_09168_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][23]$_DFFE_PP_  (.D(_01086_),
    .CK(clknet_leaf_320_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][23] ),
    .QN(_09167_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][24]$_DFFE_PP_  (.D(_01087_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][24] ),
    .QN(_09166_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][25]$_DFFE_PP_  (.D(_01088_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][25] ),
    .QN(_09165_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][26]$_DFFE_PP_  (.D(_01089_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][26] ),
    .QN(_09164_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][27]$_DFFE_PP_  (.D(_01090_),
    .CK(clknet_leaf_320_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][27] ),
    .QN(_09163_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][28]$_DFFE_PP_  (.D(_01091_),
    .CK(clknet_leaf_55_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][28] ),
    .QN(_09162_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][29]$_DFFE_PP_  (.D(_01092_),
    .CK(clknet_leaf_55_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][29] ),
    .QN(_09161_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][2]$_DFFE_PP_  (.D(_01093_),
    .CK(clknet_leaf_72_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][2] ),
    .QN(_09160_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][30]$_DFFE_PP_  (.D(_01094_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][30] ),
    .QN(_09159_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][31]$_DFFE_PP_  (.D(_01095_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][31] ),
    .QN(_09158_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][32]$_DFFE_PP_  (.D(_01096_),
    .CK(clknet_leaf_60_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][32] ),
    .QN(_09157_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][33]$_DFFE_PP_  (.D(_01097_),
    .CK(clknet_leaf_72_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][33] ),
    .QN(_09156_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][34]$_DFFE_PP_  (.D(_01098_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][34] ),
    .QN(_09155_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][35]$_DFFE_PP_  (.D(_01099_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][35] ),
    .QN(_09154_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][36]$_DFFE_PP_  (.D(_01100_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][36] ),
    .QN(_09153_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][37]$_DFFE_PP_  (.D(_01101_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][37] ),
    .QN(_09152_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][38]$_DFFE_PP_  (.D(_01102_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][38] ),
    .QN(_09151_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][39]$_DFFE_PP_  (.D(_01103_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][39] ),
    .QN(_09150_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][3]$_DFFE_PP_  (.D(_01104_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][3] ),
    .QN(_09149_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][40]$_DFFE_PP_  (.D(_01105_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][40] ),
    .QN(_09148_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][41]$_DFFE_PP_  (.D(_01106_),
    .CK(clknet_leaf_92_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][41] ),
    .QN(_09147_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][42]$_DFFE_PP_  (.D(_01107_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][42] ),
    .QN(_09146_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][43]$_DFFE_PP_  (.D(_01108_),
    .CK(clknet_leaf_98_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][43] ),
    .QN(_09145_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][44]$_DFFE_PP_  (.D(_01109_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][44] ),
    .QN(_09144_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][45]$_DFFE_PP_  (.D(_01110_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][45] ),
    .QN(_09143_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][46]$_DFFE_PP_  (.D(_01111_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][46] ),
    .QN(_09142_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][47]$_DFFE_PP_  (.D(_01112_),
    .CK(clknet_leaf_114_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][47] ),
    .QN(_09141_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][48]$_DFFE_PP_  (.D(_01113_),
    .CK(clknet_leaf_114_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][48] ),
    .QN(_09140_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][49]$_DFFE_PP_  (.D(_01114_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][49] ),
    .QN(_09139_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][4]$_DFFE_PP_  (.D(_01115_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][4] ),
    .QN(_09138_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][50]$_DFFE_PP_  (.D(_01116_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][50] ),
    .QN(_09137_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][51]$_DFFE_PP_  (.D(_01117_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][51] ),
    .QN(_09136_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][52]$_DFFE_PP_  (.D(_01118_),
    .CK(clknet_leaf_126_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][52] ),
    .QN(_09135_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][53]$_DFFE_PP_  (.D(_01119_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][53] ),
    .QN(_09134_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][54]$_DFFE_PP_  (.D(_01120_),
    .CK(clknet_leaf_121_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][54] ),
    .QN(_09133_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][55]$_DFFE_PP_  (.D(_01121_),
    .CK(clknet_leaf_48_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][55] ),
    .QN(_09132_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][56]$_DFFE_PP_  (.D(_01122_),
    .CK(clknet_leaf_304_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][56] ),
    .QN(_09131_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][57]$_DFFE_PP_  (.D(_01123_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][57] ),
    .QN(_09130_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][58]$_DFFE_PP_  (.D(_01124_),
    .CK(clknet_leaf_201_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][58] ),
    .QN(_09129_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][59]$_DFFE_PP_  (.D(_01125_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][59] ),
    .QN(_09128_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][5]$_DFFE_PP_  (.D(_01126_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][5] ),
    .QN(_09127_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][60]$_DFFE_PP_  (.D(_01127_),
    .CK(clknet_leaf_304_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][60] ),
    .QN(_09126_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][61]$_DFFE_PP_  (.D(_01128_),
    .CK(clknet_leaf_45_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][61] ),
    .QN(_09125_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][62]$_DFFE_PP_  (.D(_01129_),
    .CK(clknet_leaf_301_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][62] ),
    .QN(_09124_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][63]$_DFFE_PP_  (.D(_01130_),
    .CK(clknet_leaf_305_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][63] ),
    .QN(_09123_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][6]$_DFFE_PP_  (.D(_01131_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][6] ),
    .QN(_09122_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][7]$_DFFE_PP_  (.D(_01132_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][7] ),
    .QN(_09121_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][8]$_DFFE_PP_  (.D(_01133_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][8] ),
    .QN(_09120_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[15][9]$_DFFE_PP_  (.D(_01134_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[15][9] ),
    .QN(_09119_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][0]$_DFFE_PP_  (.D(_01135_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][0] ),
    .QN(_09118_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][10]$_DFFE_PP_  (.D(_01136_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][10] ),
    .QN(_09117_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][11]$_DFFE_PP_  (.D(_01137_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][11] ),
    .QN(_09116_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][12]$_DFFE_PP_  (.D(_01138_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][12] ),
    .QN(_09115_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][13]$_DFFE_PP_  (.D(_01139_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][13] ),
    .QN(_09114_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][14]$_DFFE_PP_  (.D(_01140_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][14] ),
    .QN(_09113_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][15]$_DFFE_PP_  (.D(_01141_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][15] ),
    .QN(_09112_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][16]$_DFFE_PP_  (.D(_01142_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][16] ),
    .QN(_09111_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][17]$_DFFE_PP_  (.D(_01143_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][17] ),
    .QN(_09110_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][18]$_DFFE_PP_  (.D(_01144_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][18] ),
    .QN(_09109_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][19]$_DFFE_PP_  (.D(_01145_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][19] ),
    .QN(_09108_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][1]$_DFFE_PP_  (.D(_01146_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][1] ),
    .QN(_09107_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][20]$_DFFE_PP_  (.D(_01147_),
    .CK(clknet_leaf_322_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][20] ),
    .QN(_09106_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][21]$_DFFE_PP_  (.D(_01148_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][21] ),
    .QN(_09105_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][22]$_DFFE_PP_  (.D(_01149_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][22] ),
    .QN(_09104_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][23]$_DFFE_PP_  (.D(_01150_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][23] ),
    .QN(_09103_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][24]$_DFFE_PP_  (.D(_01151_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][24] ),
    .QN(_09102_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][25]$_DFFE_PP_  (.D(_01152_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][25] ),
    .QN(_09101_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][26]$_DFFE_PP_  (.D(_01153_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][26] ),
    .QN(_09100_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][27]$_DFFE_PP_  (.D(_01154_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][27] ),
    .QN(_09099_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][28]$_DFFE_PP_  (.D(_01155_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][28] ),
    .QN(_09098_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][29]$_DFFE_PP_  (.D(_01156_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][29] ),
    .QN(_09097_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][2]$_DFFE_PP_  (.D(_01157_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][2] ),
    .QN(_09096_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][30]$_DFFE_PP_  (.D(_01158_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][30] ),
    .QN(_09095_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][31]$_DFFE_PP_  (.D(_01159_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][31] ),
    .QN(_09094_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][32]$_DFFE_PP_  (.D(_01160_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][32] ),
    .QN(_09093_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][33]$_DFFE_PP_  (.D(_01161_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][33] ),
    .QN(_09092_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][34]$_DFFE_PP_  (.D(_01162_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][34] ),
    .QN(_09091_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][35]$_DFFE_PP_  (.D(_01163_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][35] ),
    .QN(_09090_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][36]$_DFFE_PP_  (.D(_01164_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][36] ),
    .QN(_09089_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][37]$_DFFE_PP_  (.D(_01165_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][37] ),
    .QN(_09088_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][38]$_DFFE_PP_  (.D(_01166_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][38] ),
    .QN(_09087_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][39]$_DFFE_PP_  (.D(_01167_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][39] ),
    .QN(_09086_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][3]$_DFFE_PP_  (.D(_01168_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][3] ),
    .QN(_09085_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][40]$_DFFE_PP_  (.D(_01169_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][40] ),
    .QN(_09084_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][41]$_DFFE_PP_  (.D(_01170_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][41] ),
    .QN(_09083_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][42]$_DFFE_PP_  (.D(_01171_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][42] ),
    .QN(_09082_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][43]$_DFFE_PP_  (.D(_01172_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][43] ),
    .QN(_09081_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][44]$_DFFE_PP_  (.D(_01173_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][44] ),
    .QN(_09080_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][45]$_DFFE_PP_  (.D(_01174_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][45] ),
    .QN(_09079_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][46]$_DFFE_PP_  (.D(_01175_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][46] ),
    .QN(_09078_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][47]$_DFFE_PP_  (.D(_01176_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][47] ),
    .QN(_09077_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][48]$_DFFE_PP_  (.D(_01177_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][48] ),
    .QN(_09076_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][49]$_DFFE_PP_  (.D(_01178_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][49] ),
    .QN(_09075_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][4]$_DFFE_PP_  (.D(_01179_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][4] ),
    .QN(_09074_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][50]$_DFFE_PP_  (.D(_01180_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][50] ),
    .QN(_09073_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][51]$_DFFE_PP_  (.D(_01181_),
    .CK(clknet_leaf_60_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][51] ),
    .QN(_09072_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][52]$_DFFE_PP_  (.D(_01182_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][52] ),
    .QN(_09071_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][53]$_DFFE_PP_  (.D(_01183_),
    .CK(clknet_leaf_116_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][53] ),
    .QN(_09070_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][54]$_DFFE_PP_  (.D(_01184_),
    .CK(clknet_leaf_118_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][54] ),
    .QN(_09069_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][55]$_DFFE_PP_  (.D(_01185_),
    .CK(clknet_leaf_48_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][55] ),
    .QN(_09068_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][56]$_DFFE_PP_  (.D(_01186_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][56] ),
    .QN(_09067_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][57]$_DFFE_PP_  (.D(_01187_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][57] ),
    .QN(_09066_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][58]$_DFFE_PP_  (.D(_01188_),
    .CK(clknet_leaf_129_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][58] ),
    .QN(_09065_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][59]$_DFFE_PP_  (.D(_01189_),
    .CK(clknet_leaf_129_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][59] ),
    .QN(_09064_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][5]$_DFFE_PP_  (.D(_01190_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][5] ),
    .QN(_09063_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][60]$_DFFE_PP_  (.D(_01191_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][60] ),
    .QN(_09062_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][61]$_DFFE_PP_  (.D(_01192_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][61] ),
    .QN(_09061_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][62]$_DFFE_PP_  (.D(_01193_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][62] ),
    .QN(_09060_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][63]$_DFFE_PP_  (.D(_01194_),
    .CK(clknet_leaf_305_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][63] ),
    .QN(_09059_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][6]$_DFFE_PP_  (.D(_01195_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][6] ),
    .QN(_09058_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][7]$_DFFE_PP_  (.D(_01196_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][7] ),
    .QN(_09057_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][8]$_DFFE_PP_  (.D(_01197_),
    .CK(clknet_leaf_17_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][8] ),
    .QN(_09056_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[1][9]$_DFFE_PP_  (.D(_01198_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[1][9] ),
    .QN(_09055_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][0]$_DFFE_PP_  (.D(_01199_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][0] ),
    .QN(_09054_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][10]$_DFFE_PP_  (.D(_01200_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][10] ),
    .QN(_09053_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][11]$_DFFE_PP_  (.D(_01201_),
    .CK(clknet_leaf_324_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][11] ),
    .QN(_09052_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][12]$_DFFE_PP_  (.D(_01202_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][12] ),
    .QN(_09051_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][13]$_DFFE_PP_  (.D(_01203_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][13] ),
    .QN(_09050_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][14]$_DFFE_PP_  (.D(_01204_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][14] ),
    .QN(_09049_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][15]$_DFFE_PP_  (.D(_01205_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][15] ),
    .QN(_09048_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][16]$_DFFE_PP_  (.D(_01206_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][16] ),
    .QN(_09047_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][17]$_DFFE_PP_  (.D(_01207_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][17] ),
    .QN(_09046_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][18]$_DFFE_PP_  (.D(_01208_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][18] ),
    .QN(_09045_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][19]$_DFFE_PP_  (.D(_01209_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][19] ),
    .QN(_09044_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][1]$_DFFE_PP_  (.D(_01210_),
    .CK(clknet_leaf_33_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][1] ),
    .QN(_09043_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][20]$_DFFE_PP_  (.D(_01211_),
    .CK(clknet_leaf_322_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][20] ),
    .QN(_09042_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][21]$_DFFE_PP_  (.D(_01212_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][21] ),
    .QN(_09041_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][22]$_DFFE_PP_  (.D(_01213_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][22] ),
    .QN(_09040_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][23]$_DFFE_PP_  (.D(_01214_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][23] ),
    .QN(_09039_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][24]$_DFFE_PP_  (.D(_01215_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][24] ),
    .QN(_09038_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][25]$_DFFE_PP_  (.D(_01216_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][25] ),
    .QN(_09037_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][26]$_DFFE_PP_  (.D(_01217_),
    .CK(clknet_leaf_37_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][26] ),
    .QN(_09036_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][27]$_DFFE_PP_  (.D(_01218_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][27] ),
    .QN(_09035_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][28]$_DFFE_PP_  (.D(_01219_),
    .CK(clknet_leaf_71_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][28] ),
    .QN(_09034_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][29]$_DFFE_PP_  (.D(_01220_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][29] ),
    .QN(_09033_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][2]$_DFFE_PP_  (.D(_01221_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][2] ),
    .QN(_09032_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][30]$_DFFE_PP_  (.D(_01222_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][30] ),
    .QN(_09031_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][31]$_DFFE_PP_  (.D(_01223_),
    .CK(clknet_leaf_67_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][31] ),
    .QN(_09030_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][32]$_DFFE_PP_  (.D(_01224_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][32] ),
    .QN(_09029_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][33]$_DFFE_PP_  (.D(_01225_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][33] ),
    .QN(_09028_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][34]$_DFFE_PP_  (.D(_01226_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][34] ),
    .QN(_09027_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][35]$_DFFE_PP_  (.D(_01227_),
    .CK(clknet_leaf_90_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][35] ),
    .QN(_09026_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][36]$_DFFE_PP_  (.D(_01228_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][36] ),
    .QN(_09025_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][37]$_DFFE_PP_  (.D(_01229_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][37] ),
    .QN(_09024_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][38]$_DFFE_PP_  (.D(_01230_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][38] ),
    .QN(_09023_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][39]$_DFFE_PP_  (.D(_01231_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][39] ),
    .QN(_09022_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][3]$_DFFE_PP_  (.D(_01232_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][3] ),
    .QN(_09021_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][40]$_DFFE_PP_  (.D(_01233_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][40] ),
    .QN(_09020_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][41]$_DFFE_PP_  (.D(_01234_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][41] ),
    .QN(_09019_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][42]$_DFFE_PP_  (.D(_01235_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][42] ),
    .QN(_09018_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][43]$_DFFE_PP_  (.D(_01236_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][43] ),
    .QN(_09017_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][44]$_DFFE_PP_  (.D(_01237_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][44] ),
    .QN(_09016_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][45]$_DFFE_PP_  (.D(_01238_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][45] ),
    .QN(_09015_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][46]$_DFFE_PP_  (.D(_01239_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][46] ),
    .QN(_09014_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][47]$_DFFE_PP_  (.D(_01240_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][47] ),
    .QN(_09013_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][48]$_DFFE_PP_  (.D(_01241_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][48] ),
    .QN(_09012_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][49]$_DFFE_PP_  (.D(_01242_),
    .CK(clknet_leaf_112_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][49] ),
    .QN(_09011_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][4]$_DFFE_PP_  (.D(_01243_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][4] ),
    .QN(_09010_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][50]$_DFFE_PP_  (.D(_01244_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][50] ),
    .QN(_09009_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][51]$_DFFE_PP_  (.D(_01245_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][51] ),
    .QN(_09008_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][52]$_DFFE_PP_  (.D(_01246_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][52] ),
    .QN(_09007_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][53]$_DFFE_PP_  (.D(_01247_),
    .CK(clknet_leaf_121_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][53] ),
    .QN(_09006_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][54]$_DFFE_PP_  (.D(_01248_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][54] ),
    .QN(_09005_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][55]$_DFFE_PP_  (.D(_01249_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][55] ),
    .QN(_09004_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][56]$_DFFE_PP_  (.D(_01250_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][56] ),
    .QN(_09003_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][57]$_DFFE_PP_  (.D(_01251_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][57] ),
    .QN(_09002_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][58]$_DFFE_PP_  (.D(_01252_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][58] ),
    .QN(_09001_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][59]$_DFFE_PP_  (.D(_01253_),
    .CK(clknet_leaf_50_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][59] ),
    .QN(_09000_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][5]$_DFFE_PP_  (.D(_01254_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][5] ),
    .QN(_08999_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][60]$_DFFE_PP_  (.D(_01255_),
    .CK(clknet_leaf_302_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][60] ),
    .QN(_08998_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][61]$_DFFE_PP_  (.D(_01256_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][61] ),
    .QN(_08997_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][62]$_DFFE_PP_  (.D(_01257_),
    .CK(clknet_leaf_302_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][62] ),
    .QN(_08996_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][63]$_DFFE_PP_  (.D(_01258_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][63] ),
    .QN(_08995_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][6]$_DFFE_PP_  (.D(_01259_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][6] ),
    .QN(_08994_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][7]$_DFFE_PP_  (.D(_01260_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][7] ),
    .QN(_08993_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][8]$_DFFE_PP_  (.D(_01261_),
    .CK(clknet_leaf_17_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][8] ),
    .QN(_08992_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[2][9]$_DFFE_PP_  (.D(_01262_),
    .CK(clknet_leaf_17_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[2][9] ),
    .QN(_08991_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][0]$_DFFE_PP_  (.D(_01263_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][0] ),
    .QN(_08990_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][10]$_DFFE_PP_  (.D(_01264_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][10] ),
    .QN(_08989_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][11]$_DFFE_PP_  (.D(_01265_),
    .CK(clknet_leaf_324_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][11] ),
    .QN(_08988_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][12]$_DFFE_PP_  (.D(_01266_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][12] ),
    .QN(_08987_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][13]$_DFFE_PP_  (.D(_01267_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][13] ),
    .QN(_08986_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][14]$_DFFE_PP_  (.D(_01268_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][14] ),
    .QN(_08985_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][15]$_DFFE_PP_  (.D(_01269_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][15] ),
    .QN(_08984_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][16]$_DFFE_PP_  (.D(_01270_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][16] ),
    .QN(_08983_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][17]$_DFFE_PP_  (.D(_01271_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][17] ),
    .QN(_08982_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][18]$_DFFE_PP_  (.D(_01272_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][18] ),
    .QN(_08981_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][19]$_DFFE_PP_  (.D(_01273_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][19] ),
    .QN(_08980_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][1]$_DFFE_PP_  (.D(_01274_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][1] ),
    .QN(_08979_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][20]$_DFFE_PP_  (.D(_01275_),
    .CK(clknet_leaf_323_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][20] ),
    .QN(_08978_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][21]$_DFFE_PP_  (.D(_01276_),
    .CK(clknet_leaf_28_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][21] ),
    .QN(_08977_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][22]$_DFFE_PP_  (.D(_01277_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][22] ),
    .QN(_08976_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][23]$_DFFE_PP_  (.D(_01278_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][23] ),
    .QN(_08975_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][24]$_DFFE_PP_  (.D(_01279_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][24] ),
    .QN(_08974_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][25]$_DFFE_PP_  (.D(_01280_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][25] ),
    .QN(_08973_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][26]$_DFFE_PP_  (.D(_01281_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][26] ),
    .QN(_08972_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][27]$_DFFE_PP_  (.D(_01282_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][27] ),
    .QN(_08971_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][28]$_DFFE_PP_  (.D(_01283_),
    .CK(clknet_leaf_71_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][28] ),
    .QN(_08970_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][29]$_DFFE_PP_  (.D(_01284_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][29] ),
    .QN(_08969_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][2]$_DFFE_PP_  (.D(_01285_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][2] ),
    .QN(_08968_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][30]$_DFFE_PP_  (.D(_01286_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][30] ),
    .QN(_08967_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][31]$_DFFE_PP_  (.D(_01287_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][31] ),
    .QN(_08966_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][32]$_DFFE_PP_  (.D(_01288_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][32] ),
    .QN(_08965_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][33]$_DFFE_PP_  (.D(_01289_),
    .CK(clknet_leaf_76_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][33] ),
    .QN(_08964_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][34]$_DFFE_PP_  (.D(_01290_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][34] ),
    .QN(_08963_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][35]$_DFFE_PP_  (.D(_01291_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][35] ),
    .QN(_08962_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][36]$_DFFE_PP_  (.D(_01292_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][36] ),
    .QN(_08961_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][37]$_DFFE_PP_  (.D(_01293_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][37] ),
    .QN(_08960_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][38]$_DFFE_PP_  (.D(_01294_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][38] ),
    .QN(_08959_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][39]$_DFFE_PP_  (.D(_01295_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][39] ),
    .QN(_08958_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][3]$_DFFE_PP_  (.D(_01296_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][3] ),
    .QN(_08957_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][40]$_DFFE_PP_  (.D(_01297_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][40] ),
    .QN(_08956_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][41]$_DFFE_PP_  (.D(_01298_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][41] ),
    .QN(_08955_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][42]$_DFFE_PP_  (.D(_01299_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][42] ),
    .QN(_08954_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][43]$_DFFE_PP_  (.D(_01300_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][43] ),
    .QN(_08953_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][44]$_DFFE_PP_  (.D(_01301_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][44] ),
    .QN(_08952_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][45]$_DFFE_PP_  (.D(_01302_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][45] ),
    .QN(_08951_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][46]$_DFFE_PP_  (.D(_01303_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][46] ),
    .QN(_08950_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][47]$_DFFE_PP_  (.D(_01304_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][47] ),
    .QN(_08949_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][48]$_DFFE_PP_  (.D(_01305_),
    .CK(clknet_leaf_107_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][48] ),
    .QN(_08948_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][49]$_DFFE_PP_  (.D(_01306_),
    .CK(clknet_leaf_114_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][49] ),
    .QN(_08947_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][4]$_DFFE_PP_  (.D(_01307_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][4] ),
    .QN(_08946_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][50]$_DFFE_PP_  (.D(_01308_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][50] ),
    .QN(_08945_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][51]$_DFFE_PP_  (.D(_01309_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][51] ),
    .QN(_08944_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][52]$_DFFE_PP_  (.D(_01310_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][52] ),
    .QN(_08943_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][53]$_DFFE_PP_  (.D(_01311_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][53] ),
    .QN(_08942_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][54]$_DFFE_PP_  (.D(_01312_),
    .CK(clknet_leaf_118_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][54] ),
    .QN(_08941_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][55]$_DFFE_PP_  (.D(_01313_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][55] ),
    .QN(_08940_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][56]$_DFFE_PP_  (.D(_01314_),
    .CK(clknet_leaf_304_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][56] ),
    .QN(_08939_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][57]$_DFFE_PP_  (.D(_01315_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][57] ),
    .QN(_08938_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][58]$_DFFE_PP_  (.D(_01316_),
    .CK(clknet_leaf_129_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][58] ),
    .QN(_08937_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][59]$_DFFE_PP_  (.D(_01317_),
    .CK(clknet_leaf_52_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][59] ),
    .QN(_08936_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][5]$_DFFE_PP_  (.D(_01318_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][5] ),
    .QN(_08935_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][60]$_DFFE_PP_  (.D(_01319_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][60] ),
    .QN(_08934_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][61]$_DFFE_PP_  (.D(_01320_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][61] ),
    .QN(_08933_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][62]$_DFFE_PP_  (.D(_01321_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][62] ),
    .QN(_08932_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][63]$_DFFE_PP_  (.D(_01322_),
    .CK(clknet_leaf_46_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][63] ),
    .QN(_08931_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][6]$_DFFE_PP_  (.D(_01323_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][6] ),
    .QN(_08930_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][7]$_DFFE_PP_  (.D(_01324_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][7] ),
    .QN(_08929_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][8]$_DFFE_PP_  (.D(_01325_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][8] ),
    .QN(_08928_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[3][9]$_DFFE_PP_  (.D(_01326_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[3][9] ),
    .QN(_08927_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][0]$_DFFE_PP_  (.D(_01327_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][0] ),
    .QN(_08926_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][10]$_DFFE_PP_  (.D(_01328_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][10] ),
    .QN(_08925_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][11]$_DFFE_PP_  (.D(_01329_),
    .CK(clknet_leaf_324_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][11] ),
    .QN(_08924_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][12]$_DFFE_PP_  (.D(_01330_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][12] ),
    .QN(_08923_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][13]$_DFFE_PP_  (.D(_01331_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][13] ),
    .QN(_08922_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][14]$_DFFE_PP_  (.D(_01332_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][14] ),
    .QN(_08921_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][15]$_DFFE_PP_  (.D(_01333_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][15] ),
    .QN(_08920_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][16]$_DFFE_PP_  (.D(_01334_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][16] ),
    .QN(_08919_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][17]$_DFFE_PP_  (.D(_01335_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][17] ),
    .QN(_08918_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][18]$_DFFE_PP_  (.D(_01336_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][18] ),
    .QN(_08917_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][19]$_DFFE_PP_  (.D(_01337_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][19] ),
    .QN(_08916_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][1]$_DFFE_PP_  (.D(_01338_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][1] ),
    .QN(_08915_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][20]$_DFFE_PP_  (.D(_01339_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][20] ),
    .QN(_08914_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][21]$_DFFE_PP_  (.D(_01340_),
    .CK(clknet_leaf_36_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][21] ),
    .QN(_08913_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][22]$_DFFE_PP_  (.D(_01341_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][22] ),
    .QN(_08912_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][23]$_DFFE_PP_  (.D(_01342_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][23] ),
    .QN(_08911_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][24]$_DFFE_PP_  (.D(_01343_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][24] ),
    .QN(_08910_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][25]$_DFFE_PP_  (.D(_01344_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][25] ),
    .QN(_08909_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][26]$_DFFE_PP_  (.D(_01345_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][26] ),
    .QN(_08908_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][27]$_DFFE_PP_  (.D(_01346_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][27] ),
    .QN(_08907_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][28]$_DFFE_PP_  (.D(_01347_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][28] ),
    .QN(_08906_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][29]$_DFFE_PP_  (.D(_01348_),
    .CK(clknet_leaf_71_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][29] ),
    .QN(_08905_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][2]$_DFFE_PP_  (.D(_01349_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][2] ),
    .QN(_08904_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][30]$_DFFE_PP_  (.D(_01350_),
    .CK(clknet_leaf_80_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][30] ),
    .QN(_08903_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][31]$_DFFE_PP_  (.D(_01351_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][31] ),
    .QN(_08902_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][32]$_DFFE_PP_  (.D(_01352_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][32] ),
    .QN(_08901_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][33]$_DFFE_PP_  (.D(_01353_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][33] ),
    .QN(_08900_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][34]$_DFFE_PP_  (.D(_01354_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][34] ),
    .QN(_08899_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][35]$_DFFE_PP_  (.D(_01355_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][35] ),
    .QN(_08898_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][36]$_DFFE_PP_  (.D(_01356_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][36] ),
    .QN(_08897_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][37]$_DFFE_PP_  (.D(_01357_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][37] ),
    .QN(_08896_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][38]$_DFFE_PP_  (.D(_01358_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][38] ),
    .QN(_08895_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][39]$_DFFE_PP_  (.D(_01359_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][39] ),
    .QN(_08894_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][3]$_DFFE_PP_  (.D(_01360_),
    .CK(clknet_leaf_78_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][3] ),
    .QN(_08893_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][40]$_DFFE_PP_  (.D(_01361_),
    .CK(clknet_leaf_102_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][40] ),
    .QN(_08892_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][41]$_DFFE_PP_  (.D(_01362_),
    .CK(clknet_leaf_92_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][41] ),
    .QN(_08891_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][42]$_DFFE_PP_  (.D(_01363_),
    .CK(clknet_leaf_82_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][42] ),
    .QN(_08890_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][43]$_DFFE_PP_  (.D(_01364_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][43] ),
    .QN(_08889_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][44]$_DFFE_PP_  (.D(_01365_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][44] ),
    .QN(_08888_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][45]$_DFFE_PP_  (.D(_01366_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][45] ),
    .QN(_08887_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][46]$_DFFE_PP_  (.D(_01367_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][46] ),
    .QN(_08886_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][47]$_DFFE_PP_  (.D(_01368_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][47] ),
    .QN(_08885_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][48]$_DFFE_PP_  (.D(_01369_),
    .CK(clknet_leaf_92_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][48] ),
    .QN(_08884_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][49]$_DFFE_PP_  (.D(_01370_),
    .CK(clknet_leaf_112_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][49] ),
    .QN(_08883_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][4]$_DFFE_PP_  (.D(_01371_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][4] ),
    .QN(_08882_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][50]$_DFFE_PP_  (.D(_01372_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][50] ),
    .QN(_08881_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][51]$_DFFE_PP_  (.D(_01373_),
    .CK(clknet_leaf_60_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][51] ),
    .QN(_08880_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][52]$_DFFE_PP_  (.D(_01374_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][52] ),
    .QN(_08879_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][53]$_DFFE_PP_  (.D(_01375_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][53] ),
    .QN(_08878_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][54]$_DFFE_PP_  (.D(_01376_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][54] ),
    .QN(_08877_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][55]$_DFFE_PP_  (.D(_01377_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][55] ),
    .QN(_08876_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][56]$_DFFE_PP_  (.D(_01378_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][56] ),
    .QN(_08875_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][57]$_DFFE_PP_  (.D(_01379_),
    .CK(clknet_leaf_42_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][57] ),
    .QN(_08874_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][58]$_DFFE_PP_  (.D(_01380_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][58] ),
    .QN(_08873_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][59]$_DFFE_PP_  (.D(_01381_),
    .CK(clknet_leaf_48_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][59] ),
    .QN(_08872_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][5]$_DFFE_PP_  (.D(_01382_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][5] ),
    .QN(_08871_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][60]$_DFFE_PP_  (.D(_01383_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][60] ),
    .QN(_08870_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][61]$_DFFE_PP_  (.D(_01384_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][61] ),
    .QN(_08869_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][62]$_DFFE_PP_  (.D(_01385_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][62] ),
    .QN(_08868_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][63]$_DFFE_PP_  (.D(_01386_),
    .CK(clknet_leaf_307_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][63] ),
    .QN(_08867_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][6]$_DFFE_PP_  (.D(_01387_),
    .CK(clknet_leaf_20_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][6] ),
    .QN(_08866_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][7]$_DFFE_PP_  (.D(_01388_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][7] ),
    .QN(_08865_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][8]$_DFFE_PP_  (.D(_01389_),
    .CK(clknet_leaf_23_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][8] ),
    .QN(_08864_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[4][9]$_DFFE_PP_  (.D(_01390_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[4][9] ),
    .QN(_08863_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][0]$_DFFE_PP_  (.D(_01391_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][0] ),
    .QN(_08862_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][10]$_DFFE_PP_  (.D(_01392_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][10] ),
    .QN(_08861_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][11]$_DFFE_PP_  (.D(_01393_),
    .CK(clknet_leaf_324_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][11] ),
    .QN(_08860_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][12]$_DFFE_PP_  (.D(_01394_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][12] ),
    .QN(_08859_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][13]$_DFFE_PP_  (.D(_01395_),
    .CK(clknet_leaf_325_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][13] ),
    .QN(_08858_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][14]$_DFFE_PP_  (.D(_01396_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][14] ),
    .QN(_08857_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][15]$_DFFE_PP_  (.D(_01397_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][15] ),
    .QN(_08856_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][16]$_DFFE_PP_  (.D(_01398_),
    .CK(clknet_leaf_325_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][16] ),
    .QN(_08855_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][17]$_DFFE_PP_  (.D(_01399_),
    .CK(clknet_leaf_325_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][17] ),
    .QN(_08854_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][18]$_DFFE_PP_  (.D(_01400_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][18] ),
    .QN(_08853_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][19]$_DFFE_PP_  (.D(_01401_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][19] ),
    .QN(_08852_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][1]$_DFFE_PP_  (.D(_01402_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][1] ),
    .QN(_08851_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][20]$_DFFE_PP_  (.D(_01403_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][20] ),
    .QN(_08850_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][21]$_DFFE_PP_  (.D(_01404_),
    .CK(clknet_leaf_40_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][21] ),
    .QN(_08849_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][22]$_DFFE_PP_  (.D(_01405_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][22] ),
    .QN(_08848_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][23]$_DFFE_PP_  (.D(_01406_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][23] ),
    .QN(_08847_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][24]$_DFFE_PP_  (.D(_01407_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][24] ),
    .QN(_08846_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][25]$_DFFE_PP_  (.D(_01408_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][25] ),
    .QN(_08845_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][26]$_DFFE_PP_  (.D(_01409_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][26] ),
    .QN(_08844_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][27]$_DFFE_PP_  (.D(_01410_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][27] ),
    .QN(_08843_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][28]$_DFFE_PP_  (.D(_01411_),
    .CK(clknet_leaf_26_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][28] ),
    .QN(_08842_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][29]$_DFFE_PP_  (.D(_01412_),
    .CK(clknet_leaf_71_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][29] ),
    .QN(_08841_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][2]$_DFFE_PP_  (.D(_01413_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][2] ),
    .QN(_08840_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][30]$_DFFE_PP_  (.D(_01414_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][30] ),
    .QN(_08839_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][31]$_DFFE_PP_  (.D(_01415_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][31] ),
    .QN(_08838_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][32]$_DFFE_PP_  (.D(_01416_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][32] ),
    .QN(_08837_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][33]$_DFFE_PP_  (.D(_01417_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][33] ),
    .QN(_08836_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][34]$_DFFE_PP_  (.D(_01418_),
    .CK(clknet_leaf_82_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][34] ),
    .QN(_08835_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][35]$_DFFE_PP_  (.D(_01419_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][35] ),
    .QN(_08834_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][36]$_DFFE_PP_  (.D(_01420_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][36] ),
    .QN(_08833_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][37]$_DFFE_PP_  (.D(_01421_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][37] ),
    .QN(_08832_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][38]$_DFFE_PP_  (.D(_01422_),
    .CK(clknet_leaf_103_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][38] ),
    .QN(_08831_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][39]$_DFFE_PP_  (.D(_01423_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][39] ),
    .QN(_08830_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][3]$_DFFE_PP_  (.D(_01424_),
    .CK(clknet_leaf_78_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][3] ),
    .QN(_08829_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][40]$_DFFE_PP_  (.D(_01425_),
    .CK(clknet_leaf_103_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][40] ),
    .QN(_08828_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][41]$_DFFE_PP_  (.D(_01426_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][41] ),
    .QN(_08827_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][42]$_DFFE_PP_  (.D(_01427_),
    .CK(clknet_leaf_82_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][42] ),
    .QN(_08826_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][43]$_DFFE_PP_  (.D(_01428_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][43] ),
    .QN(_08825_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][44]$_DFFE_PP_  (.D(_01429_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][44] ),
    .QN(_08824_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][45]$_DFFE_PP_  (.D(_01430_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][45] ),
    .QN(_08823_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][46]$_DFFE_PP_  (.D(_01431_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][46] ),
    .QN(_08822_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][47]$_DFFE_PP_  (.D(_01432_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][47] ),
    .QN(_08821_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][48]$_DFFE_PP_  (.D(_01433_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][48] ),
    .QN(_08820_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][49]$_DFFE_PP_  (.D(_01434_),
    .CK(clknet_leaf_112_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][49] ),
    .QN(_08819_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][4]$_DFFE_PP_  (.D(_01435_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][4] ),
    .QN(_08818_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][50]$_DFFE_PP_  (.D(_01436_),
    .CK(clknet_leaf_118_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][50] ),
    .QN(_08817_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][51]$_DFFE_PP_  (.D(_01437_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][51] ),
    .QN(_08816_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][52]$_DFFE_PP_  (.D(_01438_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][52] ),
    .QN(_08815_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][53]$_DFFE_PP_  (.D(_01439_),
    .CK(clknet_leaf_116_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][53] ),
    .QN(_08814_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][54]$_DFFE_PP_  (.D(_01440_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][54] ),
    .QN(_08813_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][55]$_DFFE_PP_  (.D(_01441_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][55] ),
    .QN(_08812_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][56]$_DFFE_PP_  (.D(_01442_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][56] ),
    .QN(_08811_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][57]$_DFFE_PP_  (.D(_01443_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][57] ),
    .QN(_08810_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][58]$_DFFE_PP_  (.D(_01444_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][58] ),
    .QN(_08809_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][59]$_DFFE_PP_  (.D(_01445_),
    .CK(clknet_leaf_50_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][59] ),
    .QN(_08808_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][5]$_DFFE_PP_  (.D(_01446_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][5] ),
    .QN(_08807_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][60]$_DFFE_PP_  (.D(_01447_),
    .CK(clknet_leaf_47_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][60] ),
    .QN(_08806_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][61]$_DFFE_PP_  (.D(_01448_),
    .CK(clknet_leaf_45_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][61] ),
    .QN(_08805_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][62]$_DFFE_PP_  (.D(_01449_),
    .CK(clknet_leaf_48_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][62] ),
    .QN(_08804_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][63]$_DFFE_PP_  (.D(_01450_),
    .CK(clknet_leaf_305_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][63] ),
    .QN(_08803_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][6]$_DFFE_PP_  (.D(_01451_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][6] ),
    .QN(_08802_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][7]$_DFFE_PP_  (.D(_01452_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][7] ),
    .QN(_08801_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][8]$_DFFE_PP_  (.D(_01453_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][8] ),
    .QN(_08800_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[5][9]$_DFFE_PP_  (.D(_01454_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[5][9] ),
    .QN(_08799_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][0]$_DFFE_PP_  (.D(_01455_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][0] ),
    .QN(_08798_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][10]$_DFFE_PP_  (.D(_01456_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][10] ),
    .QN(_08797_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][11]$_DFFE_PP_  (.D(_01457_),
    .CK(clknet_leaf_324_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][11] ),
    .QN(_08796_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][12]$_DFFE_PP_  (.D(_01458_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][12] ),
    .QN(_08795_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][13]$_DFFE_PP_  (.D(_01459_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][13] ),
    .QN(_08794_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][14]$_DFFE_PP_  (.D(_01460_),
    .CK(clknet_leaf_11_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][14] ),
    .QN(_08793_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][15]$_DFFE_PP_  (.D(_01461_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][15] ),
    .QN(_08792_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][16]$_DFFE_PP_  (.D(_01462_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][16] ),
    .QN(_08791_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][17]$_DFFE_PP_  (.D(_01463_),
    .CK(clknet_leaf_326_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][17] ),
    .QN(_08790_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][18]$_DFFE_PP_  (.D(_01464_),
    .CK(clknet_leaf_15_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][18] ),
    .QN(_08789_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][19]$_DFFE_PP_  (.D(_01465_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][19] ),
    .QN(_08788_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][1]$_DFFE_PP_  (.D(_01466_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][1] ),
    .QN(_08787_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][20]$_DFFE_PP_  (.D(_01467_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][20] ),
    .QN(_08786_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][21]$_DFFE_PP_  (.D(_01468_),
    .CK(clknet_leaf_36_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][21] ),
    .QN(_08785_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][22]$_DFFE_PP_  (.D(_01469_),
    .CK(clknet_leaf_315_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][22] ),
    .QN(_08784_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][23]$_DFFE_PP_  (.D(_01470_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][23] ),
    .QN(_08783_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][24]$_DFFE_PP_  (.D(_01471_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][24] ),
    .QN(_08782_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][25]$_DFFE_PP_  (.D(_01472_),
    .CK(clknet_leaf_311_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][25] ),
    .QN(_08781_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][26]$_DFFE_PP_  (.D(_01473_),
    .CK(clknet_leaf_37_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][26] ),
    .QN(_08780_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][27]$_DFFE_PP_  (.D(_01474_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][27] ),
    .QN(_08779_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][28]$_DFFE_PP_  (.D(_01475_),
    .CK(clknet_leaf_71_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][28] ),
    .QN(_08778_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][29]$_DFFE_PP_  (.D(_01476_),
    .CK(clknet_leaf_71_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][29] ),
    .QN(_08777_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][2]$_DFFE_PP_  (.D(_01477_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][2] ),
    .QN(_08776_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][30]$_DFFE_PP_  (.D(_01478_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][30] ),
    .QN(_08775_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][31]$_DFFE_PP_  (.D(_01479_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][31] ),
    .QN(_08774_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][32]$_DFFE_PP_  (.D(_01480_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][32] ),
    .QN(_08773_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][33]$_DFFE_PP_  (.D(_01481_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][33] ),
    .QN(_08772_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][34]$_DFFE_PP_  (.D(_01482_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][34] ),
    .QN(_08771_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][35]$_DFFE_PP_  (.D(_01483_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][35] ),
    .QN(_08770_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][36]$_DFFE_PP_  (.D(_01484_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][36] ),
    .QN(_08769_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][37]$_DFFE_PP_  (.D(_01485_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][37] ),
    .QN(_08768_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][38]$_DFFE_PP_  (.D(_01486_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][38] ),
    .QN(_08767_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][39]$_DFFE_PP_  (.D(_01487_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][39] ),
    .QN(_08766_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][3]$_DFFE_PP_  (.D(_01488_),
    .CK(clknet_leaf_78_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][3] ),
    .QN(_08765_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][40]$_DFFE_PP_  (.D(_01489_),
    .CK(clknet_leaf_103_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][40] ),
    .QN(_08764_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][41]$_DFFE_PP_  (.D(_01490_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][41] ),
    .QN(_08763_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][42]$_DFFE_PP_  (.D(_01491_),
    .CK(clknet_leaf_82_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][42] ),
    .QN(_08762_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][43]$_DFFE_PP_  (.D(_01492_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][43] ),
    .QN(_08761_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][44]$_DFFE_PP_  (.D(_01493_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][44] ),
    .QN(_08760_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][45]$_DFFE_PP_  (.D(_01494_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][45] ),
    .QN(_08759_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][46]$_DFFE_PP_  (.D(_01495_),
    .CK(clknet_leaf_91_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][46] ),
    .QN(_08758_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][47]$_DFFE_PP_  (.D(_01496_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][47] ),
    .QN(_08757_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][48]$_DFFE_PP_  (.D(_01497_),
    .CK(clknet_leaf_92_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][48] ),
    .QN(_08756_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][49]$_DFFE_PP_  (.D(_01498_),
    .CK(clknet_leaf_112_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][49] ),
    .QN(_08755_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][4]$_DFFE_PP_  (.D(_01499_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][4] ),
    .QN(_08754_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][50]$_DFFE_PP_  (.D(_01500_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][50] ),
    .QN(_08753_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][51]$_DFFE_PP_  (.D(_01501_),
    .CK(clknet_leaf_58_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][51] ),
    .QN(_08752_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][52]$_DFFE_PP_  (.D(_01502_),
    .CK(clknet_leaf_119_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][52] ),
    .QN(_08751_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][53]$_DFFE_PP_  (.D(_01503_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][53] ),
    .QN(_08750_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][54]$_DFFE_PP_  (.D(_01504_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][54] ),
    .QN(_08749_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][55]$_DFFE_PP_  (.D(_01505_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][55] ),
    .QN(_08748_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][56]$_DFFE_PP_  (.D(_01506_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][56] ),
    .QN(_08747_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][57]$_DFFE_PP_  (.D(_01507_),
    .CK(clknet_leaf_55_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][57] ),
    .QN(_08746_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][58]$_DFFE_PP_  (.D(_01508_),
    .CK(clknet_leaf_50_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][58] ),
    .QN(_08745_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][59]$_DFFE_PP_  (.D(_01509_),
    .CK(clknet_leaf_48_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][59] ),
    .QN(_08744_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][5]$_DFFE_PP_  (.D(_01510_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][5] ),
    .QN(_08743_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][60]$_DFFE_PP_  (.D(_01511_),
    .CK(clknet_leaf_46_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][60] ),
    .QN(_08742_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][61]$_DFFE_PP_  (.D(_01512_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][61] ),
    .QN(_08741_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][62]$_DFFE_PP_  (.D(_01513_),
    .CK(clknet_leaf_302_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][62] ),
    .QN(_08740_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][63]$_DFFE_PP_  (.D(_01514_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][63] ),
    .QN(_08739_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][6]$_DFFE_PP_  (.D(_01515_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][6] ),
    .QN(_08738_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][7]$_DFFE_PP_  (.D(_01516_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][7] ),
    .QN(_08737_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][8]$_DFFE_PP_  (.D(_01517_),
    .CK(clknet_leaf_22_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][8] ),
    .QN(_08736_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[6][9]$_DFFE_PP_  (.D(_01518_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[6][9] ),
    .QN(_08735_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][0]$_DFFE_PP_  (.D(_01519_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][0] ),
    .QN(_08734_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][10]$_DFFE_PP_  (.D(_01520_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][10] ),
    .QN(_08733_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][11]$_DFFE_PP_  (.D(_01521_),
    .CK(clknet_leaf_325_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][11] ),
    .QN(_08732_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][12]$_DFFE_PP_  (.D(_01522_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][12] ),
    .QN(_08731_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][13]$_DFFE_PP_  (.D(_01523_),
    .CK(clknet_leaf_325_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][13] ),
    .QN(_08730_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][14]$_DFFE_PP_  (.D(_01524_),
    .CK(clknet_leaf_13_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][14] ),
    .QN(_08729_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][15]$_DFFE_PP_  (.D(_01525_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][15] ),
    .QN(_08728_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][16]$_DFFE_PP_  (.D(_01526_),
    .CK(clknet_leaf_325_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][16] ),
    .QN(_08727_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][17]$_DFFE_PP_  (.D(_01527_),
    .CK(clknet_leaf_12_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][17] ),
    .QN(_08726_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][18]$_DFFE_PP_  (.D(_01528_),
    .CK(clknet_leaf_14_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][18] ),
    .QN(_08725_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][19]$_DFFE_PP_  (.D(_01529_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][19] ),
    .QN(_08724_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][1]$_DFFE_PP_  (.D(_01530_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][1] ),
    .QN(_08723_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][20]$_DFFE_PP_  (.D(_01531_),
    .CK(clknet_leaf_321_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][20] ),
    .QN(_08722_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][21]$_DFFE_PP_  (.D(_01532_),
    .CK(clknet_leaf_40_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][21] ),
    .QN(_08721_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][22]$_DFFE_PP_  (.D(_01533_),
    .CK(clknet_leaf_313_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][22] ),
    .QN(_08720_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][23]$_DFFE_PP_  (.D(_01534_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][23] ),
    .QN(_08719_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][24]$_DFFE_PP_  (.D(_01535_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][24] ),
    .QN(_08718_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][25]$_DFFE_PP_  (.D(_01536_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][25] ),
    .QN(_08717_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][26]$_DFFE_PP_  (.D(_01537_),
    .CK(clknet_leaf_37_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][26] ),
    .QN(_08716_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][27]$_DFFE_PP_  (.D(_01538_),
    .CK(clknet_leaf_319_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][27] ),
    .QN(_08715_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][28]$_DFFE_PP_  (.D(_01539_),
    .CK(clknet_leaf_72_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][28] ),
    .QN(_08714_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][29]$_DFFE_PP_  (.D(_01540_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][29] ),
    .QN(_08713_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][2]$_DFFE_PP_  (.D(_01541_),
    .CK(clknet_leaf_77_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][2] ),
    .QN(_08712_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][30]$_DFFE_PP_  (.D(_01542_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][30] ),
    .QN(_08711_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][31]$_DFFE_PP_  (.D(_01543_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][31] ),
    .QN(_08710_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][32]$_DFFE_PP_  (.D(_01544_),
    .CK(clknet_leaf_66_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][32] ),
    .QN(_08709_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][33]$_DFFE_PP_  (.D(_01545_),
    .CK(clknet_leaf_78_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][33] ),
    .QN(_08708_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][34]$_DFFE_PP_  (.D(_01546_),
    .CK(clknet_leaf_82_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][34] ),
    .QN(_08707_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][35]$_DFFE_PP_  (.D(_01547_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][35] ),
    .QN(_08706_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][36]$_DFFE_PP_  (.D(_01548_),
    .CK(clknet_leaf_89_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][36] ),
    .QN(_08705_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][37]$_DFFE_PP_  (.D(_01549_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][37] ),
    .QN(_08704_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][38]$_DFFE_PP_  (.D(_01550_),
    .CK(clknet_leaf_103_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][38] ),
    .QN(_08703_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][39]$_DFFE_PP_  (.D(_01551_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][39] ),
    .QN(_08702_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][3]$_DFFE_PP_  (.D(_01552_),
    .CK(clknet_leaf_78_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][3] ),
    .QN(_08701_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][40]$_DFFE_PP_  (.D(_01553_),
    .CK(clknet_leaf_103_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][40] ),
    .QN(_08700_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][41]$_DFFE_PP_  (.D(_01554_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][41] ),
    .QN(_08699_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][42]$_DFFE_PP_  (.D(_01555_),
    .CK(clknet_leaf_83_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][42] ),
    .QN(_08698_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][43]$_DFFE_PP_  (.D(_01556_),
    .CK(clknet_leaf_100_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][43] ),
    .QN(_08697_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][44]$_DFFE_PP_  (.D(_01557_),
    .CK(clknet_leaf_84_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][44] ),
    .QN(_08696_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][45]$_DFFE_PP_  (.D(_01558_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][45] ),
    .QN(_08695_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][46]$_DFFE_PP_  (.D(_01559_),
    .CK(clknet_leaf_92_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][46] ),
    .QN(_08694_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][47]$_DFFE_PP_  (.D(_01560_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][47] ),
    .QN(_08693_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][48]$_DFFE_PP_  (.D(_01561_),
    .CK(clknet_leaf_105_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][48] ),
    .QN(_08692_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][49]$_DFFE_PP_  (.D(_01562_),
    .CK(clknet_leaf_112_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][49] ),
    .QN(_08691_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][4]$_DFFE_PP_  (.D(_01563_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][4] ),
    .QN(_08690_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][50]$_DFFE_PP_  (.D(_01564_),
    .CK(clknet_leaf_118_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][50] ),
    .QN(_08689_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][51]$_DFFE_PP_  (.D(_01565_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][51] ),
    .QN(_08688_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][52]$_DFFE_PP_  (.D(_01566_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][52] ),
    .QN(_08687_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][53]$_DFFE_PP_  (.D(_01567_),
    .CK(clknet_leaf_116_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][53] ),
    .QN(_08686_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][54]$_DFFE_PP_  (.D(_01568_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][54] ),
    .QN(_08685_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][55]$_DFFE_PP_  (.D(_01569_),
    .CK(clknet_leaf_44_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][55] ),
    .QN(_08684_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][56]$_DFFE_PP_  (.D(_01570_),
    .CK(clknet_leaf_300_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][56] ),
    .QN(_08683_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][57]$_DFFE_PP_  (.D(_01571_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][57] ),
    .QN(_08682_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][58]$_DFFE_PP_  (.D(_01572_),
    .CK(clknet_leaf_131_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][58] ),
    .QN(_08681_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][59]$_DFFE_PP_  (.D(_01573_),
    .CK(clknet_leaf_50_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][59] ),
    .QN(_08680_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][5]$_DFFE_PP_  (.D(_01574_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][5] ),
    .QN(_08679_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][60]$_DFFE_PP_  (.D(_01575_),
    .CK(clknet_leaf_46_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][60] ),
    .QN(_08678_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][61]$_DFFE_PP_  (.D(_01576_),
    .CK(clknet_leaf_43_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][61] ),
    .QN(_08677_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][62]$_DFFE_PP_  (.D(_01577_),
    .CK(clknet_leaf_49_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][62] ),
    .QN(_08676_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][63]$_DFFE_PP_  (.D(_01578_),
    .CK(clknet_leaf_46_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][63] ),
    .QN(_08675_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][6]$_DFFE_PP_  (.D(_01579_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][6] ),
    .QN(_08674_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][7]$_DFFE_PP_  (.D(_01580_),
    .CK(clknet_leaf_19_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][7] ),
    .QN(_08673_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][8]$_DFFE_PP_  (.D(_01581_),
    .CK(clknet_leaf_17_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][8] ),
    .QN(_08672_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[7][9]$_DFFE_PP_  (.D(_01582_),
    .CK(clknet_leaf_18_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[7][9] ),
    .QN(_08671_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][0]$_DFFE_PP_  (.D(_01583_),
    .CK(clknet_leaf_30_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][0] ),
    .QN(_08670_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][10]$_DFFE_PP_  (.D(_01584_),
    .CK(clknet_leaf_6_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][10] ),
    .QN(_08669_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][11]$_DFFE_PP_  (.D(_01585_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][11] ),
    .QN(_08668_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][12]$_DFFE_PP_  (.D(_01586_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][12] ),
    .QN(_08667_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][13]$_DFFE_PP_  (.D(_01587_),
    .CK(clknet_leaf_1_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][13] ),
    .QN(_08666_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][14]$_DFFE_PP_  (.D(_01588_),
    .CK(clknet_leaf_6_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][14] ),
    .QN(_08665_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][15]$_DFFE_PP_  (.D(_01589_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][15] ),
    .QN(_08664_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][16]$_DFFE_PP_  (.D(_01590_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][16] ),
    .QN(_08663_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][17]$_DFFE_PP_  (.D(_01591_),
    .CK(clknet_leaf_2_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][17] ),
    .QN(_08662_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][18]$_DFFE_PP_  (.D(_01592_),
    .CK(clknet_leaf_7_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][18] ),
    .QN(_08661_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][19]$_DFFE_PP_  (.D(_01593_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][19] ),
    .QN(_08660_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][1]$_DFFE_PP_  (.D(_01594_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][1] ),
    .QN(_08659_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][20]$_DFFE_PP_  (.D(_01595_),
    .CK(clknet_leaf_4_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][20] ),
    .QN(_08658_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][21]$_DFFE_PP_  (.D(_01596_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][21] ),
    .QN(_08657_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][22]$_DFFE_PP_  (.D(_01597_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][22] ),
    .QN(_08656_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][23]$_DFFE_PP_  (.D(_01598_),
    .CK(clknet_leaf_309_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][23] ),
    .QN(_08655_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][24]$_DFFE_PP_  (.D(_01599_),
    .CK(clknet_leaf_316_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][24] ),
    .QN(_08654_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][25]$_DFFE_PP_  (.D(_01600_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][25] ),
    .QN(_08653_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][26]$_DFFE_PP_  (.D(_01601_),
    .CK(clknet_leaf_37_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][26] ),
    .QN(_08652_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][27]$_DFFE_PP_  (.D(_01602_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][27] ),
    .QN(_08651_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][28]$_DFFE_PP_  (.D(_01603_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][28] ),
    .QN(_08650_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][29]$_DFFE_PP_  (.D(_01604_),
    .CK(clknet_leaf_56_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][29] ),
    .QN(_08649_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][2]$_DFFE_PP_  (.D(_01605_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][2] ),
    .QN(_08648_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][30]$_DFFE_PP_  (.D(_01606_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][30] ),
    .QN(_08647_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][31]$_DFFE_PP_  (.D(_01607_),
    .CK(clknet_leaf_65_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][31] ),
    .QN(_08646_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][32]$_DFFE_PP_  (.D(_01608_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][32] ),
    .QN(_08645_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][33]$_DFFE_PP_  (.D(_01609_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][33] ),
    .QN(_08644_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][34]$_DFFE_PP_  (.D(_01610_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][34] ),
    .QN(_08643_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][35]$_DFFE_PP_  (.D(_01611_),
    .CK(clknet_leaf_88_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][35] ),
    .QN(_08642_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][36]$_DFFE_PP_  (.D(_01612_),
    .CK(clknet_leaf_61_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][36] ),
    .QN(_08641_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][37]$_DFFE_PP_  (.D(_01613_),
    .CK(clknet_leaf_94_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][37] ),
    .QN(_08640_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][38]$_DFFE_PP_  (.D(_01614_),
    .CK(clknet_leaf_97_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][38] ),
    .QN(_08639_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][39]$_DFFE_PP_  (.D(_01615_),
    .CK(clknet_leaf_86_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][39] ),
    .QN(_08638_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][3]$_DFFE_PP_  (.D(_01616_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][3] ),
    .QN(_08637_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][40]$_DFFE_PP_  (.D(_01617_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][40] ),
    .QN(_08636_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][41]$_DFFE_PP_  (.D(_01618_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][41] ),
    .QN(_08635_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][42]$_DFFE_PP_  (.D(_01619_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][42] ),
    .QN(_08634_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][43]$_DFFE_PP_  (.D(_01620_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][43] ),
    .QN(_08633_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][44]$_DFFE_PP_  (.D(_01621_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][44] ),
    .QN(_08632_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][45]$_DFFE_PP_  (.D(_01622_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][45] ),
    .QN(_08631_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][46]$_DFFE_PP_  (.D(_01623_),
    .CK(clknet_leaf_62_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][46] ),
    .QN(_08630_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][47]$_DFFE_PP_  (.D(_01624_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][47] ),
    .QN(_08629_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][48]$_DFFE_PP_  (.D(_01625_),
    .CK(clknet_leaf_115_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][48] ),
    .QN(_08628_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][49]$_DFFE_PP_  (.D(_01626_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][49] ),
    .QN(_08627_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][4]$_DFFE_PP_  (.D(_01627_),
    .CK(clknet_leaf_56_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][4] ),
    .QN(_08626_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][50]$_DFFE_PP_  (.D(_01628_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][50] ),
    .QN(_08625_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][51]$_DFFE_PP_  (.D(_01629_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][51] ),
    .QN(_08624_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][52]$_DFFE_PP_  (.D(_01630_),
    .CK(clknet_leaf_127_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][52] ),
    .QN(_08623_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][53]$_DFFE_PP_  (.D(_01631_),
    .CK(clknet_leaf_121_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][53] ),
    .QN(_08622_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][54]$_DFFE_PP_  (.D(_01632_),
    .CK(clknet_leaf_120_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][54] ),
    .QN(_08621_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][55]$_DFFE_PP_  (.D(_01633_),
    .CK(clknet_leaf_51_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][55] ),
    .QN(_08620_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][56]$_DFFE_PP_  (.D(_01634_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][56] ),
    .QN(_08619_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][57]$_DFFE_PP_  (.D(_01635_),
    .CK(clknet_leaf_51_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][57] ),
    .QN(_08618_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][58]$_DFFE_PP_  (.D(_01636_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][58] ),
    .QN(_08617_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][59]$_DFFE_PP_  (.D(_01637_),
    .CK(clknet_leaf_130_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][59] ),
    .QN(_08616_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][5]$_DFFE_PP_  (.D(_01638_),
    .CK(clknet_leaf_40_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][5] ),
    .QN(_08615_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][60]$_DFFE_PP_  (.D(_01639_),
    .CK(clknet_leaf_308_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][60] ),
    .QN(_08614_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][61]$_DFFE_PP_  (.D(_01640_),
    .CK(clknet_leaf_46_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][61] ),
    .QN(_08613_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][62]$_DFFE_PP_  (.D(_01641_),
    .CK(clknet_leaf_301_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][62] ),
    .QN(_08612_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][63]$_DFFE_PP_  (.D(_01642_),
    .CK(clknet_leaf_306_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][63] ),
    .QN(_08611_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][6]$_DFFE_PP_  (.D(_01643_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][6] ),
    .QN(_08610_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][7]$_DFFE_PP_  (.D(_01644_),
    .CK(clknet_leaf_24_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][7] ),
    .QN(_08609_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][8]$_DFFE_PP_  (.D(_01645_),
    .CK(clknet_leaf_29_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][8] ),
    .QN(_08608_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[8][9]$_DFFE_PP_  (.D(_01646_),
    .CK(clknet_leaf_23_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[8][9] ),
    .QN(_08607_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][0]$_DFFE_PP_  (.D(_01647_),
    .CK(clknet_leaf_16_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][0] ),
    .QN(_08606_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][10]$_DFFE_PP_  (.D(_01648_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][10] ),
    .QN(_08605_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][11]$_DFFE_PP_  (.D(_01649_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][11] ),
    .QN(_08604_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][12]$_DFFE_PP_  (.D(_01650_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][12] ),
    .QN(_08603_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][13]$_DFFE_PP_  (.D(_01651_),
    .CK(clknet_leaf_0_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][13] ),
    .QN(_08602_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][14]$_DFFE_PP_  (.D(_01652_),
    .CK(clknet_leaf_10_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][14] ),
    .QN(_08601_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][15]$_DFFE_PP_  (.D(_01653_),
    .CK(clknet_leaf_9_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][15] ),
    .QN(_08600_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][16]$_DFFE_PP_  (.D(_01654_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][16] ),
    .QN(_08599_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][17]$_DFFE_PP_  (.D(_01655_),
    .CK(clknet_leaf_327_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][17] ),
    .QN(_08598_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][18]$_DFFE_PP_  (.D(_01656_),
    .CK(clknet_leaf_8_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][18] ),
    .QN(_08597_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][19]$_DFFE_PP_  (.D(_01657_),
    .CK(clknet_leaf_34_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][19] ),
    .QN(_08596_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][1]$_DFFE_PP_  (.D(_01658_),
    .CK(clknet_leaf_35_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][1] ),
    .QN(_08595_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][20]$_DFFE_PP_  (.D(_01659_),
    .CK(clknet_leaf_322_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][20] ),
    .QN(_08594_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][21]$_DFFE_PP_  (.D(_01660_),
    .CK(clknet_leaf_32_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][21] ),
    .QN(_08593_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][22]$_DFFE_PP_  (.D(_01661_),
    .CK(clknet_leaf_314_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][22] ),
    .QN(_08592_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][23]$_DFFE_PP_  (.D(_01662_),
    .CK(clknet_leaf_310_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][23] ),
    .QN(_08591_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][24]$_DFFE_PP_  (.D(_01663_),
    .CK(clknet_leaf_317_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][24] ),
    .QN(_08590_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][25]$_DFFE_PP_  (.D(_01664_),
    .CK(clknet_leaf_312_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][25] ),
    .QN(_08589_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][26]$_DFFE_PP_  (.D(_01665_),
    .CK(clknet_leaf_38_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][26] ),
    .QN(_08588_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][27]$_DFFE_PP_  (.D(_01666_),
    .CK(clknet_leaf_318_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][27] ),
    .QN(_08587_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][28]$_DFFE_PP_  (.D(_01667_),
    .CK(clknet_leaf_27_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][28] ),
    .QN(_08586_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][29]$_DFFE_PP_  (.D(_01668_),
    .CK(clknet_leaf_70_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][29] ),
    .QN(_08585_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][2]$_DFFE_PP_  (.D(_01669_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][2] ),
    .QN(_08584_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][30]$_DFFE_PP_  (.D(_01670_),
    .CK(clknet_leaf_73_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][30] ),
    .QN(_08583_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][31]$_DFFE_PP_  (.D(_01671_),
    .CK(clknet_leaf_68_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][31] ),
    .QN(_08582_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][32]$_DFFE_PP_  (.D(_01672_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][32] ),
    .QN(_08581_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][33]$_DFFE_PP_  (.D(_01673_),
    .CK(clknet_leaf_75_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][33] ),
    .QN(_08580_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][34]$_DFFE_PP_  (.D(_01674_),
    .CK(clknet_leaf_81_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][34] ),
    .QN(_08579_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][35]$_DFFE_PP_  (.D(_01675_),
    .CK(clknet_leaf_87_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][35] ),
    .QN(_08578_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][36]$_DFFE_PP_  (.D(_01676_),
    .CK(clknet_leaf_64_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][36] ),
    .QN(_08577_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][37]$_DFFE_PP_  (.D(_01677_),
    .CK(clknet_leaf_104_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][37] ),
    .QN(_08576_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][38]$_DFFE_PP_  (.D(_01678_),
    .CK(clknet_leaf_95_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][38] ),
    .QN(_08575_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][39]$_DFFE_PP_  (.D(_01679_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][39] ),
    .QN(_08574_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][3]$_DFFE_PP_  (.D(_01680_),
    .CK(clknet_leaf_74_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][3] ),
    .QN(_08573_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][40]$_DFFE_PP_  (.D(_01681_),
    .CK(clknet_leaf_96_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][40] ),
    .QN(_08572_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][41]$_DFFE_PP_  (.D(_01682_),
    .CK(clknet_leaf_93_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][41] ),
    .QN(_08571_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][42]$_DFFE_PP_  (.D(_01683_),
    .CK(clknet_leaf_79_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][42] ),
    .QN(_08570_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][43]$_DFFE_PP_  (.D(_01684_),
    .CK(clknet_leaf_99_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][43] ),
    .QN(_08569_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][44]$_DFFE_PP_  (.D(_01685_),
    .CK(clknet_leaf_85_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][44] ),
    .QN(_08568_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][45]$_DFFE_PP_  (.D(_01686_),
    .CK(clknet_leaf_101_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][45] ),
    .QN(_08567_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][46]$_DFFE_PP_  (.D(_01687_),
    .CK(clknet_leaf_63_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][46] ),
    .QN(_08566_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][47]$_DFFE_PP_  (.D(_01688_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][47] ),
    .QN(_08565_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][48]$_DFFE_PP_  (.D(_01689_),
    .CK(clknet_leaf_106_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][48] ),
    .QN(_08564_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][49]$_DFFE_PP_  (.D(_01690_),
    .CK(clknet_leaf_113_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][49] ),
    .QN(_08563_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][4]$_DFFE_PP_  (.D(_01691_),
    .CK(clknet_leaf_69_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][4] ),
    .QN(_08562_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][50]$_DFFE_PP_  (.D(_01692_),
    .CK(clknet_leaf_118_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][50] ),
    .QN(_08561_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][51]$_DFFE_PP_  (.D(_01693_),
    .CK(clknet_leaf_118_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][51] ),
    .QN(_08560_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][52]$_DFFE_PP_  (.D(_01694_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][52] ),
    .QN(_08559_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][53]$_DFFE_PP_  (.D(_01695_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][53] ),
    .QN(_08558_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][54]$_DFFE_PP_  (.D(_01696_),
    .CK(clknet_leaf_117_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][54] ),
    .QN(_08557_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][55]$_DFFE_PP_  (.D(_01697_),
    .CK(clknet_leaf_54_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][55] ),
    .QN(_08556_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][56]$_DFFE_PP_  (.D(_01698_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][56] ),
    .QN(_08555_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][57]$_DFFE_PP_  (.D(_01699_),
    .CK(clknet_leaf_53_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][57] ),
    .QN(_08554_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][58]$_DFFE_PP_  (.D(_01700_),
    .CK(clknet_leaf_129_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][58] ),
    .QN(_08553_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][59]$_DFFE_PP_  (.D(_01701_),
    .CK(clknet_leaf_128_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][59] ),
    .QN(_08552_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][5]$_DFFE_PP_  (.D(_01702_),
    .CK(clknet_leaf_41_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][5] ),
    .QN(_08551_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][60]$_DFFE_PP_  (.D(_01703_),
    .CK(clknet_leaf_304_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][60] ),
    .QN(_08550_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][61]$_DFFE_PP_  (.D(_01704_),
    .CK(clknet_leaf_39_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][61] ),
    .QN(_08549_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][62]$_DFFE_PP_  (.D(_01705_),
    .CK(clknet_leaf_303_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][62] ),
    .QN(_08548_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][63]$_DFFE_PP_  (.D(_01706_),
    .CK(clknet_leaf_305_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][63] ),
    .QN(_08547_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][6]$_DFFE_PP_  (.D(_01707_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][6] ),
    .QN(_08546_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][7]$_DFFE_PP_  (.D(_01708_),
    .CK(clknet_leaf_21_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][7] ),
    .QN(_08545_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][8]$_DFFE_PP_  (.D(_01709_),
    .CK(clknet_leaf_23_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][8] ),
    .QN(_08544_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.storage_data_f[9][9]$_DFFE_PP_  (.D(_01710_),
    .CK(clknet_leaf_23_clk),
    .Q(\dynamic_node_top.proc_input.NIB.storage_data_f[9][9] ),
    .QN(_08543_));
 DFF_X2 \dynamic_node_top.proc_input.NIB.tail_ptr_f[0]$_SDFFE_PP0N_  (.D(_01711_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.tail_ptr_f[0] ),
    .QN(\dynamic_node_top.proc_input.NIB.tail_ptr_next[0] ));
 DFF_X2 \dynamic_node_top.proc_input.NIB.tail_ptr_f[1]$_SDFFE_PP0N_  (.D(_01712_),
    .CK(clknet_leaf_57_clk),
    .Q(\dynamic_node_top.proc_input.NIB.tail_ptr_f[1] ),
    .QN(_10593_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.tail_ptr_f[2]$_SDFFE_PP0N_  (.D(_01713_),
    .CK(clknet_leaf_59_clk),
    .Q(\dynamic_node_top.proc_input.NIB.tail_ptr_f[2] ),
    .QN(_08542_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.tail_ptr_f[3]$_SDFFE_PP0N_  (.D(_01714_),
    .CK(clknet_leaf_60_clk),
    .Q(\dynamic_node_top.proc_input.NIB.tail_ptr_f[3] ),
    .QN(_08541_));
 DFF_X1 \dynamic_node_top.proc_input.NIB.yummy_out_f$_SDFF_PP0_  (.D(_01715_),
    .CK(clknet_leaf_112_clk),
    .Q(net628),
    .QN(_08540_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[0]$_SDFF_PP0_  (.D(_01716_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[0] ),
    .QN(_10531_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[1]$_SDFF_PP0_  (.D(_01717_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[1] ),
    .QN(_10532_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[2]$_SDFF_PP0_  (.D(_01718_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[2] ),
    .QN(_08539_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[3]$_SDFF_PP0_  (.D(_01719_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[3] ),
    .QN(_08538_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[4]$_SDFF_PP0_  (.D(_01720_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[4] ),
    .QN(_08537_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[5]$_SDFF_PP0_  (.D(_01721_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[5] ),
    .QN(_08536_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[6]$_SDFF_PP0_  (.D(_01722_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[6] ),
    .QN(_08535_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_f[7]$_SDFF_PP0_  (.D(_01723_),
    .CK(clknet_leaf_110_clk),
    .Q(\dynamic_node_top.proc_input.control.count_f[7] ),
    .QN(_08534_));
 DFF_X1 \dynamic_node_top.proc_input.control.count_one_f$_SDFF_PP0_  (.D(_01724_),
    .CK(clknet_leaf_111_clk),
    .Q(\dynamic_node_top.proc_input.control.count_one_f ),
    .QN(_10156_));
 DFF_X2 \dynamic_node_top.proc_input.control.header_temp$_DFF_P_  (.D(_00002_),
    .CK(clknet_leaf_109_clk),
    .Q(\dynamic_node_top.proc_input.control.header_last_temp ),
    .QN(_08533_));
 DFF_X1 \dynamic_node_top.proc_input.control.tail_last_f$_SDFF_PP0_  (.D(_01725_),
    .CK(clknet_leaf_111_clk),
    .Q(\dynamic_node_top.proc_input.control.tail_last_f ),
    .QN(_10157_));
 DFF_X1 \dynamic_node_top.proc_output.control.current_route_f[0]$_DFF_P_  (.D(_00022_),
    .CK(clknet_leaf_141_clk),
    .Q(\dynamic_node_top.proc_output.control.current_route_f[0] ),
    .QN(_00054_));
 DFF_X1 \dynamic_node_top.proc_output.control.current_route_f[1]$_DFF_P_  (.D(_00023_),
    .CK(clknet_leaf_159_clk),
    .Q(\dynamic_node_top.proc_output.control.current_route_f[1] ),
    .QN(_00053_));
 DFF_X2 \dynamic_node_top.proc_output.control.current_route_f[2]$_DFF_P_  (.D(_00024_),
    .CK(clknet_leaf_141_clk),
    .Q(\dynamic_node_top.proc_output.control.current_route_f[2] ),
    .QN(_00066_));
 DFF_X1 \dynamic_node_top.proc_output.control.current_route_f[3]$_DFF_P_  (.D(_00025_),
    .CK(clknet_leaf_141_clk),
    .Q(\dynamic_node_top.proc_output.control.current_route_f[3] ),
    .QN(_00067_));
 DFF_X2 \dynamic_node_top.proc_output.control.current_route_f[4]$_DFF_P_  (.D(_00026_),
    .CK(clknet_leaf_159_clk),
    .Q(\dynamic_node_top.proc_output.control.current_route_f[4] ),
    .QN(_00065_));
 DFF_X1 \dynamic_node_top.proc_output.control.planned_f$_SDFF_PP0_  (.D(_01726_),
    .CK(clknet_leaf_143_clk),
    .Q(\dynamic_node_top.proc_output.control.planned_f ),
    .QN(_00055_));
 DFF_X2 \dynamic_node_top.proc_output.space.count_f[0]$_SDFF_PP0_  (.D(_01727_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.proc_output.space.count_f[0] ),
    .QN(_10523_));
 DFF_X2 \dynamic_node_top.proc_output.space.count_f[1]$_SDFF_PP0_  (.D(_01728_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.proc_output.space.count_f[1] ),
    .QN(_10524_));
 DFF_X1 \dynamic_node_top.proc_output.space.count_f[2]$_SDFF_PP1_  (.D(_01729_),
    .CK(clknet_leaf_156_clk),
    .Q(\dynamic_node_top.proc_output.space.count_f[2] ),
    .QN(_00060_));
 DFF_X1 \dynamic_node_top.proc_output.space.is_one_f$_SDFF_PP0_  (.D(_01730_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.proc_output.space.is_one_f ),
    .QN(_08532_));
 DFF_X1 \dynamic_node_top.proc_output.space.is_two_or_more_f$_SDFF_PP1_  (.D(_01731_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.proc_output.space.is_two_or_more_f ),
    .QN(_08531_));
 DFF_X1 \dynamic_node_top.proc_output.space.valid_f$_SDFF_PP0_  (.D(_01732_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.proc_output.space.valid_f ),
    .QN(_10520_));
 DFF_X1 \dynamic_node_top.proc_output.space.yummy_f$_SDFF_PP0_  (.D(_01733_),
    .CK(clknet_leaf_155_clk),
    .Q(\dynamic_node_top.proc_output.space.yummy_f ),
    .QN(_10517_));
 DFF_X1 \dynamic_node_top.south_input.NIB.elements_in_array_f[0]$_SDFFE_PP0N_  (.D(_01734_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.south_input.NIB.elements_in_array_f[0] ),
    .QN(\dynamic_node_top.south_input.NIB.elements_in_array_next[0] ));
 DFF_X1 \dynamic_node_top.south_input.NIB.elements_in_array_f[1]$_SDFFE_PP0N_  (.D(_01735_),
    .CK(clknet_leaf_143_clk),
    .Q(\dynamic_node_top.south_input.NIB.elements_in_array_f[1] ),
    .QN(_08530_));
 DFF_X1 \dynamic_node_top.south_input.NIB.elements_in_array_f[2]$_SDFFE_PP0N_  (.D(_01736_),
    .CK(clknet_leaf_148_clk),
    .Q(\dynamic_node_top.south_input.NIB.elements_in_array_f[2] ),
    .QN(_08529_));
 DFF_X1 \dynamic_node_top.south_input.NIB.head_ptr_f[0]$_SDFFE_PP0N_  (.D(_01737_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.south_input.NIB.head_ptr_f[0] ),
    .QN(\dynamic_node_top.south_input.NIB.head_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.south_input.NIB.head_ptr_f[1]$_SDFFE_PP0N_  (.D(_00080_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.south_input.NIB.head_ptr_f[1] ),
    .QN(_08528_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][0]$_DFFE_PP_  (.D(_01738_),
    .CK(clknet_leaf_271_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][0] ),
    .QN(_08527_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][10]$_DFFE_PP_  (.D(_01739_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][10] ),
    .QN(_08526_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][11]$_DFFE_PP_  (.D(_01740_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][11] ),
    .QN(_08525_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][12]$_DFFE_PP_  (.D(_01741_),
    .CK(clknet_leaf_271_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][12] ),
    .QN(_08524_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][13]$_DFFE_PP_  (.D(_01742_),
    .CK(clknet_leaf_271_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][13] ),
    .QN(_08523_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][14]$_DFFE_PP_  (.D(_01743_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][14] ),
    .QN(_08522_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][15]$_DFFE_PP_  (.D(_01744_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][15] ),
    .QN(_08521_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][16]$_DFFE_PP_  (.D(_01745_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][16] ),
    .QN(_08520_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][17]$_DFFE_PP_  (.D(_01746_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][17] ),
    .QN(_08519_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][18]$_DFFE_PP_  (.D(_01747_),
    .CK(clknet_leaf_271_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][18] ),
    .QN(_08518_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][19]$_DFFE_PP_  (.D(_01748_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][19] ),
    .QN(_08517_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][1]$_DFFE_PP_  (.D(_01749_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][1] ),
    .QN(_08516_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][20]$_DFFE_PP_  (.D(_01750_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][20] ),
    .QN(_08515_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][21]$_DFFE_PP_  (.D(_01751_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][21] ),
    .QN(_08514_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][22]$_DFFE_PP_  (.D(_01752_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][22] ),
    .QN(_08513_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][23]$_DFFE_PP_  (.D(_01753_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][23] ),
    .QN(_08512_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][24]$_DFFE_PP_  (.D(_01754_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][24] ),
    .QN(_08511_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][25]$_DFFE_PP_  (.D(_01755_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][25] ),
    .QN(_08510_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][26]$_DFFE_PP_  (.D(_01756_),
    .CK(clknet_leaf_269_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][26] ),
    .QN(_08509_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][27]$_DFFE_PP_  (.D(_01757_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][27] ),
    .QN(_08508_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][28]$_DFFE_PP_  (.D(_01758_),
    .CK(clknet_leaf_249_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][28] ),
    .QN(_08507_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][29]$_DFFE_PP_  (.D(_01759_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][29] ),
    .QN(_08506_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][2]$_DFFE_PP_  (.D(_01760_),
    .CK(clknet_leaf_254_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][2] ),
    .QN(_08505_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][30]$_DFFE_PP_  (.D(_01761_),
    .CK(clknet_leaf_249_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][30] ),
    .QN(_08504_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][31]$_DFFE_PP_  (.D(_01762_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][31] ),
    .QN(_08503_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][32]$_DFFE_PP_  (.D(_01763_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][32] ),
    .QN(_08502_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][33]$_DFFE_PP_  (.D(_01764_),
    .CK(clknet_leaf_254_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][33] ),
    .QN(_08501_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][34]$_DFFE_PP_  (.D(_01765_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][34] ),
    .QN(_08500_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][35]$_DFFE_PP_  (.D(_01766_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][35] ),
    .QN(_08499_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][36]$_DFFE_PP_  (.D(_01767_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][36] ),
    .QN(_08498_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][37]$_DFFE_PP_  (.D(_01768_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][37] ),
    .QN(_08497_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][38]$_DFFE_PP_  (.D(_01769_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][38] ),
    .QN(_08496_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][39]$_DFFE_PP_  (.D(_01770_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][39] ),
    .QN(_08495_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][3]$_DFFE_PP_  (.D(_01771_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][3] ),
    .QN(_08494_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][40]$_DFFE_PP_  (.D(_01772_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][40] ),
    .QN(_08493_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][41]$_DFFE_PP_  (.D(_01773_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][41] ),
    .QN(_08492_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][42]$_DFFE_PP_  (.D(_01774_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][42] ),
    .QN(_08491_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][43]$_DFFE_PP_  (.D(_01775_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][43] ),
    .QN(_08490_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][44]$_DFFE_PP_  (.D(_01776_),
    .CK(clknet_leaf_262_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][44] ),
    .QN(_08489_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][45]$_DFFE_PP_  (.D(_01777_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][45] ),
    .QN(_08488_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][46]$_DFFE_PP_  (.D(_01778_),
    .CK(clknet_leaf_285_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][46] ),
    .QN(_08487_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][47]$_DFFE_PP_  (.D(_01779_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][47] ),
    .QN(_08486_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][48]$_DFFE_PP_  (.D(_01780_),
    .CK(clknet_leaf_285_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][48] ),
    .QN(_08485_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][49]$_DFFE_PP_  (.D(_01781_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][49] ),
    .QN(_08484_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][4]$_DFFE_PP_  (.D(_01782_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][4] ),
    .QN(_08483_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][50]$_DFFE_PP_  (.D(_01783_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][50] ),
    .QN(_08482_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][51]$_DFFE_PP_  (.D(_01784_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][51] ),
    .QN(_08481_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][52]$_DFFE_PP_  (.D(_01785_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][52] ),
    .QN(_08480_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][53]$_DFFE_PP_  (.D(_01786_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][53] ),
    .QN(_08479_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][54]$_DFFE_PP_  (.D(_01787_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][54] ),
    .QN(_08478_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][55]$_DFFE_PP_  (.D(_01788_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][55] ),
    .QN(_08477_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][56]$_DFFE_PP_  (.D(_01789_),
    .CK(clknet_leaf_294_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][56] ),
    .QN(_08476_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][57]$_DFFE_PP_  (.D(_01790_),
    .CK(clknet_leaf_293_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][57] ),
    .QN(_08475_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][58]$_DFFE_PP_  (.D(_01791_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][58] ),
    .QN(_08474_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][59]$_DFFE_PP_  (.D(_01792_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][59] ),
    .QN(_08473_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][5]$_DFFE_PP_  (.D(_01793_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][5] ),
    .QN(_08472_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][60]$_DFFE_PP_  (.D(_01794_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][60] ),
    .QN(_08471_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][61]$_DFFE_PP_  (.D(_01795_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][61] ),
    .QN(_08470_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][62]$_DFFE_PP_  (.D(_01796_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][62] ),
    .QN(_08469_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][63]$_DFFE_PP_  (.D(_01797_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][63] ),
    .QN(_08468_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][6]$_DFFE_PP_  (.D(_01798_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][6] ),
    .QN(_08467_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][7]$_DFFE_PP_  (.D(_01799_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][7] ),
    .QN(_08466_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][8]$_DFFE_PP_  (.D(_01800_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][8] ),
    .QN(_08465_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[0][9]$_DFFE_PP_  (.D(_01801_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[0][9] ),
    .QN(_08464_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][0]$_DFFE_PP_  (.D(_01802_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][0] ),
    .QN(_08463_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][10]$_DFFE_PP_  (.D(_01803_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][10] ),
    .QN(_08462_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][11]$_DFFE_PP_  (.D(_01804_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][11] ),
    .QN(_08461_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][12]$_DFFE_PP_  (.D(_01805_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][12] ),
    .QN(_08460_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][13]$_DFFE_PP_  (.D(_01806_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][13] ),
    .QN(_08459_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][14]$_DFFE_PP_  (.D(_01807_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][14] ),
    .QN(_08458_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][15]$_DFFE_PP_  (.D(_01808_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][15] ),
    .QN(_08457_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][16]$_DFFE_PP_  (.D(_01809_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][16] ),
    .QN(_08456_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][17]$_DFFE_PP_  (.D(_01810_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][17] ),
    .QN(_08455_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][18]$_DFFE_PP_  (.D(_01811_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][18] ),
    .QN(_08454_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][19]$_DFFE_PP_  (.D(_01812_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][19] ),
    .QN(_08453_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][1]$_DFFE_PP_  (.D(_01813_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][1] ),
    .QN(_08452_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][20]$_DFFE_PP_  (.D(_01814_),
    .CK(clknet_leaf_269_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][20] ),
    .QN(_08451_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][21]$_DFFE_PP_  (.D(_01815_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][21] ),
    .QN(_08450_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][22]$_DFFE_PP_  (.D(_01816_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][22] ),
    .QN(_08449_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][23]$_DFFE_PP_  (.D(_01817_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][23] ),
    .QN(_08448_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][24]$_DFFE_PP_  (.D(_01818_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][24] ),
    .QN(_08447_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][25]$_DFFE_PP_  (.D(_01819_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][25] ),
    .QN(_08446_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][26]$_DFFE_PP_  (.D(_01820_),
    .CK(clknet_leaf_269_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][26] ),
    .QN(_08445_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][27]$_DFFE_PP_  (.D(_01821_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][27] ),
    .QN(_08444_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][28]$_DFFE_PP_  (.D(_01822_),
    .CK(clknet_leaf_249_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][28] ),
    .QN(_08443_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][29]$_DFFE_PP_  (.D(_01823_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][29] ),
    .QN(_08442_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][2]$_DFFE_PP_  (.D(_01824_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][2] ),
    .QN(_08441_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][30]$_DFFE_PP_  (.D(_01825_),
    .CK(clknet_leaf_249_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][30] ),
    .QN(_08440_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][31]$_DFFE_PP_  (.D(_01826_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][31] ),
    .QN(_08439_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][32]$_DFFE_PP_  (.D(_01827_),
    .CK(clknet_leaf_254_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][32] ),
    .QN(_08438_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][33]$_DFFE_PP_  (.D(_01828_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][33] ),
    .QN(_08437_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][34]$_DFFE_PP_  (.D(_01829_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][34] ),
    .QN(_08436_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][35]$_DFFE_PP_  (.D(_01830_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][35] ),
    .QN(_08435_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][36]$_DFFE_PP_  (.D(_01831_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][36] ),
    .QN(_08434_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][37]$_DFFE_PP_  (.D(_01832_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][37] ),
    .QN(_08433_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][38]$_DFFE_PP_  (.D(_01833_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][38] ),
    .QN(_08432_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][39]$_DFFE_PP_  (.D(_01834_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][39] ),
    .QN(_08431_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][3]$_DFFE_PP_  (.D(_01835_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][3] ),
    .QN(_08430_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][40]$_DFFE_PP_  (.D(_01836_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][40] ),
    .QN(_08429_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][41]$_DFFE_PP_  (.D(_01837_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][41] ),
    .QN(_08428_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][42]$_DFFE_PP_  (.D(_01838_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][42] ),
    .QN(_08427_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][43]$_DFFE_PP_  (.D(_01839_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][43] ),
    .QN(_08426_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][44]$_DFFE_PP_  (.D(_01840_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][44] ),
    .QN(_08425_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][45]$_DFFE_PP_  (.D(_01841_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][45] ),
    .QN(_08424_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][46]$_DFFE_PP_  (.D(_01842_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][46] ),
    .QN(_08423_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][47]$_DFFE_PP_  (.D(_01843_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][47] ),
    .QN(_08422_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][48]$_DFFE_PP_  (.D(_01844_),
    .CK(clknet_leaf_285_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][48] ),
    .QN(_08421_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][49]$_DFFE_PP_  (.D(_01845_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][49] ),
    .QN(_08420_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][4]$_DFFE_PP_  (.D(_01846_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][4] ),
    .QN(_08419_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][50]$_DFFE_PP_  (.D(_01847_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][50] ),
    .QN(_08418_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][51]$_DFFE_PP_  (.D(_01848_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][51] ),
    .QN(_08417_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][52]$_DFFE_PP_  (.D(_01849_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][52] ),
    .QN(_08416_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][53]$_DFFE_PP_  (.D(_01850_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][53] ),
    .QN(_08415_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][54]$_DFFE_PP_  (.D(_01851_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][54] ),
    .QN(_08414_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][55]$_DFFE_PP_  (.D(_01852_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][55] ),
    .QN(_08413_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][56]$_DFFE_PP_  (.D(_01853_),
    .CK(clknet_leaf_294_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][56] ),
    .QN(_08412_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][57]$_DFFE_PP_  (.D(_01854_),
    .CK(clknet_leaf_294_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][57] ),
    .QN(_08411_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][58]$_DFFE_PP_  (.D(_01855_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][58] ),
    .QN(_08410_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][59]$_DFFE_PP_  (.D(_01856_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][59] ),
    .QN(_08409_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][5]$_DFFE_PP_  (.D(_01857_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][5] ),
    .QN(_08408_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][60]$_DFFE_PP_  (.D(_01858_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][60] ),
    .QN(_08407_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][61]$_DFFE_PP_  (.D(_01859_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][61] ),
    .QN(_08406_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][62]$_DFFE_PP_  (.D(_01860_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][62] ),
    .QN(_08405_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][63]$_DFFE_PP_  (.D(_01861_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][63] ),
    .QN(_08404_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][6]$_DFFE_PP_  (.D(_01862_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][6] ),
    .QN(_08403_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][7]$_DFFE_PP_  (.D(_01863_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][7] ),
    .QN(_08402_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][8]$_DFFE_PP_  (.D(_01864_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][8] ),
    .QN(_08401_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[1][9]$_DFFE_PP_  (.D(_01865_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[1][9] ),
    .QN(_08400_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][0]$_DFFE_PP_  (.D(_01866_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][0] ),
    .QN(_08399_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][10]$_DFFE_PP_  (.D(_01867_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][10] ),
    .QN(_08398_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][11]$_DFFE_PP_  (.D(_01868_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][11] ),
    .QN(_08397_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][12]$_DFFE_PP_  (.D(_01869_),
    .CK(clknet_leaf_271_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][12] ),
    .QN(_08396_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][13]$_DFFE_PP_  (.D(_01870_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][13] ),
    .QN(_08395_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][14]$_DFFE_PP_  (.D(_01871_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][14] ),
    .QN(_08394_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][15]$_DFFE_PP_  (.D(_01872_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][15] ),
    .QN(_08393_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][16]$_DFFE_PP_  (.D(_01873_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][16] ),
    .QN(_08392_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][17]$_DFFE_PP_  (.D(_01874_),
    .CK(clknet_leaf_272_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][17] ),
    .QN(_08391_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][18]$_DFFE_PP_  (.D(_01875_),
    .CK(clknet_leaf_271_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][18] ),
    .QN(_08390_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][19]$_DFFE_PP_  (.D(_01876_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][19] ),
    .QN(_08389_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][1]$_DFFE_PP_  (.D(_01877_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][1] ),
    .QN(_08388_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][20]$_DFFE_PP_  (.D(_01878_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][20] ),
    .QN(_08387_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][21]$_DFFE_PP_  (.D(_01879_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][21] ),
    .QN(_08386_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][22]$_DFFE_PP_  (.D(_01880_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][22] ),
    .QN(_08385_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][23]$_DFFE_PP_  (.D(_01881_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][23] ),
    .QN(_08384_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][24]$_DFFE_PP_  (.D(_01882_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][24] ),
    .QN(_08383_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][25]$_DFFE_PP_  (.D(_01883_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][25] ),
    .QN(_08382_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][26]$_DFFE_PP_  (.D(_01884_),
    .CK(clknet_leaf_269_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][26] ),
    .QN(_08381_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][27]$_DFFE_PP_  (.D(_01885_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][27] ),
    .QN(_08380_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][28]$_DFFE_PP_  (.D(_01886_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][28] ),
    .QN(_08379_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][29]$_DFFE_PP_  (.D(_01887_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][29] ),
    .QN(_08378_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][2]$_DFFE_PP_  (.D(_01888_),
    .CK(clknet_leaf_254_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][2] ),
    .QN(_08377_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][30]$_DFFE_PP_  (.D(_01889_),
    .CK(clknet_leaf_249_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][30] ),
    .QN(_08376_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][31]$_DFFE_PP_  (.D(_01890_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][31] ),
    .QN(_08375_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][32]$_DFFE_PP_  (.D(_01891_),
    .CK(clknet_leaf_254_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][32] ),
    .QN(_08374_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][33]$_DFFE_PP_  (.D(_01892_),
    .CK(clknet_leaf_254_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][33] ),
    .QN(_08373_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][34]$_DFFE_PP_  (.D(_01893_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][34] ),
    .QN(_08372_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][35]$_DFFE_PP_  (.D(_01894_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][35] ),
    .QN(_08371_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][36]$_DFFE_PP_  (.D(_01895_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][36] ),
    .QN(_08370_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][37]$_DFFE_PP_  (.D(_01896_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][37] ),
    .QN(_08369_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][38]$_DFFE_PP_  (.D(_01897_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][38] ),
    .QN(_08368_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][39]$_DFFE_PP_  (.D(_01898_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][39] ),
    .QN(_08367_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][3]$_DFFE_PP_  (.D(_01899_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][3] ),
    .QN(_08366_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][40]$_DFFE_PP_  (.D(_01900_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][40] ),
    .QN(_08365_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][41]$_DFFE_PP_  (.D(_01901_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][41] ),
    .QN(_08364_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][42]$_DFFE_PP_  (.D(_01902_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][42] ),
    .QN(_08363_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][43]$_DFFE_PP_  (.D(_01903_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][43] ),
    .QN(_08362_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][44]$_DFFE_PP_  (.D(_01904_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][44] ),
    .QN(_08361_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][45]$_DFFE_PP_  (.D(_01905_),
    .CK(clknet_leaf_258_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][45] ),
    .QN(_08360_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][46]$_DFFE_PP_  (.D(_01906_),
    .CK(clknet_leaf_285_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][46] ),
    .QN(_08359_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][47]$_DFFE_PP_  (.D(_01907_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][47] ),
    .QN(_08358_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][48]$_DFFE_PP_  (.D(_01908_),
    .CK(clknet_leaf_285_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][48] ),
    .QN(_08357_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][49]$_DFFE_PP_  (.D(_01909_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][49] ),
    .QN(_08356_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][4]$_DFFE_PP_  (.D(_01910_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][4] ),
    .QN(_08355_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][50]$_DFFE_PP_  (.D(_01911_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][50] ),
    .QN(_08354_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][51]$_DFFE_PP_  (.D(_01912_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][51] ),
    .QN(_08353_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][52]$_DFFE_PP_  (.D(_01913_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][52] ),
    .QN(_08352_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][53]$_DFFE_PP_  (.D(_01914_),
    .CK(clknet_leaf_284_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][53] ),
    .QN(_08351_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][54]$_DFFE_PP_  (.D(_01915_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][54] ),
    .QN(_08350_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][55]$_DFFE_PP_  (.D(_01916_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][55] ),
    .QN(_08349_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][56]$_DFFE_PP_  (.D(_01917_),
    .CK(clknet_leaf_294_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][56] ),
    .QN(_08348_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][57]$_DFFE_PP_  (.D(_01918_),
    .CK(clknet_leaf_293_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][57] ),
    .QN(_08347_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][58]$_DFFE_PP_  (.D(_01919_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][58] ),
    .QN(_08346_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][59]$_DFFE_PP_  (.D(_01920_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][59] ),
    .QN(_08345_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][5]$_DFFE_PP_  (.D(_01921_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][5] ),
    .QN(_08344_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][60]$_DFFE_PP_  (.D(_01922_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][60] ),
    .QN(_08343_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][61]$_DFFE_PP_  (.D(_01923_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][61] ),
    .QN(_08342_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][62]$_DFFE_PP_  (.D(_01924_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][62] ),
    .QN(_08341_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][63]$_DFFE_PP_  (.D(_01925_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][63] ),
    .QN(_08340_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][6]$_DFFE_PP_  (.D(_01926_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][6] ),
    .QN(_08339_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][7]$_DFFE_PP_  (.D(_01927_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][7] ),
    .QN(_08338_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][8]$_DFFE_PP_  (.D(_01928_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][8] ),
    .QN(_08337_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[2][9]$_DFFE_PP_  (.D(_01929_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[2][9] ),
    .QN(_08336_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][0]$_DFFE_PP_  (.D(_01930_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][0] ),
    .QN(_08335_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][10]$_DFFE_PP_  (.D(_01931_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][10] ),
    .QN(_08334_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][11]$_DFFE_PP_  (.D(_01932_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][11] ),
    .QN(_08333_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][12]$_DFFE_PP_  (.D(_01933_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][12] ),
    .QN(_08332_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][13]$_DFFE_PP_  (.D(_01934_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][13] ),
    .QN(_08331_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][14]$_DFFE_PP_  (.D(_01935_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][14] ),
    .QN(_08330_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][15]$_DFFE_PP_  (.D(_01936_),
    .CK(clknet_leaf_276_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][15] ),
    .QN(_08329_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][16]$_DFFE_PP_  (.D(_01937_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][16] ),
    .QN(_08328_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][17]$_DFFE_PP_  (.D(_01938_),
    .CK(clknet_leaf_274_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][17] ),
    .QN(_08327_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][18]$_DFFE_PP_  (.D(_01939_),
    .CK(clknet_leaf_275_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][18] ),
    .QN(_08326_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][19]$_DFFE_PP_  (.D(_01940_),
    .CK(clknet_leaf_269_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][19] ),
    .QN(_08325_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][1]$_DFFE_PP_  (.D(_01941_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][1] ),
    .QN(_08324_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][20]$_DFFE_PP_  (.D(_01942_),
    .CK(clknet_leaf_269_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][20] ),
    .QN(_08323_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][21]$_DFFE_PP_  (.D(_01943_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][21] ),
    .QN(_08322_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][22]$_DFFE_PP_  (.D(_01944_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][22] ),
    .QN(_08321_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][23]$_DFFE_PP_  (.D(_01945_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][23] ),
    .QN(_08320_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][24]$_DFFE_PP_  (.D(_01946_),
    .CK(clknet_leaf_251_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][24] ),
    .QN(_08319_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][25]$_DFFE_PP_  (.D(_01947_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][25] ),
    .QN(_08318_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][26]$_DFFE_PP_  (.D(_01948_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][26] ),
    .QN(_08317_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][27]$_DFFE_PP_  (.D(_01949_),
    .CK(clknet_leaf_247_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][27] ),
    .QN(_08316_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][28]$_DFFE_PP_  (.D(_01950_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][28] ),
    .QN(_08315_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][29]$_DFFE_PP_  (.D(_01951_),
    .CK(clknet_leaf_250_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][29] ),
    .QN(_08314_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][2]$_DFFE_PP_  (.D(_01952_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][2] ),
    .QN(_08313_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][30]$_DFFE_PP_  (.D(_01953_),
    .CK(clknet_leaf_249_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][30] ),
    .QN(_08312_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][31]$_DFFE_PP_  (.D(_01954_),
    .CK(clknet_leaf_248_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][31] ),
    .QN(_08311_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][32]$_DFFE_PP_  (.D(_01955_),
    .CK(clknet_leaf_252_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][32] ),
    .QN(_08310_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][33]$_DFFE_PP_  (.D(_01956_),
    .CK(clknet_leaf_253_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][33] ),
    .QN(_08309_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][34]$_DFFE_PP_  (.D(_01957_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][34] ),
    .QN(_08308_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][35]$_DFFE_PP_  (.D(_01958_),
    .CK(clknet_leaf_257_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][35] ),
    .QN(_08307_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][36]$_DFFE_PP_  (.D(_01959_),
    .CK(clknet_leaf_256_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][36] ),
    .QN(_08306_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][37]$_DFFE_PP_  (.D(_01960_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][37] ),
    .QN(_08305_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][38]$_DFFE_PP_  (.D(_01961_),
    .CK(clknet_leaf_255_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][38] ),
    .QN(_08304_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][39]$_DFFE_PP_  (.D(_01962_),
    .CK(clknet_leaf_264_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][39] ),
    .QN(_08303_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][3]$_DFFE_PP_  (.D(_01963_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][3] ),
    .QN(_08302_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][40]$_DFFE_PP_  (.D(_01964_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][40] ),
    .QN(_08301_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][41]$_DFFE_PP_  (.D(_01965_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][41] ),
    .QN(_08300_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][42]$_DFFE_PP_  (.D(_01966_),
    .CK(clknet_leaf_266_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][42] ),
    .QN(_08299_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][43]$_DFFE_PP_  (.D(_01967_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][43] ),
    .QN(_08298_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][44]$_DFFE_PP_  (.D(_01968_),
    .CK(clknet_leaf_263_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][44] ),
    .QN(_08297_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][45]$_DFFE_PP_  (.D(_01969_),
    .CK(clknet_leaf_259_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][45] ),
    .QN(_08296_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][46]$_DFFE_PP_  (.D(_01970_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][46] ),
    .QN(_08295_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][47]$_DFFE_PP_  (.D(_01971_),
    .CK(clknet_leaf_265_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][47] ),
    .QN(_08294_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][48]$_DFFE_PP_  (.D(_01972_),
    .CK(clknet_leaf_286_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][48] ),
    .QN(_08293_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][49]$_DFFE_PP_  (.D(_01973_),
    .CK(clknet_leaf_278_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][49] ),
    .QN(_08292_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][4]$_DFFE_PP_  (.D(_01974_),
    .CK(clknet_leaf_273_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][4] ),
    .QN(_08291_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][50]$_DFFE_PP_  (.D(_01975_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][50] ),
    .QN(_08290_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][51]$_DFFE_PP_  (.D(_01976_),
    .CK(clknet_leaf_285_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][51] ),
    .QN(_08289_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][52]$_DFFE_PP_  (.D(_01977_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][52] ),
    .QN(_08288_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][53]$_DFFE_PP_  (.D(_01978_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][53] ),
    .QN(_08287_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][54]$_DFFE_PP_  (.D(_01979_),
    .CK(clknet_leaf_283_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][54] ),
    .QN(_08286_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][55]$_DFFE_PP_  (.D(_01980_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][55] ),
    .QN(_08285_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][56]$_DFFE_PP_  (.D(_01981_),
    .CK(clknet_leaf_294_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][56] ),
    .QN(_08284_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][57]$_DFFE_PP_  (.D(_01982_),
    .CK(clknet_leaf_294_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][57] ),
    .QN(_08283_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][58]$_DFFE_PP_  (.D(_01983_),
    .CK(clknet_leaf_281_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][58] ),
    .QN(_08282_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][59]$_DFFE_PP_  (.D(_01984_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][59] ),
    .QN(_08281_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][5]$_DFFE_PP_  (.D(_01985_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][5] ),
    .QN(_08280_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][60]$_DFFE_PP_  (.D(_01986_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][60] ),
    .QN(_08279_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][61]$_DFFE_PP_  (.D(_01987_),
    .CK(clknet_leaf_279_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][61] ),
    .QN(_08278_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][62]$_DFFE_PP_  (.D(_01988_),
    .CK(clknet_leaf_282_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][62] ),
    .QN(_08277_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][63]$_DFFE_PP_  (.D(_01989_),
    .CK(clknet_leaf_280_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][63] ),
    .QN(_08276_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][6]$_DFFE_PP_  (.D(_01990_),
    .CK(clknet_leaf_270_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][6] ),
    .QN(_08275_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][7]$_DFFE_PP_  (.D(_01991_),
    .CK(clknet_leaf_267_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][7] ),
    .QN(_08274_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][8]$_DFFE_PP_  (.D(_01992_),
    .CK(clknet_leaf_277_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][8] ),
    .QN(_08273_));
 DFF_X1 \dynamic_node_top.south_input.NIB.storage_data_f[3][9]$_DFFE_PP_  (.D(_01993_),
    .CK(clknet_leaf_268_clk),
    .Q(\dynamic_node_top.south_input.NIB.storage_data_f[3][9] ),
    .QN(_08272_));
 DFF_X1 \dynamic_node_top.south_input.NIB.tail_ptr_f[0]$_SDFFE_PP0N_  (.D(_01994_),
    .CK(clknet_leaf_292_clk),
    .Q(\dynamic_node_top.south_input.NIB.tail_ptr_f[0] ),
    .QN(\dynamic_node_top.south_input.NIB.tail_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.south_input.NIB.tail_ptr_f[1]$_SDFFE_PP0N_  (.D(_01995_),
    .CK(clknet_leaf_293_clk),
    .Q(\dynamic_node_top.south_input.NIB.tail_ptr_f[1] ),
    .QN(_10601_));
 DFF_X1 \dynamic_node_top.south_input.NIB.yummy_out_f$_SDFF_PP0_  (.D(_01996_),
    .CK(clknet_leaf_154_clk),
    .Q(net629),
    .QN(_08271_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[0]$_SDFF_PP0_  (.D(_01997_),
    .CK(clknet_leaf_142_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[0] ),
    .QN(_10513_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[1]$_SDFF_PP0_  (.D(_01998_),
    .CK(clknet_leaf_142_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[1] ),
    .QN(_10514_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[2]$_SDFF_PP0_  (.D(_01999_),
    .CK(clknet_leaf_140_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[2] ),
    .QN(_08270_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[3]$_SDFF_PP0_  (.D(_02000_),
    .CK(clknet_leaf_140_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[3] ),
    .QN(_08269_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[4]$_SDFF_PP0_  (.D(_02001_),
    .CK(clknet_leaf_140_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[4] ),
    .QN(_08268_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[5]$_SDFF_PP0_  (.D(_02002_),
    .CK(clknet_leaf_141_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[5] ),
    .QN(_08267_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[6]$_SDFF_PP0_  (.D(_02003_),
    .CK(clknet_leaf_141_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[6] ),
    .QN(_08266_));
 DFF_X1 \dynamic_node_top.south_input.control.count_f[7]$_SDFF_PP0_  (.D(_02004_),
    .CK(clknet_leaf_141_clk),
    .Q(\dynamic_node_top.south_input.control.count_f[7] ),
    .QN(_08265_));
 DFF_X1 \dynamic_node_top.south_input.control.count_one_f$_SDFF_PP0_  (.D(_02005_),
    .CK(clknet_leaf_158_clk),
    .Q(\dynamic_node_top.south_input.control.count_one_f ),
    .QN(_10158_));
 DFF_X1 \dynamic_node_top.south_input.control.header_temp$_DFF_P_  (.D(_00003_),
    .CK(clknet_leaf_142_clk),
    .Q(\dynamic_node_top.south_input.control.header_last_temp ),
    .QN(_08264_));
 DFF_X1 \dynamic_node_top.south_input.control.tail_last_f$_SDFF_PP0_  (.D(_02006_),
    .CK(clknet_leaf_158_clk),
    .Q(\dynamic_node_top.south_input.control.tail_last_f ),
    .QN(_10159_));
 DFF_X1 \dynamic_node_top.south_output.control.current_route_f[0]$_DFF_P_  (.D(_00027_),
    .CK(clknet_leaf_157_clk),
    .Q(\dynamic_node_top.south_output.control.current_route_f[0] ),
    .QN(_00048_));
 DFF_X1 \dynamic_node_top.south_output.control.current_route_f[1]$_DFF_P_  (.D(_00028_),
    .CK(clknet_leaf_157_clk),
    .Q(\dynamic_node_top.south_output.control.current_route_f[1] ),
    .QN(_00047_));
 DFF_X1 \dynamic_node_top.south_output.control.current_route_f[2]$_DFF_P_  (.D(_00029_),
    .CK(clknet_leaf_160_clk),
    .Q(\dynamic_node_top.south_output.control.current_route_f[2] ),
    .QN(_00069_));
 DFF_X1 \dynamic_node_top.south_output.control.current_route_f[3]$_DFF_P_  (.D(_00030_),
    .CK(clknet_leaf_160_clk),
    .Q(\dynamic_node_top.south_output.control.current_route_f[3] ),
    .QN(_00070_));
 DFF_X1 \dynamic_node_top.south_output.control.current_route_f[4]$_DFF_P_  (.D(_00031_),
    .CK(clknet_leaf_162_clk),
    .Q(\dynamic_node_top.south_output.control.current_route_f[4] ),
    .QN(_00068_));
 DFF_X1 \dynamic_node_top.south_output.control.planned_f$_SDFF_PP0_  (.D(_02007_),
    .CK(clknet_leaf_163_clk),
    .Q(\dynamic_node_top.south_output.control.planned_f ),
    .QN(_00049_));
 DFF_X2 \dynamic_node_top.south_output.space.count_f[0]$_SDFF_PP0_  (.D(_02008_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.south_output.space.count_f[0] ),
    .QN(_10489_));
 DFF_X2 \dynamic_node_top.south_output.space.count_f[1]$_SDFF_PP0_  (.D(_02009_),
    .CK(clknet_leaf_166_clk),
    .Q(\dynamic_node_top.south_output.space.count_f[1] ),
    .QN(_10490_));
 DFF_X1 \dynamic_node_top.south_output.space.count_f[2]$_SDFF_PP1_  (.D(_02010_),
    .CK(clknet_leaf_166_clk),
    .Q(\dynamic_node_top.south_output.space.count_f[2] ),
    .QN(_00059_));
 DFF_X1 \dynamic_node_top.south_output.space.is_one_f$_SDFF_PP0_  (.D(_02011_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.south_output.space.is_one_f ),
    .QN(_08263_));
 DFF_X1 \dynamic_node_top.south_output.space.is_two_or_more_f$_SDFF_PP1_  (.D(_02012_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.south_output.space.is_two_or_more_f ),
    .QN(_08262_));
 DFF_X1 \dynamic_node_top.south_output.space.valid_f$_SDFF_PP0_  (.D(_02013_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.south_output.space.valid_f ),
    .QN(_10486_));
 DFF_X1 \dynamic_node_top.south_output.space.yummy_f$_SDFF_PP0_  (.D(_02014_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.south_output.space.yummy_f ),
    .QN(_10483_));
 DFF_X1 \dynamic_node_top.west_input.NIB.elements_in_array_f[0]$_SDFFE_PP0N_  (.D(_02015_),
    .CK(clknet_leaf_167_clk),
    .Q(\dynamic_node_top.west_input.NIB.elements_in_array_f[0] ),
    .QN(\dynamic_node_top.west_input.NIB.elements_in_array_next[0] ));
 DFF_X1 \dynamic_node_top.west_input.NIB.elements_in_array_f[1]$_SDFFE_PP0N_  (.D(_02016_),
    .CK(clknet_leaf_167_clk),
    .Q(\dynamic_node_top.west_input.NIB.elements_in_array_f[1] ),
    .QN(_08261_));
 DFF_X1 \dynamic_node_top.west_input.NIB.elements_in_array_f[2]$_SDFFE_PP0N_  (.D(_02017_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.west_input.NIB.elements_in_array_f[2] ),
    .QN(_08260_));
 DFF_X1 \dynamic_node_top.west_input.NIB.head_ptr_f[0]$_SDFFE_PP0N_  (.D(_02018_),
    .CK(clknet_leaf_167_clk),
    .Q(\dynamic_node_top.west_input.NIB.head_ptr_f[0] ),
    .QN(\dynamic_node_top.west_input.NIB.head_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.west_input.NIB.head_ptr_f[1]$_SDFFE_PP0N_  (.D(_00078_),
    .CK(clknet_leaf_175_clk),
    .Q(\dynamic_node_top.west_input.NIB.head_ptr_f[1] ),
    .QN(_08259_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][0]$_DFFE_PP_  (.D(_02019_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][0] ),
    .QN(_08258_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][10]$_DFFE_PP_  (.D(_02020_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][10] ),
    .QN(_08257_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][11]$_DFFE_PP_  (.D(_02021_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][11] ),
    .QN(_08256_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][12]$_DFFE_PP_  (.D(_02022_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][12] ),
    .QN(_08255_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][13]$_DFFE_PP_  (.D(_02023_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][13] ),
    .QN(_08254_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][14]$_DFFE_PP_  (.D(_02024_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][14] ),
    .QN(_08253_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][15]$_DFFE_PP_  (.D(_02025_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][15] ),
    .QN(_08252_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][16]$_DFFE_PP_  (.D(_02026_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][16] ),
    .QN(_08251_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][17]$_DFFE_PP_  (.D(_02027_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][17] ),
    .QN(_08250_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][18]$_DFFE_PP_  (.D(_02028_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][18] ),
    .QN(_08249_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][19]$_DFFE_PP_  (.D(_02029_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][19] ),
    .QN(_08248_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][1]$_DFFE_PP_  (.D(_02030_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][1] ),
    .QN(_08247_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][20]$_DFFE_PP_  (.D(_02031_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][20] ),
    .QN(_08246_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][21]$_DFFE_PP_  (.D(_02032_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][21] ),
    .QN(_08245_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][22]$_DFFE_PP_  (.D(_02033_),
    .CK(clknet_leaf_166_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][22] ),
    .QN(_08244_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][23]$_DFFE_PP_  (.D(_02034_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][23] ),
    .QN(_08243_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][24]$_DFFE_PP_  (.D(_02035_),
    .CK(clknet_leaf_166_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][24] ),
    .QN(_08242_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][25]$_DFFE_PP_  (.D(_02036_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][25] ),
    .QN(_08241_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][26]$_DFFE_PP_  (.D(_02037_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][26] ),
    .QN(_08240_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][27]$_DFFE_PP_  (.D(_02038_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][27] ),
    .QN(_08239_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][28]$_DFFE_PP_  (.D(_02039_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][28] ),
    .QN(_08238_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][29]$_DFFE_PP_  (.D(_02040_),
    .CK(clknet_leaf_171_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][29] ),
    .QN(_08237_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][2]$_DFFE_PP_  (.D(_02041_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][2] ),
    .QN(_08236_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][30]$_DFFE_PP_  (.D(_02042_),
    .CK(clknet_leaf_171_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][30] ),
    .QN(_08235_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][31]$_DFFE_PP_  (.D(_02043_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][31] ),
    .QN(_08234_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][32]$_DFFE_PP_  (.D(_02044_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][32] ),
    .QN(_08233_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][33]$_DFFE_PP_  (.D(_02045_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][33] ),
    .QN(_08232_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][34]$_DFFE_PP_  (.D(_02046_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][34] ),
    .QN(_08231_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][35]$_DFFE_PP_  (.D(_02047_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][35] ),
    .QN(_08230_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][36]$_DFFE_PP_  (.D(_02048_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][36] ),
    .QN(_08229_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][37]$_DFFE_PP_  (.D(_02049_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][37] ),
    .QN(_08228_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][38]$_DFFE_PP_  (.D(_02050_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][38] ),
    .QN(_08227_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][39]$_DFFE_PP_  (.D(_02051_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][39] ),
    .QN(_08226_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][3]$_DFFE_PP_  (.D(_02052_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][3] ),
    .QN(_08225_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][40]$_DFFE_PP_  (.D(_02053_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][40] ),
    .QN(_08224_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][41]$_DFFE_PP_  (.D(_02054_),
    .CK(clknet_leaf_185_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][41] ),
    .QN(_08223_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][42]$_DFFE_PP_  (.D(_02055_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][42] ),
    .QN(_08222_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][43]$_DFFE_PP_  (.D(_02056_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][43] ),
    .QN(_08221_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][44]$_DFFE_PP_  (.D(_02057_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][44] ),
    .QN(_08220_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][45]$_DFFE_PP_  (.D(_02058_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][45] ),
    .QN(_08219_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][46]$_DFFE_PP_  (.D(_02059_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][46] ),
    .QN(_08218_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][47]$_DFFE_PP_  (.D(_02060_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][47] ),
    .QN(_08217_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][48]$_DFFE_PP_  (.D(_02061_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][48] ),
    .QN(_08216_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][49]$_DFFE_PP_  (.D(_02062_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][49] ),
    .QN(_08215_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][4]$_DFFE_PP_  (.D(_02063_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][4] ),
    .QN(_08214_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][50]$_DFFE_PP_  (.D(_02064_),
    .CK(clknet_leaf_193_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][50] ),
    .QN(_08213_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][51]$_DFFE_PP_  (.D(_02065_),
    .CK(clknet_leaf_196_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][51] ),
    .QN(_08212_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][52]$_DFFE_PP_  (.D(_02066_),
    .CK(clknet_leaf_193_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][52] ),
    .QN(_08211_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][53]$_DFFE_PP_  (.D(_02067_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][53] ),
    .QN(_08210_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][54]$_DFFE_PP_  (.D(_02068_),
    .CK(clknet_leaf_195_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][54] ),
    .QN(_08209_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][55]$_DFFE_PP_  (.D(_02069_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][55] ),
    .QN(_08208_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][56]$_DFFE_PP_  (.D(_02070_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][56] ),
    .QN(_08207_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][57]$_DFFE_PP_  (.D(_02071_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][57] ),
    .QN(_08206_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][58]$_DFFE_PP_  (.D(_02072_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][58] ),
    .QN(_08205_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][59]$_DFFE_PP_  (.D(_02073_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][59] ),
    .QN(_08204_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][5]$_DFFE_PP_  (.D(_02074_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][5] ),
    .QN(_08203_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][60]$_DFFE_PP_  (.D(_02075_),
    .CK(clknet_leaf_190_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][60] ),
    .QN(_08202_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][61]$_DFFE_PP_  (.D(_02076_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][61] ),
    .QN(_08201_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][62]$_DFFE_PP_  (.D(_02077_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][62] ),
    .QN(_08200_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][63]$_DFFE_PP_  (.D(_02078_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][63] ),
    .QN(_08199_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][6]$_DFFE_PP_  (.D(_02079_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][6] ),
    .QN(_08198_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][7]$_DFFE_PP_  (.D(_02080_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][7] ),
    .QN(_08197_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][8]$_DFFE_PP_  (.D(_02081_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][8] ),
    .QN(_08196_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[0][9]$_DFFE_PP_  (.D(_02082_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[0][9] ),
    .QN(_08195_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][0]$_DFFE_PP_  (.D(_02083_),
    .CK(clknet_leaf_221_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][0] ),
    .QN(_08194_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][10]$_DFFE_PP_  (.D(_02084_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][10] ),
    .QN(_08193_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][11]$_DFFE_PP_  (.D(_02085_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][11] ),
    .QN(_08192_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][12]$_DFFE_PP_  (.D(_02086_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][12] ),
    .QN(_08191_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][13]$_DFFE_PP_  (.D(_02087_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][13] ),
    .QN(_08190_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][14]$_DFFE_PP_  (.D(_02088_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][14] ),
    .QN(_08189_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][15]$_DFFE_PP_  (.D(_02089_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][15] ),
    .QN(_08188_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][16]$_DFFE_PP_  (.D(_02090_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][16] ),
    .QN(_08187_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][17]$_DFFE_PP_  (.D(_02091_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][17] ),
    .QN(_08186_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][18]$_DFFE_PP_  (.D(_02092_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][18] ),
    .QN(_08185_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][19]$_DFFE_PP_  (.D(_02093_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][19] ),
    .QN(_08184_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][1]$_DFFE_PP_  (.D(_02094_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][1] ),
    .QN(_08183_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][20]$_DFFE_PP_  (.D(_02095_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][20] ),
    .QN(_08182_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][21]$_DFFE_PP_  (.D(_02096_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][21] ),
    .QN(_08181_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][22]$_DFFE_PP_  (.D(_02097_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][22] ),
    .QN(_08180_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][23]$_DFFE_PP_  (.D(_02098_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][23] ),
    .QN(_08179_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][24]$_DFFE_PP_  (.D(_02099_),
    .CK(clknet_leaf_167_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][24] ),
    .QN(_08178_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][25]$_DFFE_PP_  (.D(_02100_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][25] ),
    .QN(_08177_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][26]$_DFFE_PP_  (.D(_02101_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][26] ),
    .QN(_08176_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][27]$_DFFE_PP_  (.D(_02102_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][27] ),
    .QN(_08175_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][28]$_DFFE_PP_  (.D(_02103_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][28] ),
    .QN(_08174_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][29]$_DFFE_PP_  (.D(_02104_),
    .CK(clknet_leaf_171_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][29] ),
    .QN(_08173_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][2]$_DFFE_PP_  (.D(_02105_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][2] ),
    .QN(_08172_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][30]$_DFFE_PP_  (.D(_02106_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][30] ),
    .QN(_08171_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][31]$_DFFE_PP_  (.D(_02107_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][31] ),
    .QN(_08170_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][32]$_DFFE_PP_  (.D(_02108_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][32] ),
    .QN(_08169_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][33]$_DFFE_PP_  (.D(_02109_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][33] ),
    .QN(_08168_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][34]$_DFFE_PP_  (.D(_02110_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][34] ),
    .QN(_08167_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][35]$_DFFE_PP_  (.D(_02111_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][35] ),
    .QN(_08166_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][36]$_DFFE_PP_  (.D(_02112_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][36] ),
    .QN(_08165_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][37]$_DFFE_PP_  (.D(_02113_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][37] ),
    .QN(_08164_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][38]$_DFFE_PP_  (.D(_02114_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][38] ),
    .QN(_08163_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][39]$_DFFE_PP_  (.D(_02115_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][39] ),
    .QN(_08162_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][3]$_DFFE_PP_  (.D(_02116_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][3] ),
    .QN(_08161_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][40]$_DFFE_PP_  (.D(_02117_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][40] ),
    .QN(_08160_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][41]$_DFFE_PP_  (.D(_02118_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][41] ),
    .QN(_08159_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][42]$_DFFE_PP_  (.D(_02119_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][42] ),
    .QN(_08158_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][43]$_DFFE_PP_  (.D(_02120_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][43] ),
    .QN(_08157_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][44]$_DFFE_PP_  (.D(_02121_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][44] ),
    .QN(_08156_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][45]$_DFFE_PP_  (.D(_02122_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][45] ),
    .QN(_08155_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][46]$_DFFE_PP_  (.D(_02123_),
    .CK(clknet_leaf_178_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][46] ),
    .QN(_08154_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][47]$_DFFE_PP_  (.D(_02124_),
    .CK(clknet_leaf_178_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][47] ),
    .QN(_08153_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][48]$_DFFE_PP_  (.D(_02125_),
    .CK(clknet_leaf_185_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][48] ),
    .QN(_08152_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][49]$_DFFE_PP_  (.D(_02126_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][49] ),
    .QN(_08151_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][4]$_DFFE_PP_  (.D(_02127_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][4] ),
    .QN(_08150_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][50]$_DFFE_PP_  (.D(_02128_),
    .CK(clknet_leaf_193_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][50] ),
    .QN(_08149_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][51]$_DFFE_PP_  (.D(_02129_),
    .CK(clknet_leaf_195_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][51] ),
    .QN(_08148_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][52]$_DFFE_PP_  (.D(_02130_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][52] ),
    .QN(_08147_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][53]$_DFFE_PP_  (.D(_02131_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][53] ),
    .QN(_08146_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][54]$_DFFE_PP_  (.D(_02132_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][54] ),
    .QN(_08145_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][55]$_DFFE_PP_  (.D(_02133_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][55] ),
    .QN(_08144_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][56]$_DFFE_PP_  (.D(_02134_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][56] ),
    .QN(_08143_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][57]$_DFFE_PP_  (.D(_02135_),
    .CK(clknet_leaf_190_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][57] ),
    .QN(_08142_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][58]$_DFFE_PP_  (.D(_02136_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][58] ),
    .QN(_08141_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][59]$_DFFE_PP_  (.D(_02137_),
    .CK(clknet_leaf_210_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][59] ),
    .QN(_08140_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][5]$_DFFE_PP_  (.D(_02138_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][5] ),
    .QN(_08139_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][60]$_DFFE_PP_  (.D(_02139_),
    .CK(clknet_leaf_190_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][60] ),
    .QN(_08138_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][61]$_DFFE_PP_  (.D(_02140_),
    .CK(clknet_leaf_195_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][61] ),
    .QN(_08137_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][62]$_DFFE_PP_  (.D(_02141_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][62] ),
    .QN(_08136_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][63]$_DFFE_PP_  (.D(_02142_),
    .CK(clknet_leaf_212_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][63] ),
    .QN(_08135_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][6]$_DFFE_PP_  (.D(_02143_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][6] ),
    .QN(_08134_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][7]$_DFFE_PP_  (.D(_02144_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][7] ),
    .QN(_08133_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][8]$_DFFE_PP_  (.D(_02145_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][8] ),
    .QN(_08132_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[1][9]$_DFFE_PP_  (.D(_02146_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[1][9] ),
    .QN(_08131_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][0]$_DFFE_PP_  (.D(_02147_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][0] ),
    .QN(_08130_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][10]$_DFFE_PP_  (.D(_02148_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][10] ),
    .QN(_08129_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][11]$_DFFE_PP_  (.D(_02149_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][11] ),
    .QN(_08128_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][12]$_DFFE_PP_  (.D(_02150_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][12] ),
    .QN(_08127_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][13]$_DFFE_PP_  (.D(_02151_),
    .CK(clknet_leaf_226_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][13] ),
    .QN(_08126_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][14]$_DFFE_PP_  (.D(_02152_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][14] ),
    .QN(_08125_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][15]$_DFFE_PP_  (.D(_02153_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][15] ),
    .QN(_08124_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][16]$_DFFE_PP_  (.D(_02154_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][16] ),
    .QN(_08123_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][17]$_DFFE_PP_  (.D(_02155_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][17] ),
    .QN(_08122_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][18]$_DFFE_PP_  (.D(_02156_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][18] ),
    .QN(_08121_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][19]$_DFFE_PP_  (.D(_02157_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][19] ),
    .QN(_08120_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][1]$_DFFE_PP_  (.D(_02158_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][1] ),
    .QN(_08119_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][20]$_DFFE_PP_  (.D(_02159_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][20] ),
    .QN(_08118_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][21]$_DFFE_PP_  (.D(_02160_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][21] ),
    .QN(_08117_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][22]$_DFFE_PP_  (.D(_02161_),
    .CK(clknet_leaf_166_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][22] ),
    .QN(_08116_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][23]$_DFFE_PP_  (.D(_02162_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][23] ),
    .QN(_08115_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][24]$_DFFE_PP_  (.D(_02163_),
    .CK(clknet_leaf_166_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][24] ),
    .QN(_08114_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][25]$_DFFE_PP_  (.D(_02164_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][25] ),
    .QN(_08113_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][26]$_DFFE_PP_  (.D(_02165_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][26] ),
    .QN(_08112_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][27]$_DFFE_PP_  (.D(_02166_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][27] ),
    .QN(_08111_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][28]$_DFFE_PP_  (.D(_02167_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][28] ),
    .QN(_08110_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][29]$_DFFE_PP_  (.D(_02168_),
    .CK(clknet_leaf_171_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][29] ),
    .QN(_08109_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][2]$_DFFE_PP_  (.D(_02169_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][2] ),
    .QN(_08108_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][30]$_DFFE_PP_  (.D(_02170_),
    .CK(clknet_leaf_170_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][30] ),
    .QN(_08107_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][31]$_DFFE_PP_  (.D(_02171_),
    .CK(clknet_leaf_174_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][31] ),
    .QN(_08106_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][32]$_DFFE_PP_  (.D(_02172_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][32] ),
    .QN(_08105_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][33]$_DFFE_PP_  (.D(_02173_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][33] ),
    .QN(_08104_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][34]$_DFFE_PP_  (.D(_02174_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][34] ),
    .QN(_08103_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][35]$_DFFE_PP_  (.D(_02175_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][35] ),
    .QN(_08102_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][36]$_DFFE_PP_  (.D(_02176_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][36] ),
    .QN(_08101_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][37]$_DFFE_PP_  (.D(_02177_),
    .CK(clknet_leaf_181_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][37] ),
    .QN(_08100_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][38]$_DFFE_PP_  (.D(_02178_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][38] ),
    .QN(_08099_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][39]$_DFFE_PP_  (.D(_02179_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][39] ),
    .QN(_08098_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][3]$_DFFE_PP_  (.D(_02180_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][3] ),
    .QN(_08097_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][40]$_DFFE_PP_  (.D(_02181_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][40] ),
    .QN(_08096_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][41]$_DFFE_PP_  (.D(_02182_),
    .CK(clknet_leaf_185_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][41] ),
    .QN(_08095_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][42]$_DFFE_PP_  (.D(_02183_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][42] ),
    .QN(_08094_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][43]$_DFFE_PP_  (.D(_02184_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][43] ),
    .QN(_08093_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][44]$_DFFE_PP_  (.D(_02185_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][44] ),
    .QN(_08092_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][45]$_DFFE_PP_  (.D(_02186_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][45] ),
    .QN(_08091_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][46]$_DFFE_PP_  (.D(_02187_),
    .CK(clknet_leaf_178_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][46] ),
    .QN(_08090_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][47]$_DFFE_PP_  (.D(_02188_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][47] ),
    .QN(_08089_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][48]$_DFFE_PP_  (.D(_02189_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][48] ),
    .QN(_08088_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][49]$_DFFE_PP_  (.D(_02190_),
    .CK(clknet_leaf_185_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][49] ),
    .QN(_08087_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][4]$_DFFE_PP_  (.D(_02191_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][4] ),
    .QN(_08086_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][50]$_DFFE_PP_  (.D(_02192_),
    .CK(clknet_leaf_193_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][50] ),
    .QN(_08085_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][51]$_DFFE_PP_  (.D(_02193_),
    .CK(clknet_leaf_177_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][51] ),
    .QN(_08084_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][52]$_DFFE_PP_  (.D(_02194_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][52] ),
    .QN(_08083_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][53]$_DFFE_PP_  (.D(_02195_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][53] ),
    .QN(_08082_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][54]$_DFFE_PP_  (.D(_02196_),
    .CK(clknet_leaf_195_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][54] ),
    .QN(_08081_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][55]$_DFFE_PP_  (.D(_02197_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][55] ),
    .QN(_08080_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][56]$_DFFE_PP_  (.D(_02198_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][56] ),
    .QN(_08079_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][57]$_DFFE_PP_  (.D(_02199_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][57] ),
    .QN(_08078_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][58]$_DFFE_PP_  (.D(_02200_),
    .CK(clknet_leaf_213_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][58] ),
    .QN(_08077_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][59]$_DFFE_PP_  (.D(_02201_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][59] ),
    .QN(_08076_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][5]$_DFFE_PP_  (.D(_02202_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][5] ),
    .QN(_08075_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][60]$_DFFE_PP_  (.D(_02203_),
    .CK(clknet_leaf_190_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][60] ),
    .QN(_08074_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][61]$_DFFE_PP_  (.D(_02204_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][61] ),
    .QN(_08073_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][62]$_DFFE_PP_  (.D(_02205_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][62] ),
    .QN(_08072_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][63]$_DFFE_PP_  (.D(_02206_),
    .CK(clknet_leaf_211_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][63] ),
    .QN(_08071_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][6]$_DFFE_PP_  (.D(_02207_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][6] ),
    .QN(_08070_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][7]$_DFFE_PP_  (.D(_02208_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][7] ),
    .QN(_08069_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][8]$_DFFE_PP_  (.D(_02209_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][8] ),
    .QN(_08068_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[2][9]$_DFFE_PP_  (.D(_02210_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[2][9] ),
    .QN(_08067_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][0]$_DFFE_PP_  (.D(_02211_),
    .CK(clknet_leaf_221_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][0] ),
    .QN(_08066_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][10]$_DFFE_PP_  (.D(_02212_),
    .CK(clknet_leaf_224_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][10] ),
    .QN(_08065_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][11]$_DFFE_PP_  (.D(_02213_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][11] ),
    .QN(_08064_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][12]$_DFFE_PP_  (.D(_02214_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][12] ),
    .QN(_08063_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][13]$_DFFE_PP_  (.D(_02215_),
    .CK(clknet_leaf_225_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][13] ),
    .QN(_08062_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][14]$_DFFE_PP_  (.D(_02216_),
    .CK(clknet_leaf_220_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][14] ),
    .QN(_08061_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][15]$_DFFE_PP_  (.D(_02217_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][15] ),
    .QN(_08060_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][16]$_DFFE_PP_  (.D(_02218_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][16] ),
    .QN(_08059_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][17]$_DFFE_PP_  (.D(_02219_),
    .CK(clknet_leaf_223_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][17] ),
    .QN(_08058_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][18]$_DFFE_PP_  (.D(_02220_),
    .CK(clknet_leaf_219_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][18] ),
    .QN(_08057_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][19]$_DFFE_PP_  (.D(_02221_),
    .CK(clknet_leaf_188_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][19] ),
    .QN(_08056_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][1]$_DFFE_PP_  (.D(_02222_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][1] ),
    .QN(_08055_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][20]$_DFFE_PP_  (.D(_02223_),
    .CK(clknet_leaf_189_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][20] ),
    .QN(_08054_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][21]$_DFFE_PP_  (.D(_02224_),
    .CK(clknet_leaf_217_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][21] ),
    .QN(_08053_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][22]$_DFFE_PP_  (.D(_02225_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][22] ),
    .QN(_08052_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][23]$_DFFE_PP_  (.D(_02226_),
    .CK(clknet_leaf_168_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][23] ),
    .QN(_08051_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][24]$_DFFE_PP_  (.D(_02227_),
    .CK(clknet_leaf_167_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][24] ),
    .QN(_08050_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][25]$_DFFE_PP_  (.D(_02228_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][25] ),
    .QN(_08049_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][26]$_DFFE_PP_  (.D(_02229_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][26] ),
    .QN(_08048_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][27]$_DFFE_PP_  (.D(_02230_),
    .CK(clknet_leaf_169_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][27] ),
    .QN(_08047_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][28]$_DFFE_PP_  (.D(_02231_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][28] ),
    .QN(_08046_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][29]$_DFFE_PP_  (.D(_02232_),
    .CK(clknet_leaf_171_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][29] ),
    .QN(_08045_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][2]$_DFFE_PP_  (.D(_02233_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][2] ),
    .QN(_08044_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][30]$_DFFE_PP_  (.D(_02234_),
    .CK(clknet_leaf_171_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][30] ),
    .QN(_08043_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][31]$_DFFE_PP_  (.D(_02235_),
    .CK(clknet_leaf_175_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][31] ),
    .QN(_08042_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][32]$_DFFE_PP_  (.D(_02236_),
    .CK(clknet_leaf_173_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][32] ),
    .QN(_08041_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][33]$_DFFE_PP_  (.D(_02237_),
    .CK(clknet_leaf_187_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][33] ),
    .QN(_08040_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][34]$_DFFE_PP_  (.D(_02238_),
    .CK(clknet_leaf_172_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][34] ),
    .QN(_08039_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][35]$_DFFE_PP_  (.D(_02239_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][35] ),
    .QN(_08038_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][36]$_DFFE_PP_  (.D(_02240_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][36] ),
    .QN(_08037_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][37]$_DFFE_PP_  (.D(_02241_),
    .CK(clknet_leaf_178_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][37] ),
    .QN(_08036_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][38]$_DFFE_PP_  (.D(_02242_),
    .CK(clknet_leaf_179_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][38] ),
    .QN(_08035_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][39]$_DFFE_PP_  (.D(_02243_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][39] ),
    .QN(_08034_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][3]$_DFFE_PP_  (.D(_02244_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][3] ),
    .QN(_08033_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][40]$_DFFE_PP_  (.D(_02245_),
    .CK(clknet_leaf_180_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][40] ),
    .QN(_08032_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][41]$_DFFE_PP_  (.D(_02246_),
    .CK(clknet_leaf_186_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][41] ),
    .QN(_08031_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][42]$_DFFE_PP_  (.D(_02247_),
    .CK(clknet_leaf_184_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][42] ),
    .QN(_08030_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][43]$_DFFE_PP_  (.D(_02248_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][43] ),
    .QN(_08029_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][44]$_DFFE_PP_  (.D(_02249_),
    .CK(clknet_leaf_182_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][44] ),
    .QN(_08028_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][45]$_DFFE_PP_  (.D(_02250_),
    .CK(clknet_leaf_183_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][45] ),
    .QN(_08027_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][46]$_DFFE_PP_  (.D(_02251_),
    .CK(clknet_leaf_178_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][46] ),
    .QN(_08026_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][47]$_DFFE_PP_  (.D(_02252_),
    .CK(clknet_leaf_178_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][47] ),
    .QN(_08025_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][48]$_DFFE_PP_  (.D(_02253_),
    .CK(clknet_leaf_185_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][48] ),
    .QN(_08024_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][49]$_DFFE_PP_  (.D(_02254_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][49] ),
    .QN(_08023_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][4]$_DFFE_PP_  (.D(_02255_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][4] ),
    .QN(_08022_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][50]$_DFFE_PP_  (.D(_02256_),
    .CK(clknet_leaf_193_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][50] ),
    .QN(_08021_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][51]$_DFFE_PP_  (.D(_02257_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][51] ),
    .QN(_08020_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][52]$_DFFE_PP_  (.D(_02258_),
    .CK(clknet_leaf_193_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][52] ),
    .QN(_08019_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][53]$_DFFE_PP_  (.D(_02259_),
    .CK(clknet_leaf_191_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][53] ),
    .QN(_08018_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][54]$_DFFE_PP_  (.D(_02260_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][54] ),
    .QN(_08017_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][55]$_DFFE_PP_  (.D(_02261_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][55] ),
    .QN(_08016_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][56]$_DFFE_PP_  (.D(_02262_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][56] ),
    .QN(_08015_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][57]$_DFFE_PP_  (.D(_02263_),
    .CK(clknet_leaf_190_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][57] ),
    .QN(_08014_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][58]$_DFFE_PP_  (.D(_02264_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][58] ),
    .QN(_08013_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][59]$_DFFE_PP_  (.D(_02265_),
    .CK(clknet_leaf_210_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][59] ),
    .QN(_08012_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][5]$_DFFE_PP_  (.D(_02266_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][5] ),
    .QN(_08011_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][60]$_DFFE_PP_  (.D(_02267_),
    .CK(clknet_leaf_190_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][60] ),
    .QN(_08010_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][61]$_DFFE_PP_  (.D(_02268_),
    .CK(clknet_leaf_194_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][61] ),
    .QN(_08009_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][62]$_DFFE_PP_  (.D(_02269_),
    .CK(clknet_leaf_215_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][62] ),
    .QN(_08008_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][63]$_DFFE_PP_  (.D(_02270_),
    .CK(clknet_leaf_210_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][63] ),
    .QN(_08007_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][6]$_DFFE_PP_  (.D(_02271_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][6] ),
    .QN(_08006_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][7]$_DFFE_PP_  (.D(_02272_),
    .CK(clknet_leaf_214_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][7] ),
    .QN(_08005_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][8]$_DFFE_PP_  (.D(_02273_),
    .CK(clknet_leaf_216_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][8] ),
    .QN(_08004_));
 DFF_X1 \dynamic_node_top.west_input.NIB.storage_data_f[3][9]$_DFFE_PP_  (.D(_02274_),
    .CK(clknet_leaf_218_clk),
    .Q(\dynamic_node_top.west_input.NIB.storage_data_f[3][9] ),
    .QN(_08003_));
 DFF_X1 \dynamic_node_top.west_input.NIB.tail_ptr_f[0]$_SDFFE_PP0N_  (.D(_02275_),
    .CK(clknet_leaf_192_clk),
    .Q(\dynamic_node_top.west_input.NIB.tail_ptr_f[0] ),
    .QN(\dynamic_node_top.west_input.NIB.tail_ptr_next[0] ));
 DFF_X1 \dynamic_node_top.west_input.NIB.tail_ptr_f[1]$_SDFFE_PP0N_  (.D(_02276_),
    .CK(clknet_leaf_185_clk),
    .Q(\dynamic_node_top.west_input.NIB.tail_ptr_f[1] ),
    .QN(_10609_));
 DFF_X1 \dynamic_node_top.west_input.NIB.yummy_out_f$_SDFF_PP0_  (.D(_02277_),
    .CK(clknet_leaf_162_clk),
    .Q(net630),
    .QN(_08002_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[0]$_SDFF_PP0_  (.D(_02278_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[0] ),
    .QN(_10479_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[1]$_SDFF_PP0_  (.D(_02279_),
    .CK(clknet_leaf_162_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[1] ),
    .QN(_10480_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[2]$_SDFF_PP0_  (.D(_02280_),
    .CK(clknet_leaf_165_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[2] ),
    .QN(_08001_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[3]$_SDFF_PP0_  (.D(_02281_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[3] ),
    .QN(_08000_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[4]$_SDFF_PP0_  (.D(_02282_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[4] ),
    .QN(_07999_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[5]$_SDFF_PP0_  (.D(_02283_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[5] ),
    .QN(_07998_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[6]$_SDFF_PP0_  (.D(_02284_),
    .CK(clknet_leaf_176_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[6] ),
    .QN(_07997_));
 DFF_X1 \dynamic_node_top.west_input.control.count_f[7]$_SDFF_PP0_  (.D(_02285_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.west_input.control.count_f[7] ),
    .QN(_07996_));
 DFF_X1 \dynamic_node_top.west_input.control.count_one_f$_SDFF_PP0_  (.D(_02286_),
    .CK(clknet_leaf_161_clk),
    .Q(\dynamic_node_top.west_input.control.count_one_f ),
    .QN(_10160_));
 DFF_X2 \dynamic_node_top.west_input.control.header_temp$_DFF_P_  (.D(_00004_),
    .CK(clknet_leaf_162_clk),
    .Q(\dynamic_node_top.west_input.control.header_last_temp ),
    .QN(_07995_));
 DFF_X1 \dynamic_node_top.west_input.control.tail_last_f$_SDFF_PP0_  (.D(_02287_),
    .CK(clknet_leaf_160_clk),
    .Q(\dynamic_node_top.west_input.control.tail_last_f ),
    .QN(_10161_));
 DFF_X2 \dynamic_node_top.west_output.control.current_route_f[0]$_DFF_P_  (.D(_00032_),
    .CK(clknet_leaf_142_clk),
    .Q(\dynamic_node_top.west_output.control.current_route_f[0] ),
    .QN(_00051_));
 DFF_X1 \dynamic_node_top.west_output.control.current_route_f[1]$_DFF_P_  (.D(_00033_),
    .CK(clknet_leaf_158_clk),
    .Q(\dynamic_node_top.west_output.control.current_route_f[1] ),
    .QN(_00050_));
 DFF_X1 \dynamic_node_top.west_output.control.current_route_f[2]$_DFF_P_  (.D(_00034_),
    .CK(clknet_leaf_142_clk),
    .Q(\dynamic_node_top.west_output.control.current_route_f[2] ),
    .QN(_00063_));
 DFF_X1 \dynamic_node_top.west_output.control.current_route_f[3]$_DFF_P_  (.D(_00035_),
    .CK(clknet_leaf_142_clk),
    .Q(\dynamic_node_top.west_output.control.current_route_f[3] ),
    .QN(_00064_));
 DFF_X1 \dynamic_node_top.west_output.control.current_route_f[4]$_DFF_P_  (.D(_00036_),
    .CK(clknet_leaf_143_clk),
    .Q(\dynamic_node_top.west_output.control.current_route_f[4] ),
    .QN(_00062_));
 DFF_X2 \dynamic_node_top.west_output.control.planned_f$_SDFF_PP0_  (.D(_02288_),
    .CK(clknet_leaf_158_clk),
    .Q(\dynamic_node_top.west_output.control.planned_f ),
    .QN(_00052_));
 DFF_X2 \dynamic_node_top.west_output.space.count_f[0]$_SDFF_PP0_  (.D(_02289_),
    .CK(clknet_leaf_164_clk),
    .Q(\dynamic_node_top.west_output.space.count_f[0] ),
    .QN(_10448_));
 DFF_X2 \dynamic_node_top.west_output.space.count_f[1]$_SDFF_PP0_  (.D(_02290_),
    .CK(clknet_leaf_164_clk),
    .Q(\dynamic_node_top.west_output.space.count_f[1] ),
    .QN(_10449_));
 DFF_X1 \dynamic_node_top.west_output.space.count_f[2]$_SDFF_PP1_  (.D(_02291_),
    .CK(clknet_leaf_164_clk),
    .Q(\dynamic_node_top.west_output.space.count_f[2] ),
    .QN(_00058_));
 DFF_X1 \dynamic_node_top.west_output.space.is_one_f$_SDFF_PP0_  (.D(_02292_),
    .CK(clknet_leaf_163_clk),
    .Q(\dynamic_node_top.west_output.space.is_one_f ),
    .QN(_07994_));
 DFF_X1 \dynamic_node_top.west_output.space.is_two_or_more_f$_SDFF_PP1_  (.D(_02293_),
    .CK(clknet_leaf_163_clk),
    .Q(\dynamic_node_top.west_output.space.is_two_or_more_f ),
    .QN(_07993_));
 DFF_X1 \dynamic_node_top.west_output.space.valid_f$_SDFF_PP0_  (.D(_02294_),
    .CK(clknet_leaf_163_clk),
    .Q(\dynamic_node_top.west_output.space.valid_f ),
    .QN(_10445_));
 DFF_X1 \dynamic_node_top.west_output.space.yummy_f$_SDFF_PP0_  (.D(_02295_),
    .CK(clknet_leaf_163_clk),
    .Q(\dynamic_node_top.west_output.space.yummy_f ),
    .QN(_10442_));
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_420 ();
 BUF_X1 input1 (.A(dataIn_E[0]),
    .Z(net3));
 BUF_X1 input2 (.A(dataIn_E[10]),
    .Z(net4));
 BUF_X1 input3 (.A(dataIn_E[11]),
    .Z(net5));
 BUF_X1 input4 (.A(dataIn_E[12]),
    .Z(net6));
 BUF_X1 input5 (.A(dataIn_E[13]),
    .Z(net7));
 BUF_X1 input6 (.A(dataIn_E[14]),
    .Z(net8));
 BUF_X1 input7 (.A(dataIn_E[15]),
    .Z(net9));
 BUF_X1 input8 (.A(dataIn_E[16]),
    .Z(net10));
 BUF_X1 input9 (.A(dataIn_E[17]),
    .Z(net11));
 BUF_X1 input10 (.A(dataIn_E[18]),
    .Z(net12));
 BUF_X1 input11 (.A(dataIn_E[19]),
    .Z(net13));
 BUF_X1 input12 (.A(dataIn_E[1]),
    .Z(net14));
 BUF_X1 input13 (.A(dataIn_E[20]),
    .Z(net15));
 BUF_X1 input14 (.A(dataIn_E[21]),
    .Z(net16));
 BUF_X1 input15 (.A(dataIn_E[22]),
    .Z(net17));
 BUF_X1 input16 (.A(dataIn_E[23]),
    .Z(net18));
 BUF_X1 input17 (.A(dataIn_E[24]),
    .Z(net19));
 BUF_X1 input18 (.A(dataIn_E[25]),
    .Z(net20));
 BUF_X1 input19 (.A(dataIn_E[26]),
    .Z(net21));
 BUF_X1 input20 (.A(dataIn_E[27]),
    .Z(net22));
 BUF_X1 input21 (.A(dataIn_E[28]),
    .Z(net23));
 BUF_X1 input22 (.A(dataIn_E[29]),
    .Z(net24));
 BUF_X1 input23 (.A(dataIn_E[2]),
    .Z(net25));
 BUF_X1 input24 (.A(dataIn_E[30]),
    .Z(net26));
 BUF_X1 input25 (.A(dataIn_E[31]),
    .Z(net27));
 BUF_X1 input26 (.A(dataIn_E[32]),
    .Z(net28));
 BUF_X1 input27 (.A(dataIn_E[33]),
    .Z(net29));
 BUF_X1 input28 (.A(dataIn_E[34]),
    .Z(net30));
 BUF_X1 input29 (.A(dataIn_E[35]),
    .Z(net31));
 BUF_X1 input30 (.A(dataIn_E[36]),
    .Z(net32));
 BUF_X1 input31 (.A(dataIn_E[37]),
    .Z(net33));
 BUF_X1 input32 (.A(dataIn_E[38]),
    .Z(net34));
 BUF_X1 input33 (.A(dataIn_E[39]),
    .Z(net35));
 BUF_X1 input34 (.A(dataIn_E[3]),
    .Z(net36));
 BUF_X1 input35 (.A(dataIn_E[40]),
    .Z(net37));
 BUF_X1 input36 (.A(dataIn_E[41]),
    .Z(net38));
 BUF_X1 input37 (.A(dataIn_E[42]),
    .Z(net39));
 BUF_X1 input38 (.A(dataIn_E[43]),
    .Z(net40));
 BUF_X1 input39 (.A(dataIn_E[44]),
    .Z(net41));
 BUF_X1 input40 (.A(dataIn_E[45]),
    .Z(net42));
 CLKBUF_X2 input41 (.A(dataIn_E[46]),
    .Z(net43));
 BUF_X1 input42 (.A(dataIn_E[47]),
    .Z(net44));
 BUF_X1 input43 (.A(dataIn_E[48]),
    .Z(net45));
 BUF_X1 input44 (.A(dataIn_E[49]),
    .Z(net46));
 BUF_X1 input45 (.A(dataIn_E[4]),
    .Z(net47));
 BUF_X2 input46 (.A(dataIn_E[50]),
    .Z(net48));
 BUF_X2 input47 (.A(dataIn_E[51]),
    .Z(net49));
 BUF_X2 input48 (.A(dataIn_E[52]),
    .Z(net50));
 BUF_X1 input49 (.A(dataIn_E[53]),
    .Z(net51));
 CLKBUF_X2 input50 (.A(dataIn_E[54]),
    .Z(net52));
 CLKBUF_X2 input51 (.A(dataIn_E[55]),
    .Z(net53));
 BUF_X1 input52 (.A(dataIn_E[56]),
    .Z(net54));
 CLKBUF_X2 input53 (.A(dataIn_E[57]),
    .Z(net55));
 BUF_X1 input54 (.A(dataIn_E[58]),
    .Z(net56));
 BUF_X1 input55 (.A(dataIn_E[59]),
    .Z(net57));
 CLKBUF_X2 input56 (.A(dataIn_E[5]),
    .Z(net58));
 BUF_X1 input57 (.A(dataIn_E[60]),
    .Z(net59));
 BUF_X1 input58 (.A(dataIn_E[61]),
    .Z(net60));
 BUF_X1 input59 (.A(dataIn_E[62]),
    .Z(net61));
 BUF_X1 input60 (.A(dataIn_E[63]),
    .Z(net62));
 BUF_X1 input61 (.A(dataIn_E[6]),
    .Z(net63));
 BUF_X1 input62 (.A(dataIn_E[7]),
    .Z(net64));
 BUF_X1 input63 (.A(dataIn_E[8]),
    .Z(net65));
 BUF_X1 input64 (.A(dataIn_E[9]),
    .Z(net66));
 CLKBUF_X2 input65 (.A(dataIn_N[0]),
    .Z(net67));
 BUF_X2 input66 (.A(dataIn_N[10]),
    .Z(net68));
 BUF_X2 input67 (.A(dataIn_N[11]),
    .Z(net69));
 CLKBUF_X2 input68 (.A(dataIn_N[12]),
    .Z(net70));
 BUF_X2 input69 (.A(dataIn_N[13]),
    .Z(net71));
 CLKBUF_X2 input70 (.A(dataIn_N[14]),
    .Z(net72));
 CLKBUF_X2 input71 (.A(dataIn_N[15]),
    .Z(net73));
 BUF_X2 input72 (.A(dataIn_N[16]),
    .Z(net74));
 BUF_X2 input73 (.A(dataIn_N[17]),
    .Z(net75));
 BUF_X2 input74 (.A(dataIn_N[18]),
    .Z(net76));
 BUF_X2 input75 (.A(dataIn_N[19]),
    .Z(net77));
 BUF_X2 input76 (.A(dataIn_N[1]),
    .Z(net78));
 BUF_X2 input77 (.A(dataIn_N[20]),
    .Z(net79));
 BUF_X2 input78 (.A(dataIn_N[21]),
    .Z(net80));
 BUF_X1 input79 (.A(dataIn_N[22]),
    .Z(net81));
 BUF_X1 input80 (.A(dataIn_N[23]),
    .Z(net82));
 BUF_X1 input81 (.A(dataIn_N[24]),
    .Z(net83));
 BUF_X1 input82 (.A(dataIn_N[25]),
    .Z(net84));
 BUF_X1 input83 (.A(dataIn_N[26]),
    .Z(net85));
 BUF_X1 input84 (.A(dataIn_N[27]),
    .Z(net86));
 BUF_X1 input85 (.A(dataIn_N[28]),
    .Z(net87));
 BUF_X1 input86 (.A(dataIn_N[29]),
    .Z(net88));
 CLKBUF_X2 input87 (.A(dataIn_N[2]),
    .Z(net89));
 BUF_X1 input88 (.A(dataIn_N[30]),
    .Z(net90));
 BUF_X1 input89 (.A(dataIn_N[31]),
    .Z(net91));
 BUF_X1 input90 (.A(dataIn_N[32]),
    .Z(net92));
 CLKBUF_X2 input91 (.A(dataIn_N[33]),
    .Z(net93));
 CLKBUF_X2 input92 (.A(dataIn_N[34]),
    .Z(net94));
 CLKBUF_X2 input93 (.A(dataIn_N[35]),
    .Z(net95));
 BUF_X1 input94 (.A(dataIn_N[36]),
    .Z(net96));
 CLKBUF_X2 input95 (.A(dataIn_N[37]),
    .Z(net97));
 CLKBUF_X2 input96 (.A(dataIn_N[38]),
    .Z(net98));
 CLKBUF_X2 input97 (.A(dataIn_N[39]),
    .Z(net99));
 BUF_X2 input98 (.A(dataIn_N[3]),
    .Z(net100));
 BUF_X1 input99 (.A(dataIn_N[40]),
    .Z(net101));
 BUF_X2 input100 (.A(dataIn_N[41]),
    .Z(net102));
 CLKBUF_X2 input101 (.A(dataIn_N[42]),
    .Z(net103));
 BUF_X2 input102 (.A(dataIn_N[43]),
    .Z(net104));
 CLKBUF_X2 input103 (.A(dataIn_N[44]),
    .Z(net105));
 CLKBUF_X2 input104 (.A(dataIn_N[45]),
    .Z(net106));
 BUF_X2 input105 (.A(dataIn_N[46]),
    .Z(net107));
 BUF_X2 input106 (.A(dataIn_N[47]),
    .Z(net108));
 BUF_X2 input107 (.A(dataIn_N[48]),
    .Z(net109));
 BUF_X2 input108 (.A(dataIn_N[49]),
    .Z(net110));
 BUF_X2 input109 (.A(dataIn_N[4]),
    .Z(net111));
 BUF_X2 input110 (.A(dataIn_N[50]),
    .Z(net112));
 BUF_X2 input111 (.A(dataIn_N[51]),
    .Z(net113));
 BUF_X2 input112 (.A(dataIn_N[52]),
    .Z(net114));
 BUF_X2 input113 (.A(dataIn_N[53]),
    .Z(net115));
 BUF_X2 input114 (.A(dataIn_N[54]),
    .Z(net116));
 BUF_X2 input115 (.A(dataIn_N[55]),
    .Z(net117));
 BUF_X2 input116 (.A(dataIn_N[56]),
    .Z(net118));
 BUF_X2 input117 (.A(dataIn_N[57]),
    .Z(net119));
 BUF_X2 input118 (.A(dataIn_N[58]),
    .Z(net120));
 BUF_X2 input119 (.A(dataIn_N[59]),
    .Z(net121));
 CLKBUF_X3 input120 (.A(dataIn_N[5]),
    .Z(net122));
 BUF_X2 input121 (.A(dataIn_N[60]),
    .Z(net123));
 BUF_X2 input122 (.A(dataIn_N[61]),
    .Z(net124));
 BUF_X2 input123 (.A(dataIn_N[62]),
    .Z(net125));
 BUF_X2 input124 (.A(dataIn_N[63]),
    .Z(net126));
 BUF_X2 input125 (.A(dataIn_N[6]),
    .Z(net127));
 BUF_X2 input126 (.A(dataIn_N[7]),
    .Z(net128));
 BUF_X2 input127 (.A(dataIn_N[8]),
    .Z(net129));
 BUF_X2 input128 (.A(dataIn_N[9]),
    .Z(net130));
 BUF_X1 input129 (.A(dataIn_S[0]),
    .Z(net131));
 BUF_X1 input130 (.A(dataIn_S[10]),
    .Z(net132));
 BUF_X1 input131 (.A(dataIn_S[11]),
    .Z(net133));
 BUF_X1 input132 (.A(dataIn_S[12]),
    .Z(net134));
 BUF_X1 input133 (.A(dataIn_S[13]),
    .Z(net135));
 BUF_X1 input134 (.A(dataIn_S[14]),
    .Z(net136));
 BUF_X1 input135 (.A(dataIn_S[15]),
    .Z(net137));
 BUF_X1 input136 (.A(dataIn_S[16]),
    .Z(net138));
 BUF_X1 input137 (.A(dataIn_S[17]),
    .Z(net139));
 BUF_X1 input138 (.A(dataIn_S[18]),
    .Z(net140));
 BUF_X1 input139 (.A(dataIn_S[19]),
    .Z(net141));
 BUF_X1 input140 (.A(dataIn_S[1]),
    .Z(net142));
 BUF_X1 input141 (.A(dataIn_S[20]),
    .Z(net143));
 BUF_X1 input142 (.A(dataIn_S[21]),
    .Z(net144));
 BUF_X1 input143 (.A(dataIn_S[22]),
    .Z(net145));
 BUF_X1 input144 (.A(dataIn_S[23]),
    .Z(net146));
 BUF_X1 input145 (.A(dataIn_S[24]),
    .Z(net147));
 BUF_X1 input146 (.A(dataIn_S[25]),
    .Z(net148));
 BUF_X1 input147 (.A(dataIn_S[26]),
    .Z(net149));
 BUF_X1 input148 (.A(dataIn_S[27]),
    .Z(net150));
 BUF_X1 input149 (.A(dataIn_S[28]),
    .Z(net151));
 BUF_X1 input150 (.A(dataIn_S[29]),
    .Z(net152));
 BUF_X1 input151 (.A(dataIn_S[2]),
    .Z(net153));
 BUF_X1 input152 (.A(dataIn_S[30]),
    .Z(net154));
 BUF_X1 input153 (.A(dataIn_S[31]),
    .Z(net155));
 BUF_X1 input154 (.A(dataIn_S[32]),
    .Z(net156));
 BUF_X1 input155 (.A(dataIn_S[33]),
    .Z(net157));
 BUF_X1 input156 (.A(dataIn_S[34]),
    .Z(net158));
 BUF_X1 input157 (.A(dataIn_S[35]),
    .Z(net159));
 BUF_X1 input158 (.A(dataIn_S[36]),
    .Z(net160));
 BUF_X1 input159 (.A(dataIn_S[37]),
    .Z(net161));
 BUF_X1 input160 (.A(dataIn_S[38]),
    .Z(net162));
 BUF_X1 input161 (.A(dataIn_S[39]),
    .Z(net163));
 BUF_X1 input162 (.A(dataIn_S[3]),
    .Z(net164));
 CLKBUF_X2 input163 (.A(dataIn_S[40]),
    .Z(net165));
 BUF_X1 input164 (.A(dataIn_S[41]),
    .Z(net166));
 BUF_X1 input165 (.A(dataIn_S[42]),
    .Z(net167));
 CLKBUF_X2 input166 (.A(dataIn_S[43]),
    .Z(net168));
 CLKBUF_X2 input167 (.A(dataIn_S[44]),
    .Z(net169));
 BUF_X1 input168 (.A(dataIn_S[45]),
    .Z(net170));
 BUF_X1 input169 (.A(dataIn_S[46]),
    .Z(net171));
 CLKBUF_X2 input170 (.A(dataIn_S[47]),
    .Z(net172));
 BUF_X1 input171 (.A(dataIn_S[48]),
    .Z(net173));
 BUF_X1 input172 (.A(dataIn_S[49]),
    .Z(net174));
 BUF_X1 input173 (.A(dataIn_S[4]),
    .Z(net175));
 BUF_X1 input174 (.A(dataIn_S[50]),
    .Z(net176));
 BUF_X1 input175 (.A(dataIn_S[51]),
    .Z(net177));
 BUF_X1 input176 (.A(dataIn_S[52]),
    .Z(net178));
 BUF_X1 input177 (.A(dataIn_S[53]),
    .Z(net179));
 BUF_X1 input178 (.A(dataIn_S[54]),
    .Z(net180));
 BUF_X1 input179 (.A(dataIn_S[55]),
    .Z(net181));
 BUF_X1 input180 (.A(dataIn_S[56]),
    .Z(net182));
 BUF_X2 input181 (.A(dataIn_S[57]),
    .Z(net183));
 BUF_X1 input182 (.A(dataIn_S[58]),
    .Z(net184));
 CLKBUF_X2 input183 (.A(dataIn_S[59]),
    .Z(net185));
 BUF_X1 input184 (.A(dataIn_S[5]),
    .Z(net186));
 BUF_X1 input185 (.A(dataIn_S[60]),
    .Z(net187));
 BUF_X1 input186 (.A(dataIn_S[61]),
    .Z(net188));
 BUF_X1 input187 (.A(dataIn_S[62]),
    .Z(net189));
 BUF_X1 input188 (.A(dataIn_S[63]),
    .Z(net190));
 BUF_X1 input189 (.A(dataIn_S[6]),
    .Z(net191));
 BUF_X1 input190 (.A(dataIn_S[7]),
    .Z(net192));
 BUF_X1 input191 (.A(dataIn_S[8]),
    .Z(net193));
 BUF_X1 input192 (.A(dataIn_S[9]),
    .Z(net194));
 BUF_X1 input193 (.A(dataIn_W[0]),
    .Z(net195));
 BUF_X1 input194 (.A(dataIn_W[10]),
    .Z(net196));
 BUF_X1 input195 (.A(dataIn_W[11]),
    .Z(net197));
 BUF_X1 input196 (.A(dataIn_W[12]),
    .Z(net198));
 BUF_X1 input197 (.A(dataIn_W[13]),
    .Z(net199));
 BUF_X1 input198 (.A(dataIn_W[14]),
    .Z(net200));
 BUF_X1 input199 (.A(dataIn_W[15]),
    .Z(net201));
 BUF_X1 input200 (.A(dataIn_W[16]),
    .Z(net202));
 BUF_X1 input201 (.A(dataIn_W[17]),
    .Z(net203));
 BUF_X1 input202 (.A(dataIn_W[18]),
    .Z(net204));
 BUF_X1 input203 (.A(dataIn_W[19]),
    .Z(net205));
 BUF_X1 input204 (.A(dataIn_W[1]),
    .Z(net206));
 BUF_X1 input205 (.A(dataIn_W[20]),
    .Z(net207));
 BUF_X1 input206 (.A(dataIn_W[21]),
    .Z(net208));
 BUF_X1 input207 (.A(dataIn_W[22]),
    .Z(net209));
 BUF_X1 input208 (.A(dataIn_W[23]),
    .Z(net210));
 BUF_X1 input209 (.A(dataIn_W[24]),
    .Z(net211));
 BUF_X1 input210 (.A(dataIn_W[25]),
    .Z(net212));
 BUF_X1 input211 (.A(dataIn_W[26]),
    .Z(net213));
 BUF_X1 input212 (.A(dataIn_W[27]),
    .Z(net214));
 BUF_X1 input213 (.A(dataIn_W[28]),
    .Z(net215));
 BUF_X1 input214 (.A(dataIn_W[29]),
    .Z(net216));
 BUF_X1 input215 (.A(dataIn_W[2]),
    .Z(net217));
 BUF_X1 input216 (.A(dataIn_W[30]),
    .Z(net218));
 BUF_X1 input217 (.A(dataIn_W[31]),
    .Z(net219));
 BUF_X1 input218 (.A(dataIn_W[32]),
    .Z(net220));
 BUF_X1 input219 (.A(dataIn_W[33]),
    .Z(net221));
 BUF_X1 input220 (.A(dataIn_W[34]),
    .Z(net222));
 BUF_X1 input221 (.A(dataIn_W[35]),
    .Z(net223));
 BUF_X1 input222 (.A(dataIn_W[36]),
    .Z(net224));
 BUF_X1 input223 (.A(dataIn_W[37]),
    .Z(net225));
 BUF_X1 input224 (.A(dataIn_W[38]),
    .Z(net226));
 BUF_X1 input225 (.A(dataIn_W[39]),
    .Z(net227));
 BUF_X1 input226 (.A(dataIn_W[3]),
    .Z(net228));
 BUF_X1 input227 (.A(dataIn_W[40]),
    .Z(net229));
 CLKBUF_X2 input228 (.A(dataIn_W[41]),
    .Z(net230));
 BUF_X1 input229 (.A(dataIn_W[42]),
    .Z(net231));
 CLKBUF_X2 input230 (.A(dataIn_W[43]),
    .Z(net232));
 BUF_X1 input231 (.A(dataIn_W[44]),
    .Z(net233));
 BUF_X1 input232 (.A(dataIn_W[45]),
    .Z(net234));
 BUF_X1 input233 (.A(dataIn_W[46]),
    .Z(net235));
 BUF_X1 input234 (.A(dataIn_W[47]),
    .Z(net236));
 BUF_X1 input235 (.A(dataIn_W[48]),
    .Z(net237));
 BUF_X1 input236 (.A(dataIn_W[49]),
    .Z(net238));
 BUF_X2 input237 (.A(dataIn_W[4]),
    .Z(net239));
 BUF_X1 input238 (.A(dataIn_W[50]),
    .Z(net240));
 BUF_X1 input239 (.A(dataIn_W[51]),
    .Z(net241));
 BUF_X1 input240 (.A(dataIn_W[52]),
    .Z(net242));
 BUF_X1 input241 (.A(dataIn_W[53]),
    .Z(net243));
 BUF_X2 input242 (.A(dataIn_W[54]),
    .Z(net244));
 BUF_X1 input243 (.A(dataIn_W[55]),
    .Z(net245));
 BUF_X1 input244 (.A(dataIn_W[56]),
    .Z(net246));
 BUF_X1 input245 (.A(dataIn_W[57]),
    .Z(net247));
 BUF_X1 input246 (.A(dataIn_W[58]),
    .Z(net248));
 BUF_X1 input247 (.A(dataIn_W[59]),
    .Z(net249));
 BUF_X1 input248 (.A(dataIn_W[5]),
    .Z(net250));
 BUF_X1 input249 (.A(dataIn_W[60]),
    .Z(net251));
 BUF_X1 input250 (.A(dataIn_W[61]),
    .Z(net252));
 BUF_X1 input251 (.A(dataIn_W[62]),
    .Z(net253));
 BUF_X1 input252 (.A(dataIn_W[63]),
    .Z(net254));
 BUF_X1 input253 (.A(dataIn_W[6]),
    .Z(net255));
 BUF_X1 input254 (.A(dataIn_W[7]),
    .Z(net256));
 BUF_X1 input255 (.A(dataIn_W[8]),
    .Z(net257));
 BUF_X1 input256 (.A(dataIn_W[9]),
    .Z(net258));
 BUF_X1 input257 (.A(myChipID[0]),
    .Z(net259));
 BUF_X1 input258 (.A(myChipID[10]),
    .Z(net260));
 BUF_X1 input259 (.A(myChipID[11]),
    .Z(net261));
 BUF_X1 input260 (.A(myChipID[12]),
    .Z(net262));
 CLKBUF_X2 input261 (.A(myChipID[13]),
    .Z(net263));
 BUF_X1 input262 (.A(myChipID[1]),
    .Z(net264));
 BUF_X1 input263 (.A(myChipID[2]),
    .Z(net265));
 BUF_X1 input264 (.A(myChipID[3]),
    .Z(net266));
 BUF_X1 input265 (.A(myChipID[4]),
    .Z(net267));
 BUF_X1 input266 (.A(myChipID[5]),
    .Z(net268));
 CLKBUF_X2 input267 (.A(myChipID[6]),
    .Z(net269));
 BUF_X1 input268 (.A(myChipID[7]),
    .Z(net270));
 BUF_X1 input269 (.A(myChipID[8]),
    .Z(net271));
 BUF_X1 input270 (.A(myChipID[9]),
    .Z(net272));
 BUF_X1 input271 (.A(myLocX[0]),
    .Z(net273));
 BUF_X1 input272 (.A(myLocX[1]),
    .Z(net274));
 BUF_X1 input273 (.A(myLocX[2]),
    .Z(net275));
 BUF_X1 input274 (.A(myLocX[3]),
    .Z(net276));
 BUF_X1 input275 (.A(myLocX[4]),
    .Z(net277));
 BUF_X1 input276 (.A(myLocX[5]),
    .Z(net278));
 BUF_X1 input277 (.A(myLocX[6]),
    .Z(net279));
 BUF_X1 input278 (.A(myLocX[7]),
    .Z(net280));
 BUF_X1 input279 (.A(myLocY[0]),
    .Z(net281));
 BUF_X1 input280 (.A(myLocY[1]),
    .Z(net282));
 BUF_X1 input281 (.A(myLocY[2]),
    .Z(net283));
 BUF_X1 input282 (.A(myLocY[3]),
    .Z(net284));
 BUF_X1 input283 (.A(myLocY[4]),
    .Z(net285));
 BUF_X1 input284 (.A(myLocY[5]),
    .Z(net286));
 BUF_X1 input285 (.A(myLocY[6]),
    .Z(net287));
 BUF_X1 input286 (.A(myLocY[7]),
    .Z(net288));
 BUF_X1 input287 (.A(reset_in),
    .Z(net289));
 CLKBUF_X2 input288 (.A(validIn_E),
    .Z(net290));
 BUF_X1 input289 (.A(validIn_N),
    .Z(net291));
 BUF_X1 input290 (.A(validIn_P),
    .Z(net292));
 CLKBUF_X2 input291 (.A(validIn_S),
    .Z(net293));
 BUF_X1 input292 (.A(validIn_W),
    .Z(net294));
 BUF_X1 input293 (.A(yummyIn_E),
    .Z(net295));
 BUF_X1 input294 (.A(yummyIn_N),
    .Z(net296));
 BUF_X1 input295 (.A(yummyIn_P),
    .Z(net297));
 BUF_X1 input296 (.A(yummyIn_S),
    .Z(net298));
 BUF_X1 input297 (.A(yummyIn_W),
    .Z(net299));
 BUF_X1 output298 (.A(net300),
    .Z(dataOut_E[0]));
 BUF_X1 output299 (.A(net301),
    .Z(dataOut_E[10]));
 BUF_X1 output300 (.A(net302),
    .Z(dataOut_E[11]));
 BUF_X1 output301 (.A(net303),
    .Z(dataOut_E[12]));
 BUF_X1 output302 (.A(net304),
    .Z(dataOut_E[13]));
 BUF_X1 output303 (.A(net305),
    .Z(dataOut_E[14]));
 BUF_X1 output304 (.A(net306),
    .Z(dataOut_E[15]));
 BUF_X1 output305 (.A(net307),
    .Z(dataOut_E[16]));
 BUF_X1 output306 (.A(net308),
    .Z(dataOut_E[17]));
 BUF_X1 output307 (.A(net309),
    .Z(dataOut_E[18]));
 BUF_X1 output308 (.A(net310),
    .Z(dataOut_E[19]));
 BUF_X1 output309 (.A(net311),
    .Z(dataOut_E[1]));
 BUF_X1 output310 (.A(net312),
    .Z(dataOut_E[20]));
 BUF_X1 output311 (.A(net313),
    .Z(dataOut_E[21]));
 BUF_X1 output312 (.A(net314),
    .Z(dataOut_E[22]));
 BUF_X1 output313 (.A(net315),
    .Z(dataOut_E[23]));
 BUF_X1 output314 (.A(net316),
    .Z(dataOut_E[24]));
 BUF_X1 output315 (.A(net317),
    .Z(dataOut_E[25]));
 BUF_X1 output316 (.A(net318),
    .Z(dataOut_E[26]));
 BUF_X1 output317 (.A(net319),
    .Z(dataOut_E[27]));
 BUF_X1 output318 (.A(net320),
    .Z(dataOut_E[28]));
 BUF_X1 output319 (.A(net321),
    .Z(dataOut_E[29]));
 BUF_X1 output320 (.A(net322),
    .Z(dataOut_E[2]));
 BUF_X1 output321 (.A(net323),
    .Z(dataOut_E[30]));
 BUF_X1 output322 (.A(net324),
    .Z(dataOut_E[31]));
 BUF_X1 output323 (.A(net325),
    .Z(dataOut_E[32]));
 BUF_X1 output324 (.A(net326),
    .Z(dataOut_E[33]));
 BUF_X1 output325 (.A(net327),
    .Z(dataOut_E[34]));
 BUF_X1 output326 (.A(net328),
    .Z(dataOut_E[35]));
 BUF_X1 output327 (.A(net329),
    .Z(dataOut_E[36]));
 BUF_X1 output328 (.A(net330),
    .Z(dataOut_E[37]));
 BUF_X1 output329 (.A(net331),
    .Z(dataOut_E[38]));
 BUF_X1 output330 (.A(net332),
    .Z(dataOut_E[39]));
 BUF_X1 output331 (.A(net333),
    .Z(dataOut_E[3]));
 BUF_X1 output332 (.A(net334),
    .Z(dataOut_E[40]));
 BUF_X1 output333 (.A(net335),
    .Z(dataOut_E[41]));
 BUF_X1 output334 (.A(net336),
    .Z(dataOut_E[42]));
 BUF_X1 output335 (.A(net337),
    .Z(dataOut_E[43]));
 BUF_X1 output336 (.A(net338),
    .Z(dataOut_E[44]));
 BUF_X1 output337 (.A(net339),
    .Z(dataOut_E[45]));
 BUF_X1 output338 (.A(net340),
    .Z(dataOut_E[46]));
 BUF_X1 output339 (.A(net341),
    .Z(dataOut_E[47]));
 BUF_X1 output340 (.A(net342),
    .Z(dataOut_E[48]));
 BUF_X1 output341 (.A(net343),
    .Z(dataOut_E[49]));
 BUF_X1 output342 (.A(net344),
    .Z(dataOut_E[4]));
 BUF_X1 output343 (.A(net345),
    .Z(dataOut_E[50]));
 BUF_X1 output344 (.A(net346),
    .Z(dataOut_E[51]));
 BUF_X1 output345 (.A(net347),
    .Z(dataOut_E[52]));
 BUF_X1 output346 (.A(net348),
    .Z(dataOut_E[53]));
 BUF_X1 output347 (.A(net349),
    .Z(dataOut_E[54]));
 BUF_X1 output348 (.A(net350),
    .Z(dataOut_E[55]));
 BUF_X1 output349 (.A(net351),
    .Z(dataOut_E[56]));
 BUF_X1 output350 (.A(net352),
    .Z(dataOut_E[57]));
 BUF_X1 output351 (.A(net353),
    .Z(dataOut_E[58]));
 BUF_X1 output352 (.A(net354),
    .Z(dataOut_E[59]));
 BUF_X1 output353 (.A(net355),
    .Z(dataOut_E[5]));
 BUF_X1 output354 (.A(net356),
    .Z(dataOut_E[60]));
 BUF_X1 output355 (.A(net357),
    .Z(dataOut_E[61]));
 BUF_X1 output356 (.A(net358),
    .Z(dataOut_E[62]));
 BUF_X1 output357 (.A(net359),
    .Z(dataOut_E[63]));
 BUF_X1 output358 (.A(net360),
    .Z(dataOut_E[6]));
 BUF_X1 output359 (.A(net361),
    .Z(dataOut_E[7]));
 BUF_X1 output360 (.A(net362),
    .Z(dataOut_E[8]));
 BUF_X1 output361 (.A(net363),
    .Z(dataOut_E[9]));
 BUF_X1 output362 (.A(net364),
    .Z(dataOut_N[0]));
 BUF_X1 output363 (.A(net365),
    .Z(dataOut_N[10]));
 BUF_X1 output364 (.A(net366),
    .Z(dataOut_N[11]));
 BUF_X1 output365 (.A(net367),
    .Z(dataOut_N[12]));
 BUF_X1 output366 (.A(net368),
    .Z(dataOut_N[13]));
 BUF_X1 output367 (.A(net369),
    .Z(dataOut_N[14]));
 BUF_X1 output368 (.A(net370),
    .Z(dataOut_N[15]));
 BUF_X1 output369 (.A(net371),
    .Z(dataOut_N[16]));
 BUF_X1 output370 (.A(net372),
    .Z(dataOut_N[17]));
 BUF_X1 output371 (.A(net373),
    .Z(dataOut_N[18]));
 BUF_X1 output372 (.A(net374),
    .Z(dataOut_N[19]));
 BUF_X1 output373 (.A(net375),
    .Z(dataOut_N[1]));
 BUF_X1 output374 (.A(net376),
    .Z(dataOut_N[20]));
 BUF_X1 output375 (.A(net377),
    .Z(dataOut_N[21]));
 BUF_X1 output376 (.A(net378),
    .Z(dataOut_N[22]));
 BUF_X1 output377 (.A(net379),
    .Z(dataOut_N[23]));
 BUF_X1 output378 (.A(net380),
    .Z(dataOut_N[24]));
 BUF_X1 output379 (.A(net381),
    .Z(dataOut_N[25]));
 BUF_X1 output380 (.A(net382),
    .Z(dataOut_N[26]));
 BUF_X1 output381 (.A(net383),
    .Z(dataOut_N[27]));
 BUF_X1 output382 (.A(net384),
    .Z(dataOut_N[28]));
 BUF_X1 output383 (.A(net385),
    .Z(dataOut_N[29]));
 BUF_X1 output384 (.A(net386),
    .Z(dataOut_N[2]));
 BUF_X1 output385 (.A(net387),
    .Z(dataOut_N[30]));
 BUF_X1 output386 (.A(net388),
    .Z(dataOut_N[31]));
 BUF_X1 output387 (.A(net389),
    .Z(dataOut_N[32]));
 BUF_X1 output388 (.A(net390),
    .Z(dataOut_N[33]));
 BUF_X1 output389 (.A(net391),
    .Z(dataOut_N[34]));
 BUF_X1 output390 (.A(net392),
    .Z(dataOut_N[35]));
 BUF_X1 output391 (.A(net393),
    .Z(dataOut_N[36]));
 BUF_X1 output392 (.A(net394),
    .Z(dataOut_N[37]));
 BUF_X1 output393 (.A(net395),
    .Z(dataOut_N[38]));
 BUF_X1 output394 (.A(net396),
    .Z(dataOut_N[39]));
 BUF_X1 output395 (.A(net397),
    .Z(dataOut_N[3]));
 BUF_X1 output396 (.A(net398),
    .Z(dataOut_N[40]));
 BUF_X1 output397 (.A(net399),
    .Z(dataOut_N[41]));
 BUF_X1 output398 (.A(net400),
    .Z(dataOut_N[42]));
 BUF_X1 output399 (.A(net401),
    .Z(dataOut_N[43]));
 BUF_X1 output400 (.A(net402),
    .Z(dataOut_N[44]));
 BUF_X1 output401 (.A(net403),
    .Z(dataOut_N[45]));
 BUF_X1 output402 (.A(net404),
    .Z(dataOut_N[46]));
 BUF_X1 output403 (.A(net405),
    .Z(dataOut_N[47]));
 BUF_X1 output404 (.A(net406),
    .Z(dataOut_N[48]));
 BUF_X1 output405 (.A(net407),
    .Z(dataOut_N[49]));
 BUF_X1 output406 (.A(net408),
    .Z(dataOut_N[4]));
 BUF_X1 output407 (.A(net409),
    .Z(dataOut_N[50]));
 BUF_X1 output408 (.A(net410),
    .Z(dataOut_N[51]));
 BUF_X1 output409 (.A(net411),
    .Z(dataOut_N[52]));
 BUF_X1 output410 (.A(net412),
    .Z(dataOut_N[53]));
 BUF_X1 output411 (.A(net413),
    .Z(dataOut_N[54]));
 BUF_X1 output412 (.A(net414),
    .Z(dataOut_N[55]));
 BUF_X1 output413 (.A(net415),
    .Z(dataOut_N[56]));
 BUF_X1 output414 (.A(net416),
    .Z(dataOut_N[57]));
 BUF_X1 output415 (.A(net417),
    .Z(dataOut_N[58]));
 BUF_X1 output416 (.A(net418),
    .Z(dataOut_N[59]));
 BUF_X1 output417 (.A(net419),
    .Z(dataOut_N[5]));
 BUF_X1 output418 (.A(net420),
    .Z(dataOut_N[60]));
 BUF_X1 output419 (.A(net421),
    .Z(dataOut_N[61]));
 BUF_X1 output420 (.A(net422),
    .Z(dataOut_N[62]));
 BUF_X1 output421 (.A(net423),
    .Z(dataOut_N[63]));
 BUF_X1 output422 (.A(net424),
    .Z(dataOut_N[6]));
 BUF_X1 output423 (.A(net425),
    .Z(dataOut_N[7]));
 BUF_X1 output424 (.A(net426),
    .Z(dataOut_N[8]));
 BUF_X1 output425 (.A(net427),
    .Z(dataOut_N[9]));
 BUF_X1 output426 (.A(net428),
    .Z(dataOut_P[0]));
 BUF_X1 output427 (.A(net429),
    .Z(dataOut_P[10]));
 BUF_X1 output428 (.A(net430),
    .Z(dataOut_P[11]));
 BUF_X1 output429 (.A(net431),
    .Z(dataOut_P[12]));
 BUF_X1 output430 (.A(net432),
    .Z(dataOut_P[13]));
 BUF_X1 output431 (.A(net433),
    .Z(dataOut_P[14]));
 BUF_X1 output432 (.A(net434),
    .Z(dataOut_P[15]));
 BUF_X1 output433 (.A(net435),
    .Z(dataOut_P[16]));
 BUF_X1 output434 (.A(net436),
    .Z(dataOut_P[17]));
 BUF_X1 output435 (.A(net437),
    .Z(dataOut_P[18]));
 BUF_X1 output436 (.A(net438),
    .Z(dataOut_P[19]));
 BUF_X1 output437 (.A(net439),
    .Z(dataOut_P[1]));
 BUF_X1 output438 (.A(net440),
    .Z(dataOut_P[20]));
 BUF_X1 output439 (.A(net441),
    .Z(dataOut_P[21]));
 BUF_X1 output440 (.A(net442),
    .Z(dataOut_P[22]));
 BUF_X1 output441 (.A(net443),
    .Z(dataOut_P[23]));
 BUF_X1 output442 (.A(net444),
    .Z(dataOut_P[24]));
 BUF_X1 output443 (.A(net445),
    .Z(dataOut_P[25]));
 BUF_X1 output444 (.A(net446),
    .Z(dataOut_P[26]));
 BUF_X1 output445 (.A(net447),
    .Z(dataOut_P[27]));
 BUF_X1 output446 (.A(net448),
    .Z(dataOut_P[28]));
 BUF_X1 output447 (.A(net449),
    .Z(dataOut_P[29]));
 BUF_X1 output448 (.A(net450),
    .Z(dataOut_P[2]));
 BUF_X1 output449 (.A(net451),
    .Z(dataOut_P[30]));
 BUF_X1 output450 (.A(net452),
    .Z(dataOut_P[31]));
 BUF_X1 output451 (.A(net453),
    .Z(dataOut_P[32]));
 BUF_X1 output452 (.A(net454),
    .Z(dataOut_P[33]));
 BUF_X1 output453 (.A(net455),
    .Z(dataOut_P[34]));
 BUF_X1 output454 (.A(net456),
    .Z(dataOut_P[35]));
 BUF_X1 output455 (.A(net457),
    .Z(dataOut_P[36]));
 BUF_X1 output456 (.A(net458),
    .Z(dataOut_P[37]));
 BUF_X1 output457 (.A(net459),
    .Z(dataOut_P[38]));
 BUF_X1 output458 (.A(net460),
    .Z(dataOut_P[39]));
 BUF_X1 output459 (.A(net461),
    .Z(dataOut_P[3]));
 BUF_X1 output460 (.A(net462),
    .Z(dataOut_P[40]));
 BUF_X1 output461 (.A(net463),
    .Z(dataOut_P[41]));
 BUF_X1 output462 (.A(net464),
    .Z(dataOut_P[42]));
 BUF_X1 output463 (.A(net465),
    .Z(dataOut_P[43]));
 BUF_X1 output464 (.A(net466),
    .Z(dataOut_P[44]));
 BUF_X1 output465 (.A(net467),
    .Z(dataOut_P[45]));
 BUF_X1 output466 (.A(net468),
    .Z(dataOut_P[46]));
 BUF_X1 output467 (.A(net469),
    .Z(dataOut_P[47]));
 BUF_X1 output468 (.A(net470),
    .Z(dataOut_P[48]));
 BUF_X1 output469 (.A(net471),
    .Z(dataOut_P[49]));
 BUF_X1 output470 (.A(net472),
    .Z(dataOut_P[4]));
 BUF_X1 output471 (.A(net473),
    .Z(dataOut_P[50]));
 BUF_X1 output472 (.A(net474),
    .Z(dataOut_P[51]));
 BUF_X1 output473 (.A(net475),
    .Z(dataOut_P[52]));
 BUF_X1 output474 (.A(net476),
    .Z(dataOut_P[53]));
 BUF_X1 output475 (.A(net477),
    .Z(dataOut_P[54]));
 BUF_X1 output476 (.A(net478),
    .Z(dataOut_P[55]));
 BUF_X1 output477 (.A(net479),
    .Z(dataOut_P[56]));
 BUF_X1 output478 (.A(net480),
    .Z(dataOut_P[57]));
 BUF_X1 output479 (.A(net481),
    .Z(dataOut_P[58]));
 BUF_X1 output480 (.A(net482),
    .Z(dataOut_P[59]));
 BUF_X1 output481 (.A(net483),
    .Z(dataOut_P[5]));
 BUF_X1 output482 (.A(net484),
    .Z(dataOut_P[60]));
 BUF_X1 output483 (.A(net485),
    .Z(dataOut_P[61]));
 BUF_X1 output484 (.A(net486),
    .Z(dataOut_P[62]));
 BUF_X1 output485 (.A(net487),
    .Z(dataOut_P[63]));
 BUF_X1 output486 (.A(net488),
    .Z(dataOut_P[6]));
 BUF_X1 output487 (.A(net489),
    .Z(dataOut_P[7]));
 BUF_X1 output488 (.A(net490),
    .Z(dataOut_P[8]));
 BUF_X1 output489 (.A(net491),
    .Z(dataOut_P[9]));
 BUF_X1 output490 (.A(net492),
    .Z(dataOut_S[0]));
 BUF_X1 output491 (.A(net493),
    .Z(dataOut_S[10]));
 BUF_X1 output492 (.A(net494),
    .Z(dataOut_S[11]));
 BUF_X1 output493 (.A(net495),
    .Z(dataOut_S[12]));
 BUF_X1 output494 (.A(net496),
    .Z(dataOut_S[13]));
 BUF_X1 output495 (.A(net497),
    .Z(dataOut_S[14]));
 BUF_X1 output496 (.A(net498),
    .Z(dataOut_S[15]));
 BUF_X1 output497 (.A(net499),
    .Z(dataOut_S[16]));
 BUF_X1 output498 (.A(net500),
    .Z(dataOut_S[17]));
 BUF_X1 output499 (.A(net501),
    .Z(dataOut_S[18]));
 BUF_X1 output500 (.A(net502),
    .Z(dataOut_S[19]));
 BUF_X1 output501 (.A(net503),
    .Z(dataOut_S[1]));
 BUF_X1 output502 (.A(net504),
    .Z(dataOut_S[20]));
 BUF_X1 output503 (.A(net505),
    .Z(dataOut_S[21]));
 BUF_X1 output504 (.A(net506),
    .Z(dataOut_S[22]));
 BUF_X1 output505 (.A(net507),
    .Z(dataOut_S[23]));
 BUF_X1 output506 (.A(net508),
    .Z(dataOut_S[24]));
 BUF_X1 output507 (.A(net509),
    .Z(dataOut_S[25]));
 BUF_X1 output508 (.A(net510),
    .Z(dataOut_S[26]));
 BUF_X1 output509 (.A(net511),
    .Z(dataOut_S[27]));
 BUF_X1 output510 (.A(net512),
    .Z(dataOut_S[28]));
 BUF_X1 output511 (.A(net513),
    .Z(dataOut_S[29]));
 BUF_X1 output512 (.A(net514),
    .Z(dataOut_S[2]));
 BUF_X1 output513 (.A(net515),
    .Z(dataOut_S[30]));
 BUF_X1 output514 (.A(net516),
    .Z(dataOut_S[31]));
 BUF_X1 output515 (.A(net517),
    .Z(dataOut_S[32]));
 BUF_X1 output516 (.A(net518),
    .Z(dataOut_S[33]));
 BUF_X1 output517 (.A(net519),
    .Z(dataOut_S[34]));
 BUF_X1 output518 (.A(net520),
    .Z(dataOut_S[35]));
 BUF_X1 output519 (.A(net521),
    .Z(dataOut_S[36]));
 BUF_X1 output520 (.A(net522),
    .Z(dataOut_S[37]));
 BUF_X1 output521 (.A(net523),
    .Z(dataOut_S[38]));
 BUF_X1 output522 (.A(net524),
    .Z(dataOut_S[39]));
 BUF_X1 output523 (.A(net525),
    .Z(dataOut_S[3]));
 BUF_X1 output524 (.A(net526),
    .Z(dataOut_S[40]));
 BUF_X1 output525 (.A(net527),
    .Z(dataOut_S[41]));
 BUF_X1 output526 (.A(net528),
    .Z(dataOut_S[42]));
 BUF_X1 output527 (.A(net529),
    .Z(dataOut_S[43]));
 BUF_X1 output528 (.A(net530),
    .Z(dataOut_S[44]));
 BUF_X1 output529 (.A(net531),
    .Z(dataOut_S[45]));
 BUF_X1 output530 (.A(net532),
    .Z(dataOut_S[46]));
 BUF_X1 output531 (.A(net533),
    .Z(dataOut_S[47]));
 BUF_X1 output532 (.A(net534),
    .Z(dataOut_S[48]));
 BUF_X1 output533 (.A(net535),
    .Z(dataOut_S[49]));
 BUF_X1 output534 (.A(net536),
    .Z(dataOut_S[4]));
 BUF_X1 output535 (.A(net537),
    .Z(dataOut_S[50]));
 BUF_X1 output536 (.A(net538),
    .Z(dataOut_S[51]));
 BUF_X1 output537 (.A(net539),
    .Z(dataOut_S[52]));
 BUF_X1 output538 (.A(net540),
    .Z(dataOut_S[53]));
 BUF_X1 output539 (.A(net541),
    .Z(dataOut_S[54]));
 BUF_X1 output540 (.A(net542),
    .Z(dataOut_S[55]));
 BUF_X1 output541 (.A(net543),
    .Z(dataOut_S[56]));
 BUF_X1 output542 (.A(net544),
    .Z(dataOut_S[57]));
 BUF_X1 output543 (.A(net545),
    .Z(dataOut_S[58]));
 BUF_X1 output544 (.A(net546),
    .Z(dataOut_S[59]));
 BUF_X1 output545 (.A(net547),
    .Z(dataOut_S[5]));
 BUF_X1 output546 (.A(net548),
    .Z(dataOut_S[60]));
 BUF_X1 output547 (.A(net549),
    .Z(dataOut_S[61]));
 BUF_X1 output548 (.A(net550),
    .Z(dataOut_S[62]));
 BUF_X1 output549 (.A(net551),
    .Z(dataOut_S[63]));
 BUF_X1 output550 (.A(net552),
    .Z(dataOut_S[6]));
 BUF_X1 output551 (.A(net553),
    .Z(dataOut_S[7]));
 BUF_X1 output552 (.A(net554),
    .Z(dataOut_S[8]));
 BUF_X1 output553 (.A(net555),
    .Z(dataOut_S[9]));
 BUF_X1 output554 (.A(net556),
    .Z(dataOut_W[0]));
 BUF_X1 output555 (.A(net557),
    .Z(dataOut_W[10]));
 BUF_X1 output556 (.A(net558),
    .Z(dataOut_W[11]));
 BUF_X1 output557 (.A(net559),
    .Z(dataOut_W[12]));
 BUF_X1 output558 (.A(net560),
    .Z(dataOut_W[13]));
 BUF_X1 output559 (.A(net561),
    .Z(dataOut_W[14]));
 BUF_X1 output560 (.A(net562),
    .Z(dataOut_W[15]));
 BUF_X1 output561 (.A(net563),
    .Z(dataOut_W[16]));
 BUF_X1 output562 (.A(net564),
    .Z(dataOut_W[17]));
 BUF_X1 output563 (.A(net565),
    .Z(dataOut_W[18]));
 BUF_X1 output564 (.A(net566),
    .Z(dataOut_W[19]));
 BUF_X1 output565 (.A(net567),
    .Z(dataOut_W[1]));
 BUF_X1 output566 (.A(net568),
    .Z(dataOut_W[20]));
 BUF_X1 output567 (.A(net569),
    .Z(dataOut_W[21]));
 BUF_X1 output568 (.A(net570),
    .Z(dataOut_W[22]));
 BUF_X1 output569 (.A(net571),
    .Z(dataOut_W[23]));
 BUF_X1 output570 (.A(net572),
    .Z(dataOut_W[24]));
 BUF_X1 output571 (.A(net573),
    .Z(dataOut_W[25]));
 BUF_X1 output572 (.A(net574),
    .Z(dataOut_W[26]));
 BUF_X1 output573 (.A(net575),
    .Z(dataOut_W[27]));
 BUF_X1 output574 (.A(net576),
    .Z(dataOut_W[28]));
 BUF_X1 output575 (.A(net577),
    .Z(dataOut_W[29]));
 BUF_X1 output576 (.A(net578),
    .Z(dataOut_W[2]));
 BUF_X1 output577 (.A(net579),
    .Z(dataOut_W[30]));
 BUF_X1 output578 (.A(net580),
    .Z(dataOut_W[31]));
 BUF_X1 output579 (.A(net581),
    .Z(dataOut_W[32]));
 BUF_X1 output580 (.A(net582),
    .Z(dataOut_W[33]));
 BUF_X1 output581 (.A(net583),
    .Z(dataOut_W[34]));
 BUF_X1 output582 (.A(net584),
    .Z(dataOut_W[35]));
 BUF_X1 output583 (.A(net585),
    .Z(dataOut_W[36]));
 BUF_X1 output584 (.A(net586),
    .Z(dataOut_W[37]));
 BUF_X1 output585 (.A(net587),
    .Z(dataOut_W[38]));
 BUF_X1 output586 (.A(net588),
    .Z(dataOut_W[39]));
 BUF_X1 output587 (.A(net589),
    .Z(dataOut_W[3]));
 BUF_X1 output588 (.A(net590),
    .Z(dataOut_W[40]));
 BUF_X1 output589 (.A(net591),
    .Z(dataOut_W[41]));
 BUF_X1 output590 (.A(net592),
    .Z(dataOut_W[42]));
 BUF_X1 output591 (.A(net593),
    .Z(dataOut_W[43]));
 BUF_X1 output592 (.A(net594),
    .Z(dataOut_W[44]));
 BUF_X1 output593 (.A(net595),
    .Z(dataOut_W[45]));
 BUF_X1 output594 (.A(net596),
    .Z(dataOut_W[46]));
 BUF_X1 output595 (.A(net597),
    .Z(dataOut_W[47]));
 BUF_X1 output596 (.A(net598),
    .Z(dataOut_W[48]));
 BUF_X1 output597 (.A(net599),
    .Z(dataOut_W[49]));
 BUF_X1 output598 (.A(net600),
    .Z(dataOut_W[4]));
 BUF_X1 output599 (.A(net601),
    .Z(dataOut_W[50]));
 BUF_X1 output600 (.A(net602),
    .Z(dataOut_W[51]));
 BUF_X1 output601 (.A(net603),
    .Z(dataOut_W[52]));
 BUF_X1 output602 (.A(net604),
    .Z(dataOut_W[53]));
 BUF_X1 output603 (.A(net605),
    .Z(dataOut_W[54]));
 BUF_X1 output604 (.A(net606),
    .Z(dataOut_W[55]));
 BUF_X1 output605 (.A(net607),
    .Z(dataOut_W[56]));
 BUF_X1 output606 (.A(net608),
    .Z(dataOut_W[57]));
 BUF_X1 output607 (.A(net609),
    .Z(dataOut_W[58]));
 BUF_X1 output608 (.A(net610),
    .Z(dataOut_W[59]));
 BUF_X1 output609 (.A(net611),
    .Z(dataOut_W[5]));
 BUF_X1 output610 (.A(net612),
    .Z(dataOut_W[60]));
 BUF_X1 output611 (.A(net613),
    .Z(dataOut_W[61]));
 BUF_X1 output612 (.A(net614),
    .Z(dataOut_W[62]));
 BUF_X1 output613 (.A(net615),
    .Z(dataOut_W[63]));
 BUF_X1 output614 (.A(net616),
    .Z(dataOut_W[6]));
 BUF_X1 output615 (.A(net617),
    .Z(dataOut_W[7]));
 BUF_X1 output616 (.A(net618),
    .Z(dataOut_W[8]));
 BUF_X1 output617 (.A(net619),
    .Z(dataOut_W[9]));
 BUF_X2 output618 (.A(net620),
    .Z(thanksIn_P));
 BUF_X1 output619 (.A(net621),
    .Z(validOut_E));
 BUF_X2 output620 (.A(net622),
    .Z(validOut_N));
 BUF_X1 output621 (.A(net623),
    .Z(validOut_P));
 BUF_X2 output622 (.A(net624),
    .Z(validOut_S));
 BUF_X2 output623 (.A(net756),
    .Z(validOut_W));
 BUF_X1 output624 (.A(net626),
    .Z(yummyOut_E));
 BUF_X1 output625 (.A(net627),
    .Z(yummyOut_N));
 BUF_X1 output626 (.A(net628),
    .Z(yummyOut_P));
 BUF_X1 output627 (.A(net629),
    .Z(yummyOut_S));
 BUF_X1 output628 (.A(net630),
    .Z(yummyOut_W));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_leaf_98_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_98_clk));
 CLKBUF_X3 clkbuf_leaf_99_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_99_clk));
 CLKBUF_X3 clkbuf_leaf_100_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_100_clk));
 CLKBUF_X3 clkbuf_leaf_101_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_101_clk));
 CLKBUF_X3 clkbuf_leaf_102_clk (.A(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_102_clk));
 CLKBUF_X3 clkbuf_leaf_103_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_103_clk));
 CLKBUF_X3 clkbuf_leaf_104_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_104_clk));
 CLKBUF_X3 clkbuf_leaf_105_clk (.A(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_105_clk));
 CLKBUF_X3 clkbuf_leaf_106_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_106_clk));
 CLKBUF_X3 clkbuf_leaf_107_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_107_clk));
 CLKBUF_X3 clkbuf_leaf_108_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_108_clk));
 CLKBUF_X3 clkbuf_leaf_109_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_109_clk));
 CLKBUF_X3 clkbuf_leaf_110_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_110_clk));
 CLKBUF_X3 clkbuf_leaf_111_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_111_clk));
 CLKBUF_X3 clkbuf_leaf_112_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_112_clk));
 CLKBUF_X3 clkbuf_leaf_113_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_113_clk));
 CLKBUF_X3 clkbuf_leaf_114_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_114_clk));
 CLKBUF_X3 clkbuf_leaf_115_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_115_clk));
 CLKBUF_X3 clkbuf_leaf_116_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_116_clk));
 CLKBUF_X3 clkbuf_leaf_117_clk (.A(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_117_clk));
 CLKBUF_X3 clkbuf_leaf_118_clk (.A(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_118_clk));
 CLKBUF_X3 clkbuf_leaf_119_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_119_clk));
 CLKBUF_X3 clkbuf_leaf_120_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_120_clk));
 CLKBUF_X3 clkbuf_leaf_121_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_121_clk));
 CLKBUF_X3 clkbuf_leaf_122_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_122_clk));
 CLKBUF_X3 clkbuf_leaf_123_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_123_clk));
 CLKBUF_X3 clkbuf_leaf_124_clk (.A(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_124_clk));
 CLKBUF_X3 clkbuf_leaf_125_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_125_clk));
 CLKBUF_X3 clkbuf_leaf_126_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_126_clk));
 CLKBUF_X3 clkbuf_leaf_127_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_127_clk));
 CLKBUF_X3 clkbuf_leaf_128_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_128_clk));
 CLKBUF_X3 clkbuf_leaf_129_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_129_clk));
 CLKBUF_X3 clkbuf_leaf_130_clk (.A(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_130_clk));
 CLKBUF_X3 clkbuf_leaf_131_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_131_clk));
 CLKBUF_X3 clkbuf_leaf_132_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_132_clk));
 CLKBUF_X3 clkbuf_leaf_133_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_133_clk));
 CLKBUF_X3 clkbuf_leaf_134_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_134_clk));
 CLKBUF_X3 clkbuf_leaf_135_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_135_clk));
 CLKBUF_X3 clkbuf_leaf_136_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_136_clk));
 CLKBUF_X3 clkbuf_leaf_137_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_137_clk));
 CLKBUF_X3 clkbuf_leaf_138_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_138_clk));
 CLKBUF_X3 clkbuf_leaf_139_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_139_clk));
 CLKBUF_X3 clkbuf_leaf_140_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_140_clk));
 CLKBUF_X3 clkbuf_leaf_141_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_141_clk));
 CLKBUF_X3 clkbuf_leaf_142_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_142_clk));
 CLKBUF_X3 clkbuf_leaf_143_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_143_clk));
 CLKBUF_X3 clkbuf_leaf_144_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_144_clk));
 CLKBUF_X3 clkbuf_leaf_145_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_145_clk));
 CLKBUF_X3 clkbuf_leaf_146_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_146_clk));
 CLKBUF_X3 clkbuf_leaf_147_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_147_clk));
 CLKBUF_X3 clkbuf_leaf_148_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_148_clk));
 CLKBUF_X3 clkbuf_leaf_149_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_149_clk));
 CLKBUF_X3 clkbuf_leaf_150_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_150_clk));
 CLKBUF_X3 clkbuf_leaf_151_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_151_clk));
 CLKBUF_X3 clkbuf_leaf_152_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_152_clk));
 CLKBUF_X3 clkbuf_leaf_153_clk (.A(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_153_clk));
 CLKBUF_X3 clkbuf_leaf_154_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_154_clk));
 CLKBUF_X3 clkbuf_leaf_155_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_155_clk));
 CLKBUF_X3 clkbuf_leaf_156_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_156_clk));
 CLKBUF_X3 clkbuf_leaf_157_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_157_clk));
 CLKBUF_X3 clkbuf_leaf_158_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_158_clk));
 CLKBUF_X3 clkbuf_leaf_159_clk (.A(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_159_clk));
 CLKBUF_X3 clkbuf_leaf_160_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_160_clk));
 CLKBUF_X3 clkbuf_leaf_161_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_161_clk));
 CLKBUF_X3 clkbuf_leaf_162_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_162_clk));
 CLKBUF_X3 clkbuf_leaf_163_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_163_clk));
 CLKBUF_X3 clkbuf_leaf_164_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_164_clk));
 CLKBUF_X3 clkbuf_leaf_165_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_165_clk));
 CLKBUF_X3 clkbuf_leaf_166_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_166_clk));
 CLKBUF_X3 clkbuf_leaf_167_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_167_clk));
 CLKBUF_X3 clkbuf_leaf_168_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_168_clk));
 CLKBUF_X3 clkbuf_leaf_169_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_169_clk));
 CLKBUF_X3 clkbuf_leaf_170_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_170_clk));
 CLKBUF_X3 clkbuf_leaf_171_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_171_clk));
 CLKBUF_X3 clkbuf_leaf_172_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_172_clk));
 CLKBUF_X3 clkbuf_leaf_173_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_173_clk));
 CLKBUF_X3 clkbuf_leaf_174_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_174_clk));
 CLKBUF_X3 clkbuf_leaf_175_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_175_clk));
 CLKBUF_X3 clkbuf_leaf_176_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_176_clk));
 CLKBUF_X3 clkbuf_leaf_177_clk (.A(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_177_clk));
 CLKBUF_X3 clkbuf_leaf_178_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_178_clk));
 CLKBUF_X3 clkbuf_leaf_179_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_179_clk));
 CLKBUF_X3 clkbuf_leaf_180_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_180_clk));
 CLKBUF_X3 clkbuf_leaf_181_clk (.A(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_181_clk));
 CLKBUF_X3 clkbuf_leaf_182_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_182_clk));
 CLKBUF_X3 clkbuf_leaf_183_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_183_clk));
 CLKBUF_X3 clkbuf_leaf_184_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_184_clk));
 CLKBUF_X3 clkbuf_leaf_185_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_185_clk));
 CLKBUF_X3 clkbuf_leaf_186_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_186_clk));
 CLKBUF_X3 clkbuf_leaf_187_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_187_clk));
 CLKBUF_X3 clkbuf_leaf_188_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_188_clk));
 CLKBUF_X3 clkbuf_leaf_189_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_189_clk));
 CLKBUF_X3 clkbuf_leaf_190_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_190_clk));
 CLKBUF_X3 clkbuf_leaf_191_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_191_clk));
 CLKBUF_X3 clkbuf_leaf_192_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_192_clk));
 CLKBUF_X3 clkbuf_leaf_193_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_193_clk));
 CLKBUF_X3 clkbuf_leaf_194_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_194_clk));
 CLKBUF_X3 clkbuf_leaf_195_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_195_clk));
 CLKBUF_X3 clkbuf_leaf_196_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_196_clk));
 CLKBUF_X3 clkbuf_leaf_197_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_197_clk));
 CLKBUF_X3 clkbuf_leaf_198_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_198_clk));
 CLKBUF_X3 clkbuf_leaf_199_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_199_clk));
 CLKBUF_X3 clkbuf_leaf_200_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_200_clk));
 CLKBUF_X3 clkbuf_leaf_201_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_201_clk));
 CLKBUF_X3 clkbuf_leaf_202_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_202_clk));
 CLKBUF_X3 clkbuf_leaf_203_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_203_clk));
 CLKBUF_X3 clkbuf_leaf_204_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_204_clk));
 CLKBUF_X3 clkbuf_leaf_205_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_205_clk));
 CLKBUF_X3 clkbuf_leaf_206_clk (.A(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_206_clk));
 CLKBUF_X3 clkbuf_leaf_207_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_207_clk));
 CLKBUF_X3 clkbuf_leaf_208_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_208_clk));
 CLKBUF_X3 clkbuf_leaf_209_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_209_clk));
 CLKBUF_X3 clkbuf_leaf_210_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_210_clk));
 CLKBUF_X3 clkbuf_leaf_211_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_211_clk));
 CLKBUF_X3 clkbuf_leaf_212_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_212_clk));
 CLKBUF_X3 clkbuf_leaf_213_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_213_clk));
 CLKBUF_X3 clkbuf_leaf_214_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_214_clk));
 CLKBUF_X3 clkbuf_leaf_215_clk (.A(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_215_clk));
 CLKBUF_X3 clkbuf_leaf_216_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_216_clk));
 CLKBUF_X3 clkbuf_leaf_217_clk (.A(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_217_clk));
 CLKBUF_X3 clkbuf_leaf_218_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_218_clk));
 CLKBUF_X3 clkbuf_leaf_219_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_219_clk));
 CLKBUF_X3 clkbuf_leaf_220_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_220_clk));
 CLKBUF_X3 clkbuf_leaf_221_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_221_clk));
 CLKBUF_X3 clkbuf_leaf_222_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_222_clk));
 CLKBUF_X3 clkbuf_leaf_223_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_223_clk));
 CLKBUF_X3 clkbuf_leaf_224_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_224_clk));
 CLKBUF_X3 clkbuf_leaf_225_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_225_clk));
 CLKBUF_X3 clkbuf_leaf_226_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_226_clk));
 CLKBUF_X3 clkbuf_leaf_227_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_227_clk));
 CLKBUF_X3 clkbuf_leaf_228_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_228_clk));
 CLKBUF_X3 clkbuf_leaf_229_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_229_clk));
 CLKBUF_X3 clkbuf_leaf_230_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_230_clk));
 CLKBUF_X3 clkbuf_leaf_231_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_231_clk));
 CLKBUF_X3 clkbuf_leaf_232_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_232_clk));
 CLKBUF_X3 clkbuf_leaf_233_clk (.A(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_233_clk));
 CLKBUF_X3 clkbuf_leaf_234_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_234_clk));
 CLKBUF_X3 clkbuf_leaf_235_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_235_clk));
 CLKBUF_X3 clkbuf_leaf_236_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_236_clk));
 CLKBUF_X3 clkbuf_leaf_237_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_237_clk));
 CLKBUF_X3 clkbuf_leaf_238_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_238_clk));
 CLKBUF_X3 clkbuf_leaf_239_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_239_clk));
 CLKBUF_X3 clkbuf_leaf_240_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_240_clk));
 CLKBUF_X3 clkbuf_leaf_241_clk (.A(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_241_clk));
 CLKBUF_X3 clkbuf_leaf_242_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_242_clk));
 CLKBUF_X3 clkbuf_leaf_243_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_243_clk));
 CLKBUF_X3 clkbuf_leaf_244_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_244_clk));
 CLKBUF_X3 clkbuf_leaf_245_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_245_clk));
 CLKBUF_X3 clkbuf_leaf_246_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_246_clk));
 CLKBUF_X3 clkbuf_leaf_247_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_247_clk));
 CLKBUF_X3 clkbuf_leaf_248_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_248_clk));
 CLKBUF_X3 clkbuf_leaf_249_clk (.A(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_249_clk));
 CLKBUF_X3 clkbuf_leaf_250_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_250_clk));
 CLKBUF_X3 clkbuf_leaf_251_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_251_clk));
 CLKBUF_X3 clkbuf_leaf_252_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_252_clk));
 CLKBUF_X3 clkbuf_leaf_253_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_253_clk));
 CLKBUF_X3 clkbuf_leaf_254_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_254_clk));
 CLKBUF_X3 clkbuf_leaf_255_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_255_clk));
 CLKBUF_X3 clkbuf_leaf_256_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_256_clk));
 CLKBUF_X3 clkbuf_leaf_257_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_257_clk));
 CLKBUF_X3 clkbuf_leaf_258_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_258_clk));
 CLKBUF_X3 clkbuf_leaf_259_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_259_clk));
 CLKBUF_X3 clkbuf_leaf_260_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_260_clk));
 CLKBUF_X3 clkbuf_leaf_261_clk (.A(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_261_clk));
 CLKBUF_X3 clkbuf_leaf_262_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_262_clk));
 CLKBUF_X3 clkbuf_leaf_263_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_263_clk));
 CLKBUF_X3 clkbuf_leaf_264_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_264_clk));
 CLKBUF_X3 clkbuf_leaf_265_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_265_clk));
 CLKBUF_X3 clkbuf_leaf_266_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_266_clk));
 CLKBUF_X3 clkbuf_leaf_267_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_267_clk));
 CLKBUF_X3 clkbuf_leaf_268_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_268_clk));
 CLKBUF_X3 clkbuf_leaf_269_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_269_clk));
 CLKBUF_X3 clkbuf_leaf_270_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_270_clk));
 CLKBUF_X3 clkbuf_leaf_271_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_271_clk));
 CLKBUF_X3 clkbuf_leaf_272_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_272_clk));
 CLKBUF_X3 clkbuf_leaf_273_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_273_clk));
 CLKBUF_X3 clkbuf_leaf_274_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_274_clk));
 CLKBUF_X3 clkbuf_leaf_275_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_275_clk));
 CLKBUF_X3 clkbuf_leaf_276_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_276_clk));
 CLKBUF_X3 clkbuf_leaf_277_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_277_clk));
 CLKBUF_X3 clkbuf_leaf_278_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_278_clk));
 CLKBUF_X3 clkbuf_leaf_279_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_279_clk));
 CLKBUF_X3 clkbuf_leaf_280_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_280_clk));
 CLKBUF_X3 clkbuf_leaf_281_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_281_clk));
 CLKBUF_X3 clkbuf_leaf_282_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_282_clk));
 CLKBUF_X3 clkbuf_leaf_283_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_283_clk));
 CLKBUF_X3 clkbuf_leaf_284_clk (.A(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_284_clk));
 CLKBUF_X3 clkbuf_leaf_285_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_285_clk));
 CLKBUF_X3 clkbuf_leaf_286_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_286_clk));
 CLKBUF_X3 clkbuf_leaf_287_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_287_clk));
 CLKBUF_X3 clkbuf_leaf_288_clk (.A(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_288_clk));
 CLKBUF_X3 clkbuf_leaf_289_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_289_clk));
 CLKBUF_X3 clkbuf_leaf_290_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_290_clk));
 CLKBUF_X3 clkbuf_leaf_291_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_291_clk));
 CLKBUF_X3 clkbuf_leaf_292_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_292_clk));
 CLKBUF_X3 clkbuf_leaf_293_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_293_clk));
 CLKBUF_X3 clkbuf_leaf_294_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_294_clk));
 CLKBUF_X3 clkbuf_leaf_295_clk (.A(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_295_clk));
 CLKBUF_X3 clkbuf_leaf_296_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_296_clk));
 CLKBUF_X3 clkbuf_leaf_297_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_297_clk));
 CLKBUF_X3 clkbuf_leaf_298_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_298_clk));
 CLKBUF_X3 clkbuf_leaf_299_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_299_clk));
 CLKBUF_X3 clkbuf_leaf_300_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_300_clk));
 CLKBUF_X3 clkbuf_leaf_301_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_301_clk));
 CLKBUF_X3 clkbuf_leaf_302_clk (.A(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_302_clk));
 CLKBUF_X3 clkbuf_leaf_303_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_303_clk));
 CLKBUF_X3 clkbuf_leaf_304_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_304_clk));
 CLKBUF_X3 clkbuf_leaf_305_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_305_clk));
 CLKBUF_X3 clkbuf_leaf_306_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_306_clk));
 CLKBUF_X3 clkbuf_leaf_307_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_307_clk));
 CLKBUF_X3 clkbuf_leaf_308_clk (.A(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_308_clk));
 CLKBUF_X3 clkbuf_leaf_309_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_309_clk));
 CLKBUF_X3 clkbuf_leaf_310_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_310_clk));
 CLKBUF_X3 clkbuf_leaf_311_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_311_clk));
 CLKBUF_X3 clkbuf_leaf_312_clk (.A(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_312_clk));
 CLKBUF_X3 clkbuf_leaf_313_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_313_clk));
 CLKBUF_X3 clkbuf_leaf_314_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_314_clk));
 CLKBUF_X3 clkbuf_leaf_315_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_315_clk));
 CLKBUF_X3 clkbuf_leaf_316_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_316_clk));
 CLKBUF_X3 clkbuf_leaf_317_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_317_clk));
 CLKBUF_X3 clkbuf_leaf_318_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_318_clk));
 CLKBUF_X3 clkbuf_leaf_319_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_319_clk));
 CLKBUF_X3 clkbuf_leaf_320_clk (.A(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_320_clk));
 CLKBUF_X3 clkbuf_leaf_321_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_321_clk));
 CLKBUF_X3 clkbuf_leaf_322_clk (.A(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_322_clk));
 CLKBUF_X3 clkbuf_leaf_323_clk (.A(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_323_clk));
 CLKBUF_X3 clkbuf_leaf_324_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_324_clk));
 CLKBUF_X3 clkbuf_leaf_325_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_325_clk));
 CLKBUF_X3 clkbuf_leaf_326_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_326_clk));
 CLKBUF_X3 clkbuf_leaf_327_clk (.A(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_327_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 CLKBUF_X3 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_5_0__leaf_clk));
 CLKBUF_X3 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_5_1__leaf_clk));
 CLKBUF_X3 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_5_2__leaf_clk));
 CLKBUF_X3 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_5_3__leaf_clk));
 CLKBUF_X3 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_5_4__leaf_clk));
 CLKBUF_X3 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_5_5__leaf_clk));
 CLKBUF_X3 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_5_6__leaf_clk));
 CLKBUF_X3 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_5_7__leaf_clk));
 CLKBUF_X3 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_5_8__leaf_clk));
 CLKBUF_X3 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_5_9__leaf_clk));
 CLKBUF_X3 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_5_10__leaf_clk));
 CLKBUF_X3 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_5_11__leaf_clk));
 CLKBUF_X3 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_5_12__leaf_clk));
 CLKBUF_X3 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_5_13__leaf_clk));
 CLKBUF_X3 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_5_14__leaf_clk));
 CLKBUF_X3 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_5_15__leaf_clk));
 CLKBUF_X3 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_5_16__leaf_clk));
 CLKBUF_X3 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_5_17__leaf_clk));
 CLKBUF_X3 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_5_18__leaf_clk));
 CLKBUF_X3 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_5_19__leaf_clk));
 CLKBUF_X3 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_5_20__leaf_clk));
 CLKBUF_X3 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_5_21__leaf_clk));
 CLKBUF_X3 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_5_22__leaf_clk));
 CLKBUF_X3 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_5_23__leaf_clk));
 CLKBUF_X3 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_5_24__leaf_clk));
 CLKBUF_X3 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_5_25__leaf_clk));
 CLKBUF_X3 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_5_26__leaf_clk));
 CLKBUF_X3 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_5_27__leaf_clk));
 CLKBUF_X3 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_5_28__leaf_clk));
 CLKBUF_X3 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_5_29__leaf_clk));
 CLKBUF_X3 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_5_30__leaf_clk));
 CLKBUF_X3 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_5_31__leaf_clk));
 INV_X2 clkload0 (.A(clknet_5_1__leaf_clk));
 CLKBUF_X3 clkload1 (.A(clknet_5_7__leaf_clk));
 CLKBUF_X3 clkload2 (.A(clknet_5_8__leaf_clk));
 CLKBUF_X3 clkload3 (.A(clknet_5_10__leaf_clk));
 INV_X4 clkload4 (.A(clknet_5_13__leaf_clk));
 CLKBUF_X3 clkload5 (.A(clknet_5_15__leaf_clk));
 CLKBUF_X3 clkload6 (.A(clknet_5_16__leaf_clk));
 INV_X4 clkload7 (.A(clknet_5_19__leaf_clk));
 INV_X4 clkload8 (.A(clknet_5_21__leaf_clk));
 INV_X4 clkload9 (.A(clknet_5_25__leaf_clk));
 INV_X2 clkload10 (.A(clknet_5_27__leaf_clk));
 INV_X2 clkload11 (.A(clknet_5_28__leaf_clk));
 INV_X2 clkload12 (.A(clknet_5_30__leaf_clk));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_9_clk));
 CLKBUF_X1 clkload14 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload15 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_13_clk));
 INV_X1 clkload17 (.A(clknet_leaf_324_clk));
 INV_X1 clkload18 (.A(clknet_leaf_325_clk));
 CLKBUF_X1 clkload19 (.A(clknet_leaf_326_clk));
 CLKBUF_X1 clkload20 (.A(clknet_leaf_327_clk));
 CLKBUF_X1 clkload21 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_2_clk));
 INV_X1 clkload23 (.A(clknet_leaf_3_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_5_clk));
 INV_X1 clkload25 (.A(clknet_leaf_6_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_8_clk));
 CLKBUF_X1 clkload27 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_323_clk));
 INV_X1 clkload29 (.A(clknet_leaf_17_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_18_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_21_clk));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_76_clk));
 CLKBUF_X1 clkload35 (.A(clknet_leaf_77_clk));
 INV_X1 clkload36 (.A(clknet_leaf_23_clk));
 CLKBUF_X1 clkload37 (.A(clknet_leaf_24_clk));
 INV_X1 clkload38 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload39 (.A(clknet_leaf_29_clk));
 INV_X1 clkload40 (.A(clknet_leaf_30_clk));
 INV_X1 clkload41 (.A(clknet_leaf_31_clk));
 INV_X1 clkload42 (.A(clknet_leaf_71_clk));
 INV_X1 clkload43 (.A(clknet_leaf_72_clk));
 CLKBUF_X1 clkload44 (.A(clknet_leaf_4_clk));
 CLKBUF_X1 clkload45 (.A(clknet_leaf_317_clk));
 CLKBUF_X1 clkload46 (.A(clknet_leaf_321_clk));
 INV_X1 clkload47 (.A(clknet_leaf_322_clk));
 CLKBUF_X1 clkload48 (.A(clknet_leaf_310_clk));
 CLKBUF_X1 clkload49 (.A(clknet_leaf_311_clk));
 CLKBUF_X1 clkload50 (.A(clknet_leaf_314_clk));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_318_clk));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_319_clk));
 INV_X1 clkload53 (.A(clknet_leaf_320_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_36_clk));
 CLKBUF_X1 clkload55 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload56 (.A(clknet_leaf_40_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_45_clk));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_44_clk));
 INV_X1 clkload59 (.A(clknet_leaf_46_clk));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_47_clk));
 INV_X1 clkload61 (.A(clknet_leaf_48_clk));
 CLKBUF_X1 clkload62 (.A(clknet_leaf_49_clk));
 INV_X1 clkload63 (.A(clknet_leaf_305_clk));
 CLKBUF_X1 clkload64 (.A(clknet_leaf_306_clk));
 CLKBUF_X1 clkload65 (.A(clknet_leaf_307_clk));
 INV_X2 clkload66 (.A(clknet_leaf_78_clk));
 INV_X1 clkload67 (.A(clknet_leaf_79_clk));
 INV_X1 clkload68 (.A(clknet_leaf_80_clk));
 CLKBUF_X1 clkload69 (.A(clknet_leaf_81_clk));
 INV_X2 clkload70 (.A(clknet_leaf_82_clk));
 INV_X1 clkload71 (.A(clknet_leaf_83_clk));
 INV_X1 clkload72 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload73 (.A(clknet_leaf_68_clk));
 CLKBUF_X1 clkload74 (.A(clknet_leaf_73_clk));
 INV_X1 clkload75 (.A(clknet_leaf_74_clk));
 INV_X1 clkload76 (.A(clknet_leaf_75_clk));
 CLKBUF_X1 clkload77 (.A(clknet_leaf_88_clk));
 INV_X1 clkload78 (.A(clknet_leaf_89_clk));
 INV_X1 clkload79 (.A(clknet_leaf_86_clk));
 CLKBUF_X1 clkload80 (.A(clknet_leaf_98_clk));
 CLKBUF_X1 clkload81 (.A(clknet_leaf_90_clk));
 INV_X1 clkload82 (.A(clknet_leaf_91_clk));
 INV_X2 clkload83 (.A(clknet_leaf_92_clk));
 INV_X1 clkload84 (.A(clknet_leaf_93_clk));
 INV_X1 clkload85 (.A(clknet_leaf_94_clk));
 CLKBUF_X1 clkload86 (.A(clknet_leaf_95_clk));
 INV_X1 clkload87 (.A(clknet_leaf_97_clk));
 INV_X2 clkload88 (.A(clknet_leaf_103_clk));
 INV_X1 clkload89 (.A(clknet_leaf_104_clk));
 CLKBUF_X1 clkload90 (.A(clknet_leaf_55_clk));
 CLKBUF_X1 clkload91 (.A(clknet_leaf_56_clk));
 CLKBUF_X1 clkload92 (.A(clknet_leaf_57_clk));
 INV_X1 clkload93 (.A(clknet_leaf_60_clk));
 CLKBUF_X1 clkload94 (.A(clknet_leaf_118_clk));
 INV_X2 clkload95 (.A(clknet_leaf_50_clk));
 INV_X1 clkload96 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload97 (.A(clknet_leaf_119_clk));
 CLKBUF_X1 clkload98 (.A(clknet_leaf_126_clk));
 INV_X1 clkload99 (.A(clknet_leaf_128_clk));
 INV_X1 clkload100 (.A(clknet_leaf_129_clk));
 CLKBUF_X1 clkload101 (.A(clknet_leaf_62_clk));
 CLKBUF_X1 clkload102 (.A(clknet_leaf_63_clk));
 CLKBUF_X1 clkload103 (.A(clknet_leaf_107_clk));
 CLKBUF_X1 clkload104 (.A(clknet_leaf_112_clk));
 INV_X1 clkload105 (.A(clknet_leaf_114_clk));
 CLKBUF_X1 clkload106 (.A(clknet_leaf_115_clk));
 INV_X1 clkload107 (.A(clknet_leaf_116_clk));
 CLKBUF_X1 clkload108 (.A(clknet_leaf_117_clk));
 INV_X1 clkload109 (.A(clknet_leaf_108_clk));
 CLKBUF_X1 clkload110 (.A(clknet_leaf_109_clk));
 INV_X1 clkload111 (.A(clknet_leaf_111_clk));
 CLKBUF_X1 clkload112 (.A(clknet_leaf_121_clk));
 CLKBUF_X1 clkload113 (.A(clknet_leaf_124_clk));
 INV_X1 clkload114 (.A(clknet_leaf_271_clk));
 CLKBUF_X1 clkload115 (.A(clknet_leaf_274_clk));
 CLKBUF_X1 clkload116 (.A(clknet_leaf_275_clk));
 CLKBUF_X1 clkload117 (.A(clknet_leaf_276_clk));
 CLKBUF_X1 clkload118 (.A(clknet_leaf_277_clk));
 CLKBUF_X1 clkload119 (.A(clknet_leaf_278_clk));
 CLKBUF_X1 clkload120 (.A(clknet_leaf_284_clk));
 INV_X1 clkload121 (.A(clknet_leaf_262_clk));
 INV_X1 clkload122 (.A(clknet_leaf_263_clk));
 INV_X1 clkload123 (.A(clknet_leaf_264_clk));
 INV_X1 clkload124 (.A(clknet_leaf_265_clk));
 INV_X1 clkload125 (.A(clknet_leaf_266_clk));
 INV_X1 clkload126 (.A(clknet_leaf_268_clk));
 INV_X2 clkload127 (.A(clknet_leaf_269_clk));
 INV_X1 clkload128 (.A(clknet_leaf_270_clk));
 INV_X2 clkload129 (.A(clknet_leaf_285_clk));
 INV_X2 clkload130 (.A(clknet_leaf_286_clk));
 INV_X1 clkload131 (.A(clknet_leaf_288_clk));
 INV_X1 clkload132 (.A(clknet_leaf_204_clk));
 CLKBUF_X1 clkload133 (.A(clknet_leaf_282_clk));
 INV_X1 clkload134 (.A(clknet_leaf_294_clk));
 CLKBUF_X1 clkload135 (.A(clknet_leaf_296_clk));
 CLKBUF_X1 clkload136 (.A(clknet_leaf_298_clk));
 CLKBUF_X1 clkload137 (.A(clknet_leaf_300_clk));
 INV_X1 clkload138 (.A(clknet_leaf_301_clk));
 CLKBUF_X1 clkload139 (.A(clknet_leaf_303_clk));
 INV_X1 clkload140 (.A(clknet_leaf_304_clk));
 CLKBUF_X1 clkload141 (.A(clknet_leaf_308_clk));
 CLKBUF_X1 clkload142 (.A(clknet_leaf_205_clk));
 CLKBUF_X1 clkload143 (.A(clknet_leaf_287_clk));
 CLKBUF_X1 clkload144 (.A(clknet_leaf_289_clk));
 INV_X1 clkload145 (.A(clknet_leaf_290_clk));
 INV_X1 clkload146 (.A(clknet_leaf_293_clk));
 CLKBUF_X1 clkload147 (.A(clknet_leaf_234_clk));
 INV_X1 clkload148 (.A(clknet_leaf_235_clk));
 INV_X1 clkload149 (.A(clknet_leaf_237_clk));
 CLKBUF_X1 clkload150 (.A(clknet_leaf_250_clk));
 CLKBUF_X1 clkload151 (.A(clknet_leaf_252_clk));
 CLKBUF_X1 clkload152 (.A(clknet_leaf_253_clk));
 INV_X1 clkload153 (.A(clknet_leaf_254_clk));
 CLKBUF_X1 clkload154 (.A(clknet_leaf_255_clk));
 CLKBUF_X1 clkload155 (.A(clknet_leaf_256_clk));
 CLKBUF_X1 clkload156 (.A(clknet_leaf_258_clk));
 CLKBUF_X1 clkload157 (.A(clknet_leaf_259_clk));
 CLKBUF_X1 clkload158 (.A(clknet_leaf_236_clk));
 CLKBUF_X1 clkload159 (.A(clknet_leaf_243_clk));
 INV_X2 clkload160 (.A(clknet_leaf_246_clk));
 CLKBUF_X1 clkload161 (.A(clknet_leaf_247_clk));
 CLKBUF_X1 clkload162 (.A(clknet_leaf_248_clk));
 INV_X1 clkload163 (.A(clknet_leaf_249_clk));
 CLKBUF_X1 clkload164 (.A(clknet_leaf_207_clk));
 CLKBUF_X1 clkload165 (.A(clknet_leaf_208_clk));
 CLKBUF_X1 clkload166 (.A(clknet_leaf_209_clk));
 INV_X1 clkload167 (.A(clknet_leaf_210_clk));
 CLKBUF_X1 clkload168 (.A(clknet_leaf_212_clk));
 CLKBUF_X1 clkload169 (.A(clknet_leaf_213_clk));
 CLKBUF_X1 clkload170 (.A(clknet_leaf_214_clk));
 INV_X1 clkload171 (.A(clknet_leaf_221_clk));
 CLKBUF_X1 clkload172 (.A(clknet_leaf_222_clk));
 CLKBUF_X1 clkload173 (.A(clknet_leaf_230_clk));
 CLKBUF_X1 clkload174 (.A(clknet_leaf_231_clk));
 CLKBUF_X1 clkload175 (.A(clknet_leaf_232_clk));
 CLKBUF_X1 clkload176 (.A(clknet_leaf_218_clk));
 CLKBUF_X1 clkload177 (.A(clknet_leaf_223_clk));
 CLKBUF_X1 clkload178 (.A(clknet_leaf_224_clk));
 CLKBUF_X1 clkload179 (.A(clknet_leaf_225_clk));
 INV_X1 clkload180 (.A(clknet_leaf_228_clk));
 INV_X1 clkload181 (.A(clknet_leaf_229_clk));
 CLKBUF_X1 clkload182 (.A(clknet_leaf_239_clk));
 CLKBUF_X1 clkload183 (.A(clknet_leaf_240_clk));
 CLKBUF_X1 clkload184 (.A(clknet_leaf_131_clk));
 CLKBUF_X1 clkload185 (.A(clknet_leaf_132_clk));
 CLKBUF_X1 clkload186 (.A(clknet_leaf_133_clk));
 CLKBUF_X1 clkload187 (.A(clknet_leaf_134_clk));
 CLKBUF_X1 clkload188 (.A(clknet_leaf_135_clk));
 CLKBUF_X1 clkload189 (.A(clknet_leaf_136_clk));
 INV_X1 clkload190 (.A(clknet_leaf_139_clk));
 CLKBUF_X1 clkload191 (.A(clknet_leaf_201_clk));
 CLKBUF_X1 clkload192 (.A(clknet_leaf_202_clk));
 INV_X1 clkload193 (.A(clknet_leaf_302_clk));
 INV_X2 clkload194 (.A(clknet_leaf_196_clk));
 CLKBUF_X1 clkload195 (.A(clknet_leaf_198_clk));
 INV_X1 clkload196 (.A(clknet_leaf_199_clk));
 CLKBUF_X1 clkload197 (.A(clknet_leaf_203_clk));
 INV_X2 clkload198 (.A(clknet_leaf_206_clk));
 CLKBUF_X1 clkload199 (.A(clknet_leaf_138_clk));
 CLKBUF_X1 clkload200 (.A(clknet_leaf_144_clk));
 INV_X1 clkload201 (.A(clknet_leaf_145_clk));
 CLKBUF_X1 clkload202 (.A(clknet_leaf_147_clk));
 CLKBUF_X1 clkload203 (.A(clknet_leaf_149_clk));
 INV_X1 clkload204 (.A(clknet_leaf_150_clk));
 INV_X1 clkload205 (.A(clknet_leaf_151_clk));
 CLKBUF_X1 clkload206 (.A(clknet_leaf_152_clk));
 CLKBUF_X1 clkload207 (.A(clknet_leaf_153_clk));
 INV_X2 clkload208 (.A(clknet_leaf_140_clk));
 CLKBUF_X1 clkload209 (.A(clknet_leaf_141_clk));
 CLKBUF_X1 clkload210 (.A(clknet_leaf_142_clk));
 INV_X1 clkload211 (.A(clknet_leaf_143_clk));
 CLKBUF_X1 clkload212 (.A(clknet_leaf_155_clk));
 CLKBUF_X1 clkload213 (.A(clknet_leaf_156_clk));
 INV_X1 clkload214 (.A(clknet_leaf_157_clk));
 CLKBUF_X1 clkload215 (.A(clknet_leaf_158_clk));
 CLKBUF_X1 clkload216 (.A(clknet_leaf_159_clk));
 CLKBUF_X1 clkload217 (.A(clknet_leaf_190_clk));
 INV_X2 clkload218 (.A(clknet_leaf_195_clk));
 INV_X1 clkload219 (.A(clknet_leaf_178_clk));
 CLKBUF_X1 clkload220 (.A(clknet_leaf_182_clk));
 CLKBUF_X1 clkload221 (.A(clknet_leaf_183_clk));
 INV_X1 clkload222 (.A(clknet_leaf_185_clk));
 CLKBUF_X1 clkload223 (.A(clknet_leaf_186_clk));
 CLKBUF_X1 clkload224 (.A(clknet_leaf_187_clk));
 CLKBUF_X1 clkload225 (.A(clknet_leaf_188_clk));
 CLKBUF_X1 clkload226 (.A(clknet_leaf_189_clk));
 CLKBUF_X1 clkload227 (.A(clknet_leaf_216_clk));
 CLKBUF_X1 clkload228 (.A(clknet_leaf_217_clk));
 INV_X1 clkload229 (.A(clknet_leaf_160_clk));
 CLKBUF_X1 clkload230 (.A(clknet_leaf_162_clk));
 CLKBUF_X1 clkload231 (.A(clknet_leaf_163_clk));
 CLKBUF_X1 clkload232 (.A(clknet_leaf_164_clk));
 CLKBUF_X1 clkload233 (.A(clknet_leaf_175_clk));
 CLKBUF_X1 clkload234 (.A(clknet_leaf_176_clk));
 INV_X2 clkload235 (.A(clknet_leaf_177_clk));
 INV_X1 clkload236 (.A(clknet_leaf_166_clk));
 INV_X1 clkload237 (.A(clknet_leaf_167_clk));
 CLKBUF_X1 clkload238 (.A(clknet_leaf_168_clk));
 CLKBUF_X1 clkload239 (.A(clknet_leaf_169_clk));
 CLKBUF_X1 clkload240 (.A(clknet_leaf_170_clk));
 INV_X1 clkload241 (.A(clknet_leaf_171_clk));
 CLKBUF_X1 clkload242 (.A(clknet_leaf_172_clk));
 CLKBUF_X1 clkload243 (.A(clknet_leaf_173_clk));
 INV_X1 clkload244 (.A(clknet_leaf_174_clk));
 CLKBUF_X1 clkload245 (.A(clknet_leaf_180_clk));
 CLKBUF_X1 clkload246 (.A(clknet_leaf_181_clk));
 BUF_X1 rebuffer1 (.A(net691),
    .Z(net631));
 BUF_X1 rebuffer2 (.A(_10300_),
    .Z(net632));
 BUF_X1 rebuffer3 (.A(_10308_),
    .Z(net633));
 BUF_X1 rebuffer4 (.A(_10308_),
    .Z(net634));
 BUF_X1 rebuffer5 (.A(net661),
    .Z(net635));
 BUF_X1 rebuffer6 (.A(net635),
    .Z(net636));
 BUF_X1 rebuffer7 (.A(_10335_),
    .Z(net637));
 BUF_X1 rebuffer8 (.A(_10326_),
    .Z(net638));
 BUF_X1 rebuffer9 (.A(net638),
    .Z(net639));
 BUF_X1 rebuffer10 (.A(_10264_),
    .Z(net640));
 BUF_X1 rebuffer11 (.A(_10190_),
    .Z(net641));
 BUF_X1 rebuffer12 (.A(_10182_),
    .Z(net642));
 BUF_X1 rebuffer13 (.A(_10182_),
    .Z(net643));
 BUF_X1 rebuffer14 (.A(net643),
    .Z(net644));
 BUF_X1 rebuffer15 (.A(_10188_),
    .Z(net645));
 BUF_X1 rebuffer16 (.A(net645),
    .Z(net646));
 BUF_X1 rebuffer17 (.A(_10200_),
    .Z(net647));
 BUF_X1 rebuffer18 (.A(net647),
    .Z(net648));
 BUF_X1 rebuffer19 (.A(net692),
    .Z(net649));
 BUF_X1 rebuffer20 (.A(_10203_),
    .Z(net650));
 BUF_X1 rebuffer21 (.A(_07293_),
    .Z(net651));
 BUF_X1 rebuffer22 (.A(net651),
    .Z(net652));
 BUF_X1 rebuffer23 (.A(_10184_),
    .Z(net653));
 BUF_X1 rebuffer24 (.A(_10362_),
    .Z(net654));
 BUF_X1 rebuffer25 (.A(net654),
    .Z(net655));
 BUF_X1 rebuffer26 (.A(_10362_),
    .Z(net656));
 BUF_X1 rebuffer27 (.A(_10205_),
    .Z(net657));
 BUF_X1 rebuffer28 (.A(net696),
    .Z(net658));
 BUF_X1 rebuffer29 (.A(_10202_),
    .Z(net659));
 BUF_X1 rebuffer30 (.A(_10332_),
    .Z(net660));
 BUF_X2 rebuffer31 (.A(_10230_),
    .Z(net661));
 BUF_X1 rebuffer32 (.A(_00008_),
    .Z(net662));
 BUF_X1 rebuffer109 (.A(_00006_),
    .Z(net758));
 BUF_X1 rebuffer34 (.A(_07509_),
    .Z(net664));
 BUF_X1 rebuffer35 (.A(net664),
    .Z(net665));
 BUF_X1 rebuffer36 (.A(_05128_),
    .Z(net666));
 BUF_X2 clone37 (.A(_06120_),
    .Z(net667));
 BUF_X4 clone38 (.A(net669),
    .Z(net668));
 BUF_X1 rebuffer39 (.A(_00014_),
    .Z(net669));
 BUF_X1 rebuffer40 (.A(_10324_),
    .Z(net670));
 BUF_X2 rebuffer41 (.A(net670),
    .Z(net671));
 BUF_X1 rebuffer42 (.A(_00016_),
    .Z(net672));
 BUF_X1 rebuffer43 (.A(_07431_),
    .Z(net673));
 BUF_X1 rebuffer44 (.A(net673),
    .Z(net674));
 BUF_X1 rebuffer45 (.A(net674),
    .Z(net675));
 BUF_X1 rebuffer46 (.A(_10196_),
    .Z(net676));
 BUF_X1 rebuffer47 (.A(_05309_),
    .Z(net677));
 BUF_X1 rebuffer48 (.A(_05309_),
    .Z(net678));
 BUF_X1 rebuffer49 (.A(net733),
    .Z(net679));
 BUF_X4 clone50 (.A(net693),
    .Z(net680));
 BUF_X2 rebuffer51 (.A(_10314_),
    .Z(net681));
 BUF_X2 rebuffer52 (.A(net705),
    .Z(net682));
 BUF_X1 rebuffer53 (.A(net682),
    .Z(net683));
 BUF_X1 rebuffer54 (.A(net683),
    .Z(net684));
 BUF_X1 rebuffer55 (.A(_05138_),
    .Z(net685));
 BUF_X1 rebuffer56 (.A(_10197_),
    .Z(net686));
 BUF_X1 rebuffer57 (.A(_05129_),
    .Z(net687));
 BUF_X1 rebuffer58 (.A(_07479_),
    .Z(net688));
 BUF_X1 rebuffer59 (.A(net688),
    .Z(net689));
 BUF_X1 rebuffer60 (.A(net688),
    .Z(net690));
 BUF_X1 rebuffer68 (.A(_05455_),
    .Z(net698));
 BUF_X1 rebuffer69 (.A(_05455_),
    .Z(net699));
 BUF_X1 rebuffer70 (.A(_05455_),
    .Z(net700));
 BUF_X1 rebuffer71 (.A(net700),
    .Z(net701));
 BUF_X2 clone72 (.A(_05590_),
    .Z(net702));
 BUF_X1 rebuffer73 (.A(_10330_),
    .Z(net703));
 BUF_X1 rebuffer74 (.A(net703),
    .Z(net704));
 BUF_X1 rebuffer75 (.A(_05509_),
    .Z(net705));
 BUF_X16 clone115 (.A(_05129_),
    .Z(net765));
 BUF_X2 rebuffer114 (.A(_05129_),
    .Z(net764));
 BUF_X1 rebuffer78 (.A(net709),
    .Z(net708));
 BUF_X1 rebuffer79 (.A(net710),
    .Z(net709));
 BUF_X1 rebuffer80 (.A(net712),
    .Z(net710));
 BUF_X16 clone81 (.A(net714),
    .Z(net711));
 BUF_X2 rebuffer82 (.A(net758),
    .Z(net712));
 BUF_X1 rebuffer83 (.A(_10360_),
    .Z(net713));
 BUF_X1 rebuffer84 (.A(_05455_),
    .Z(net714));
 BUF_X1 rebuffer85 (.A(_10329_),
    .Z(net715));
 BUF_X1 rebuffer86 (.A(_10344_),
    .Z(net716));
 BUF_X16 clone87 (.A(net722),
    .Z(net717));
 BUF_X1 rebuffer88 (.A(_10353_),
    .Z(net718));
 BUF_X1 rebuffer89 (.A(_10356_),
    .Z(net719));
 BUF_X16 clone90 (.A(_05456_),
    .Z(net720));
 BUF_X16 clone91 (.A(_05458_),
    .Z(net721));
 BUF_X8 rebuffer92 (.A(_05455_),
    .Z(net722));
 BUF_X1 rebuffer93 (.A(_10339_),
    .Z(net723));
 BUF_X1 rebuffer94 (.A(_10338_),
    .Z(net724));
 BUF_X1 rebuffer95 (.A(_10359_),
    .Z(net725));
 BUF_X16 clone96 (.A(net727),
    .Z(net726));
 BUF_X1 rebuffer97 (.A(net729),
    .Z(net727));
 BUF_X16 clone98 (.A(net729),
    .Z(net728));
 BUF_X2 rebuffer99 (.A(_05309_),
    .Z(net729));
 BUF_X4 rebuffer104 (.A(_05264_),
    .Z(net734));
 BUF_X1 rebuffer105 (.A(_05141_),
    .Z(net735));
 BUF_X1 rebuffer106 (.A(_05142_),
    .Z(net736));
 BUF_X16 clone107 (.A(_05144_),
    .Z(net737));
 BUF_X16 clone108 (.A(_05143_),
    .Z(net738));
 BUF_X16 clone109 (.A(_05143_),
    .Z(net739));
 BUF_X16 clone110 (.A(net741),
    .Z(net740));
 BUF_X1 rebuffer111 (.A(_05142_),
    .Z(net741));
 AOI21_X2 clone114 (.A(_05610_),
    .B1(_05697_),
    .B2(_05696_),
    .ZN(net744));
 BUF_X1 rebuffer38 (.A(net691),
    .Z(net692));
 BUF_X1 rebuffer50 (.A(_05452_),
    .Z(net693));
 BUF_X1 rebuffer61 (.A(_07518_),
    .Z(net694));
 BUF_X1 rebuffer62 (.A(_10284_),
    .Z(net695));
 BUF_X1 rebuffer63 (.A(_00008_),
    .Z(net696));
 BUF_X1 rebuffer64 (.A(_10309_),
    .Z(net697));
 BUF_X1 rebuffer65 (.A(_10231_),
    .Z(net730));
 BUF_X1 rebuffer66 (.A(_10228_),
    .Z(net731));
 BUF_X1 rebuffer67 (.A(_10234_),
    .Z(net732));
 BUF_X1 rebuffer72 (.A(_00014_),
    .Z(net733));
 BUF_X1 rebuffer81 (.A(_07267_),
    .Z(net742));
 BUF_X16 clone82 (.A(_05130_),
    .Z(net743));
 BUF_X16 clone83 (.A(_05130_),
    .Z(net745));
 BUF_X16 clone84 (.A(net764),
    .Z(net746));
 BUF_X4 rebuffer87 (.A(_05695_),
    .Z(net747));
 BUF_X1 rebuffer90 (.A(net747),
    .Z(net748));
 BUF_X1 rebuffer91 (.A(net748),
    .Z(net749));
 BUF_X1 rebuffer96 (.A(_10231_),
    .Z(net750));
 BUF_X1 rebuffer98 (.A(net750),
    .Z(net751));
 BUF_X1 rebuffer101 (.A(net752),
    .Z(net753));
 BUF_X1 rebuffer102 (.A(net752),
    .Z(net754));
 BUF_X1 rebuffer108 (.A(net756),
    .Z(net757));
 BUF_X1 rebuffer121 (.A(_10246_),
    .Z(net771));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X16 FILLER_0_545 ();
 FILLCELL_X4 FILLER_0_564 ();
 FILLCELL_X2 FILLER_0_568 ();
 FILLCELL_X1 FILLER_0_573 ();
 FILLCELL_X2 FILLER_0_581 ();
 FILLCELL_X1 FILLER_0_583 ();
 FILLCELL_X1 FILLER_0_605 ();
 FILLCELL_X4 FILLER_0_609 ();
 FILLCELL_X1 FILLER_0_613 ();
 FILLCELL_X1 FILLER_0_639 ();
 FILLCELL_X2 FILLER_0_643 ();
 FILLCELL_X1 FILLER_0_656 ();
 FILLCELL_X2 FILLER_0_672 ();
 FILLCELL_X1 FILLER_0_674 ();
 FILLCELL_X1 FILLER_0_678 ();
 FILLCELL_X1 FILLER_0_682 ();
 FILLCELL_X1 FILLER_0_686 ();
 FILLCELL_X1 FILLER_0_708 ();
 FILLCELL_X2 FILLER_0_717 ();
 FILLCELL_X1 FILLER_0_770 ();
 FILLCELL_X2 FILLER_0_794 ();
 FILLCELL_X2 FILLER_0_809 ();
 FILLCELL_X4 FILLER_0_891 ();
 FILLCELL_X2 FILLER_0_904 ();
 FILLCELL_X1 FILLER_0_958 ();
 FILLCELL_X1 FILLER_0_978 ();
 FILLCELL_X2 FILLER_0_985 ();
 FILLCELL_X1 FILLER_0_987 ();
 FILLCELL_X1 FILLER_0_995 ();
 FILLCELL_X1 FILLER_0_999 ();
 FILLCELL_X1 FILLER_0_1043 ();
 FILLCELL_X1 FILLER_0_1047 ();
 FILLCELL_X1 FILLER_0_1054 ();
 FILLCELL_X1 FILLER_0_1061 ();
 FILLCELL_X1 FILLER_0_1069 ();
 FILLCELL_X1 FILLER_0_1131 ();
 FILLCELL_X32 FILLER_0_1154 ();
 FILLCELL_X32 FILLER_0_1186 ();
 FILLCELL_X16 FILLER_0_1218 ();
 FILLCELL_X4 FILLER_0_1234 ();
 FILLCELL_X2 FILLER_0_1238 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X4 FILLER_1_577 ();
 FILLCELL_X1 FILLER_1_581 ();
 FILLCELL_X16 FILLER_1_585 ();
 FILLCELL_X8 FILLER_1_601 ();
 FILLCELL_X2 FILLER_1_612 ();
 FILLCELL_X1 FILLER_1_614 ();
 FILLCELL_X8 FILLER_1_618 ();
 FILLCELL_X4 FILLER_1_626 ();
 FILLCELL_X1 FILLER_1_630 ();
 FILLCELL_X16 FILLER_1_639 ();
 FILLCELL_X4 FILLER_1_655 ();
 FILLCELL_X1 FILLER_1_659 ();
 FILLCELL_X8 FILLER_1_663 ();
 FILLCELL_X2 FILLER_1_680 ();
 FILLCELL_X1 FILLER_1_682 ();
 FILLCELL_X1 FILLER_1_686 ();
 FILLCELL_X1 FILLER_1_745 ();
 FILLCELL_X1 FILLER_1_757 ();
 FILLCELL_X1 FILLER_1_797 ();
 FILLCELL_X1 FILLER_1_840 ();
 FILLCELL_X1 FILLER_1_874 ();
 FILLCELL_X1 FILLER_1_899 ();
 FILLCELL_X2 FILLER_1_930 ();
 FILLCELL_X4 FILLER_1_939 ();
 FILLCELL_X1 FILLER_1_978 ();
 FILLCELL_X2 FILLER_1_1022 ();
 FILLCELL_X1 FILLER_1_1024 ();
 FILLCELL_X4 FILLER_1_1028 ();
 FILLCELL_X1 FILLER_1_1032 ();
 FILLCELL_X1 FILLER_1_1073 ();
 FILLCELL_X4 FILLER_1_1077 ();
 FILLCELL_X4 FILLER_1_1088 ();
 FILLCELL_X1 FILLER_1_1118 ();
 FILLCELL_X32 FILLER_1_1146 ();
 FILLCELL_X32 FILLER_1_1178 ();
 FILLCELL_X16 FILLER_1_1210 ();
 FILLCELL_X8 FILLER_1_1226 ();
 FILLCELL_X4 FILLER_1_1234 ();
 FILLCELL_X2 FILLER_1_1238 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X16 FILLER_2_577 ();
 FILLCELL_X8 FILLER_2_593 ();
 FILLCELL_X4 FILLER_2_601 ();
 FILLCELL_X1 FILLER_2_605 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X16 FILLER_2_632 ();
 FILLCELL_X8 FILLER_2_648 ();
 FILLCELL_X16 FILLER_2_659 ();
 FILLCELL_X8 FILLER_2_675 ();
 FILLCELL_X4 FILLER_2_683 ();
 FILLCELL_X1 FILLER_2_690 ();
 FILLCELL_X1 FILLER_2_712 ();
 FILLCELL_X1 FILLER_2_716 ();
 FILLCELL_X4 FILLER_2_782 ();
 FILLCELL_X4 FILLER_2_789 ();
 FILLCELL_X1 FILLER_2_793 ();
 FILLCELL_X2 FILLER_2_818 ();
 FILLCELL_X2 FILLER_2_830 ();
 FILLCELL_X1 FILLER_2_832 ();
 FILLCELL_X4 FILLER_2_836 ();
 FILLCELL_X8 FILLER_2_846 ();
 FILLCELL_X4 FILLER_2_884 ();
 FILLCELL_X2 FILLER_2_888 ();
 FILLCELL_X2 FILLER_2_898 ();
 FILLCELL_X8 FILLER_2_951 ();
 FILLCELL_X4 FILLER_2_959 ();
 FILLCELL_X1 FILLER_2_963 ();
 FILLCELL_X4 FILLER_2_967 ();
 FILLCELL_X2 FILLER_2_971 ();
 FILLCELL_X1 FILLER_2_973 ();
 FILLCELL_X1 FILLER_2_981 ();
 FILLCELL_X4 FILLER_2_989 ();
 FILLCELL_X8 FILLER_2_1000 ();
 FILLCELL_X4 FILLER_2_1032 ();
 FILLCELL_X4 FILLER_2_1123 ();
 FILLCELL_X32 FILLER_2_1130 ();
 FILLCELL_X32 FILLER_2_1162 ();
 FILLCELL_X32 FILLER_2_1194 ();
 FILLCELL_X8 FILLER_2_1226 ();
 FILLCELL_X4 FILLER_2_1234 ();
 FILLCELL_X2 FILLER_2_1238 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X4 FILLER_3_673 ();
 FILLCELL_X2 FILLER_3_677 ();
 FILLCELL_X1 FILLER_3_679 ();
 FILLCELL_X4 FILLER_3_704 ();
 FILLCELL_X2 FILLER_3_708 ();
 FILLCELL_X1 FILLER_3_736 ();
 FILLCELL_X1 FILLER_3_751 ();
 FILLCELL_X2 FILLER_3_766 ();
 FILLCELL_X1 FILLER_3_768 ();
 FILLCELL_X2 FILLER_3_786 ();
 FILLCELL_X1 FILLER_3_788 ();
 FILLCELL_X8 FILLER_3_815 ();
 FILLCELL_X2 FILLER_3_823 ();
 FILLCELL_X1 FILLER_3_825 ();
 FILLCELL_X8 FILLER_3_846 ();
 FILLCELL_X16 FILLER_3_857 ();
 FILLCELL_X1 FILLER_3_873 ();
 FILLCELL_X2 FILLER_3_881 ();
 FILLCELL_X8 FILLER_3_897 ();
 FILLCELL_X2 FILLER_3_905 ();
 FILLCELL_X1 FILLER_3_935 ();
 FILLCELL_X4 FILLER_3_960 ();
 FILLCELL_X1 FILLER_3_964 ();
 FILLCELL_X1 FILLER_3_991 ();
 FILLCELL_X8 FILLER_3_1016 ();
 FILLCELL_X2 FILLER_3_1072 ();
 FILLCELL_X4 FILLER_3_1081 ();
 FILLCELL_X2 FILLER_3_1092 ();
 FILLCELL_X1 FILLER_3_1104 ();
 FILLCELL_X32 FILLER_3_1119 ();
 FILLCELL_X32 FILLER_3_1151 ();
 FILLCELL_X32 FILLER_3_1183 ();
 FILLCELL_X16 FILLER_3_1215 ();
 FILLCELL_X8 FILLER_3_1231 ();
 FILLCELL_X1 FILLER_3_1239 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X16 FILLER_4_664 ();
 FILLCELL_X1 FILLER_4_680 ();
 FILLCELL_X4 FILLER_4_712 ();
 FILLCELL_X2 FILLER_4_716 ();
 FILLCELL_X4 FILLER_4_720 ();
 FILLCELL_X1 FILLER_4_724 ();
 FILLCELL_X16 FILLER_4_728 ();
 FILLCELL_X8 FILLER_4_744 ();
 FILLCELL_X2 FILLER_4_752 ();
 FILLCELL_X1 FILLER_4_771 ();
 FILLCELL_X16 FILLER_4_774 ();
 FILLCELL_X2 FILLER_4_790 ();
 FILLCELL_X2 FILLER_4_799 ();
 FILLCELL_X1 FILLER_4_818 ();
 FILLCELL_X4 FILLER_4_832 ();
 FILLCELL_X8 FILLER_4_853 ();
 FILLCELL_X2 FILLER_4_861 ();
 FILLCELL_X16 FILLER_4_865 ();
 FILLCELL_X4 FILLER_4_881 ();
 FILLCELL_X32 FILLER_4_909 ();
 FILLCELL_X4 FILLER_4_941 ();
 FILLCELL_X1 FILLER_4_945 ();
 FILLCELL_X2 FILLER_4_956 ();
 FILLCELL_X1 FILLER_4_958 ();
 FILLCELL_X1 FILLER_4_985 ();
 FILLCELL_X8 FILLER_4_989 ();
 FILLCELL_X4 FILLER_4_997 ();
 FILLCELL_X2 FILLER_4_1001 ();
 FILLCELL_X16 FILLER_4_1017 ();
 FILLCELL_X4 FILLER_4_1033 ();
 FILLCELL_X1 FILLER_4_1037 ();
 FILLCELL_X16 FILLER_4_1050 ();
 FILLCELL_X8 FILLER_4_1066 ();
 FILLCELL_X4 FILLER_4_1074 ();
 FILLCELL_X2 FILLER_4_1078 ();
 FILLCELL_X1 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1094 ();
 FILLCELL_X32 FILLER_4_1126 ();
 FILLCELL_X32 FILLER_4_1158 ();
 FILLCELL_X32 FILLER_4_1190 ();
 FILLCELL_X16 FILLER_4_1222 ();
 FILLCELL_X2 FILLER_4_1238 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X8 FILLER_5_737 ();
 FILLCELL_X4 FILLER_5_745 ();
 FILLCELL_X2 FILLER_5_749 ();
 FILLCELL_X8 FILLER_5_754 ();
 FILLCELL_X2 FILLER_5_762 ();
 FILLCELL_X1 FILLER_5_764 ();
 FILLCELL_X16 FILLER_5_791 ();
 FILLCELL_X8 FILLER_5_823 ();
 FILLCELL_X16 FILLER_5_854 ();
 FILLCELL_X8 FILLER_5_870 ();
 FILLCELL_X2 FILLER_5_883 ();
 FILLCELL_X1 FILLER_5_885 ();
 FILLCELL_X2 FILLER_5_903 ();
 FILLCELL_X1 FILLER_5_938 ();
 FILLCELL_X8 FILLER_5_964 ();
 FILLCELL_X1 FILLER_5_972 ();
 FILLCELL_X2 FILLER_5_986 ();
 FILLCELL_X1 FILLER_5_988 ();
 FILLCELL_X2 FILLER_5_1004 ();
 FILLCELL_X1 FILLER_5_1006 ();
 FILLCELL_X32 FILLER_5_1023 ();
 FILLCELL_X8 FILLER_5_1055 ();
 FILLCELL_X4 FILLER_5_1063 ();
 FILLCELL_X2 FILLER_5_1067 ();
 FILLCELL_X16 FILLER_5_1078 ();
 FILLCELL_X2 FILLER_5_1094 ();
 FILLCELL_X32 FILLER_5_1112 ();
 FILLCELL_X32 FILLER_5_1144 ();
 FILLCELL_X32 FILLER_5_1176 ();
 FILLCELL_X32 FILLER_5_1208 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X16 FILLER_6_664 ();
 FILLCELL_X8 FILLER_6_680 ();
 FILLCELL_X4 FILLER_6_688 ();
 FILLCELL_X4 FILLER_6_707 ();
 FILLCELL_X2 FILLER_6_711 ();
 FILLCELL_X1 FILLER_6_713 ();
 FILLCELL_X4 FILLER_6_719 ();
 FILLCELL_X8 FILLER_6_740 ();
 FILLCELL_X4 FILLER_6_748 ();
 FILLCELL_X1 FILLER_6_752 ();
 FILLCELL_X16 FILLER_6_770 ();
 FILLCELL_X8 FILLER_6_786 ();
 FILLCELL_X2 FILLER_6_794 ();
 FILLCELL_X1 FILLER_6_796 ();
 FILLCELL_X16 FILLER_6_804 ();
 FILLCELL_X8 FILLER_6_820 ();
 FILLCELL_X1 FILLER_6_828 ();
 FILLCELL_X2 FILLER_6_846 ();
 FILLCELL_X1 FILLER_6_848 ();
 FILLCELL_X4 FILLER_6_859 ();
 FILLCELL_X2 FILLER_6_863 ();
 FILLCELL_X4 FILLER_6_877 ();
 FILLCELL_X1 FILLER_6_881 ();
 FILLCELL_X2 FILLER_6_884 ();
 FILLCELL_X16 FILLER_6_924 ();
 FILLCELL_X1 FILLER_6_940 ();
 FILLCELL_X16 FILLER_6_965 ();
 FILLCELL_X8 FILLER_6_981 ();
 FILLCELL_X2 FILLER_6_989 ();
 FILLCELL_X1 FILLER_6_1015 ();
 FILLCELL_X32 FILLER_6_1042 ();
 FILLCELL_X8 FILLER_6_1074 ();
 FILLCELL_X4 FILLER_6_1082 ();
 FILLCELL_X1 FILLER_6_1086 ();
 FILLCELL_X4 FILLER_6_1101 ();
 FILLCELL_X2 FILLER_6_1105 ();
 FILLCELL_X32 FILLER_6_1124 ();
 FILLCELL_X32 FILLER_6_1156 ();
 FILLCELL_X32 FILLER_6_1188 ();
 FILLCELL_X16 FILLER_6_1220 ();
 FILLCELL_X4 FILLER_6_1236 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X8 FILLER_7_673 ();
 FILLCELL_X2 FILLER_7_681 ();
 FILLCELL_X1 FILLER_7_683 ();
 FILLCELL_X2 FILLER_7_718 ();
 FILLCELL_X1 FILLER_7_720 ();
 FILLCELL_X4 FILLER_7_738 ();
 FILLCELL_X2 FILLER_7_742 ();
 FILLCELL_X4 FILLER_7_761 ();
 FILLCELL_X16 FILLER_7_813 ();
 FILLCELL_X4 FILLER_7_829 ();
 FILLCELL_X1 FILLER_7_850 ();
 FILLCELL_X1 FILLER_7_864 ();
 FILLCELL_X1 FILLER_7_882 ();
 FILLCELL_X1 FILLER_7_890 ();
 FILLCELL_X16 FILLER_7_922 ();
 FILLCELL_X8 FILLER_7_938 ();
 FILLCELL_X16 FILLER_7_973 ();
 FILLCELL_X8 FILLER_7_989 ();
 FILLCELL_X2 FILLER_7_997 ();
 FILLCELL_X1 FILLER_7_999 ();
 FILLCELL_X4 FILLER_7_1017 ();
 FILLCELL_X8 FILLER_7_1042 ();
 FILLCELL_X2 FILLER_7_1050 ();
 FILLCELL_X1 FILLER_7_1052 ();
 FILLCELL_X8 FILLER_7_1070 ();
 FILLCELL_X4 FILLER_7_1078 ();
 FILLCELL_X1 FILLER_7_1082 ();
 FILLCELL_X32 FILLER_7_1124 ();
 FILLCELL_X32 FILLER_7_1156 ();
 FILLCELL_X32 FILLER_7_1188 ();
 FILLCELL_X16 FILLER_7_1220 ();
 FILLCELL_X4 FILLER_7_1236 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X16 FILLER_8_664 ();
 FILLCELL_X1 FILLER_8_680 ();
 FILLCELL_X4 FILLER_8_712 ();
 FILLCELL_X2 FILLER_8_716 ();
 FILLCELL_X1 FILLER_8_718 ();
 FILLCELL_X1 FILLER_8_726 ();
 FILLCELL_X4 FILLER_8_743 ();
 FILLCELL_X1 FILLER_8_766 ();
 FILLCELL_X2 FILLER_8_808 ();
 FILLCELL_X8 FILLER_8_817 ();
 FILLCELL_X4 FILLER_8_825 ();
 FILLCELL_X2 FILLER_8_829 ();
 FILLCELL_X2 FILLER_8_852 ();
 FILLCELL_X2 FILLER_8_878 ();
 FILLCELL_X4 FILLER_8_883 ();
 FILLCELL_X4 FILLER_8_922 ();
 FILLCELL_X2 FILLER_8_926 ();
 FILLCELL_X16 FILLER_8_952 ();
 FILLCELL_X8 FILLER_8_1009 ();
 FILLCELL_X4 FILLER_8_1017 ();
 FILLCELL_X2 FILLER_8_1038 ();
 FILLCELL_X4 FILLER_8_1078 ();
 FILLCELL_X1 FILLER_8_1082 ();
 FILLCELL_X2 FILLER_8_1107 ();
 FILLCELL_X32 FILLER_8_1116 ();
 FILLCELL_X32 FILLER_8_1148 ();
 FILLCELL_X32 FILLER_8_1180 ();
 FILLCELL_X16 FILLER_8_1212 ();
 FILLCELL_X8 FILLER_8_1228 ();
 FILLCELL_X4 FILLER_8_1236 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X4 FILLER_9_673 ();
 FILLCELL_X16 FILLER_9_715 ();
 FILLCELL_X4 FILLER_9_731 ();
 FILLCELL_X1 FILLER_9_735 ();
 FILLCELL_X1 FILLER_9_738 ();
 FILLCELL_X4 FILLER_9_747 ();
 FILLCELL_X8 FILLER_9_761 ();
 FILLCELL_X4 FILLER_9_769 ();
 FILLCELL_X1 FILLER_9_773 ();
 FILLCELL_X2 FILLER_9_784 ();
 FILLCELL_X16 FILLER_9_793 ();
 FILLCELL_X8 FILLER_9_809 ();
 FILLCELL_X16 FILLER_9_833 ();
 FILLCELL_X4 FILLER_9_849 ();
 FILLCELL_X4 FILLER_9_869 ();
 FILLCELL_X4 FILLER_9_886 ();
 FILLCELL_X1 FILLER_9_890 ();
 FILLCELL_X8 FILLER_9_917 ();
 FILLCELL_X4 FILLER_9_925 ();
 FILLCELL_X2 FILLER_9_929 ();
 FILLCELL_X1 FILLER_9_931 ();
 FILLCELL_X16 FILLER_9_949 ();
 FILLCELL_X8 FILLER_9_965 ();
 FILLCELL_X4 FILLER_9_973 ();
 FILLCELL_X1 FILLER_9_977 ();
 FILLCELL_X8 FILLER_9_992 ();
 FILLCELL_X4 FILLER_9_1000 ();
 FILLCELL_X2 FILLER_9_1004 ();
 FILLCELL_X8 FILLER_9_1031 ();
 FILLCELL_X2 FILLER_9_1039 ();
 FILLCELL_X1 FILLER_9_1041 ();
 FILLCELL_X8 FILLER_9_1059 ();
 FILLCELL_X8 FILLER_9_1083 ();
 FILLCELL_X4 FILLER_9_1091 ();
 FILLCELL_X32 FILLER_9_1104 ();
 FILLCELL_X32 FILLER_9_1136 ();
 FILLCELL_X32 FILLER_9_1168 ();
 FILLCELL_X32 FILLER_9_1200 ();
 FILLCELL_X8 FILLER_9_1232 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X4 FILLER_10_735 ();
 FILLCELL_X2 FILLER_10_756 ();
 FILLCELL_X8 FILLER_10_771 ();
 FILLCELL_X4 FILLER_10_779 ();
 FILLCELL_X2 FILLER_10_783 ();
 FILLCELL_X32 FILLER_10_815 ();
 FILLCELL_X16 FILLER_10_847 ();
 FILLCELL_X8 FILLER_10_863 ();
 FILLCELL_X1 FILLER_10_871 ();
 FILLCELL_X16 FILLER_10_879 ();
 FILLCELL_X4 FILLER_10_895 ();
 FILLCELL_X2 FILLER_10_899 ();
 FILLCELL_X1 FILLER_10_901 ();
 FILLCELL_X16 FILLER_10_918 ();
 FILLCELL_X4 FILLER_10_950 ();
 FILLCELL_X16 FILLER_10_957 ();
 FILLCELL_X8 FILLER_10_973 ();
 FILLCELL_X2 FILLER_10_981 ();
 FILLCELL_X16 FILLER_10_1024 ();
 FILLCELL_X2 FILLER_10_1040 ();
 FILLCELL_X32 FILLER_10_1074 ();
 FILLCELL_X32 FILLER_10_1106 ();
 FILLCELL_X32 FILLER_10_1138 ();
 FILLCELL_X32 FILLER_10_1170 ();
 FILLCELL_X32 FILLER_10_1202 ();
 FILLCELL_X4 FILLER_10_1234 ();
 FILLCELL_X2 FILLER_10_1238 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X16 FILLER_11_673 ();
 FILLCELL_X2 FILLER_11_694 ();
 FILLCELL_X2 FILLER_11_703 ();
 FILLCELL_X2 FILLER_11_712 ();
 FILLCELL_X2 FILLER_11_721 ();
 FILLCELL_X2 FILLER_11_754 ();
 FILLCELL_X1 FILLER_11_756 ();
 FILLCELL_X16 FILLER_11_781 ();
 FILLCELL_X4 FILLER_11_828 ();
 FILLCELL_X16 FILLER_11_866 ();
 FILLCELL_X8 FILLER_11_882 ();
 FILLCELL_X2 FILLER_11_890 ();
 FILLCELL_X1 FILLER_11_892 ();
 FILLCELL_X1 FILLER_11_900 ();
 FILLCELL_X8 FILLER_11_922 ();
 FILLCELL_X4 FILLER_11_930 ();
 FILLCELL_X2 FILLER_11_934 ();
 FILLCELL_X1 FILLER_11_936 ();
 FILLCELL_X4 FILLER_11_974 ();
 FILLCELL_X2 FILLER_11_978 ();
 FILLCELL_X1 FILLER_11_980 ();
 FILLCELL_X16 FILLER_11_1004 ();
 FILLCELL_X8 FILLER_11_1020 ();
 FILLCELL_X4 FILLER_11_1028 ();
 FILLCELL_X16 FILLER_11_1039 ();
 FILLCELL_X4 FILLER_11_1055 ();
 FILLCELL_X4 FILLER_11_1066 ();
 FILLCELL_X2 FILLER_11_1070 ();
 FILLCELL_X1 FILLER_11_1072 ();
 FILLCELL_X32 FILLER_11_1112 ();
 FILLCELL_X32 FILLER_11_1144 ();
 FILLCELL_X32 FILLER_11_1176 ();
 FILLCELL_X32 FILLER_11_1208 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X16 FILLER_12_664 ();
 FILLCELL_X8 FILLER_12_680 ();
 FILLCELL_X2 FILLER_12_688 ();
 FILLCELL_X1 FILLER_12_690 ();
 FILLCELL_X2 FILLER_12_725 ();
 FILLCELL_X1 FILLER_12_727 ();
 FILLCELL_X4 FILLER_12_730 ();
 FILLCELL_X1 FILLER_12_734 ();
 FILLCELL_X16 FILLER_12_742 ();
 FILLCELL_X4 FILLER_12_758 ();
 FILLCELL_X1 FILLER_12_762 ();
 FILLCELL_X4 FILLER_12_770 ();
 FILLCELL_X8 FILLER_12_786 ();
 FILLCELL_X1 FILLER_12_794 ();
 FILLCELL_X2 FILLER_12_802 ();
 FILLCELL_X1 FILLER_12_804 ();
 FILLCELL_X8 FILLER_12_830 ();
 FILLCELL_X1 FILLER_12_838 ();
 FILLCELL_X4 FILLER_12_846 ();
 FILLCELL_X1 FILLER_12_850 ();
 FILLCELL_X1 FILLER_12_867 ();
 FILLCELL_X4 FILLER_12_881 ();
 FILLCELL_X2 FILLER_12_885 ();
 FILLCELL_X1 FILLER_12_887 ();
 FILLCELL_X2 FILLER_12_936 ();
 FILLCELL_X2 FILLER_12_962 ();
 FILLCELL_X1 FILLER_12_964 ();
 FILLCELL_X4 FILLER_12_1022 ();
 FILLCELL_X1 FILLER_12_1026 ();
 FILLCELL_X1 FILLER_12_1051 ();
 FILLCELL_X2 FILLER_12_1069 ();
 FILLCELL_X1 FILLER_12_1071 ();
 FILLCELL_X1 FILLER_12_1110 ();
 FILLCELL_X32 FILLER_12_1128 ();
 FILLCELL_X32 FILLER_12_1160 ();
 FILLCELL_X32 FILLER_12_1192 ();
 FILLCELL_X16 FILLER_12_1224 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X16 FILLER_13_705 ();
 FILLCELL_X8 FILLER_13_721 ();
 FILLCELL_X2 FILLER_13_760 ();
 FILLCELL_X4 FILLER_13_782 ();
 FILLCELL_X2 FILLER_13_786 ();
 FILLCELL_X16 FILLER_13_822 ();
 FILLCELL_X2 FILLER_13_838 ();
 FILLCELL_X1 FILLER_13_840 ();
 FILLCELL_X2 FILLER_13_878 ();
 FILLCELL_X2 FILLER_13_904 ();
 FILLCELL_X8 FILLER_13_930 ();
 FILLCELL_X4 FILLER_13_952 ();
 FILLCELL_X2 FILLER_13_956 ();
 FILLCELL_X1 FILLER_13_982 ();
 FILLCELL_X1 FILLER_13_986 ();
 FILLCELL_X16 FILLER_13_1011 ();
 FILLCELL_X2 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1124 ();
 FILLCELL_X32 FILLER_13_1156 ();
 FILLCELL_X32 FILLER_13_1188 ();
 FILLCELL_X16 FILLER_13_1220 ();
 FILLCELL_X4 FILLER_13_1236 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X16 FILLER_14_664 ();
 FILLCELL_X4 FILLER_14_680 ();
 FILLCELL_X2 FILLER_14_684 ();
 FILLCELL_X16 FILLER_14_711 ();
 FILLCELL_X8 FILLER_14_727 ();
 FILLCELL_X2 FILLER_14_735 ();
 FILLCELL_X1 FILLER_14_737 ();
 FILLCELL_X16 FILLER_14_755 ();
 FILLCELL_X4 FILLER_14_773 ();
 FILLCELL_X2 FILLER_14_777 ();
 FILLCELL_X8 FILLER_14_809 ();
 FILLCELL_X8 FILLER_14_841 ();
 FILLCELL_X2 FILLER_14_849 ();
 FILLCELL_X1 FILLER_14_851 ();
 FILLCELL_X1 FILLER_14_866 ();
 FILLCELL_X2 FILLER_14_887 ();
 FILLCELL_X4 FILLER_14_896 ();
 FILLCELL_X1 FILLER_14_900 ();
 FILLCELL_X1 FILLER_14_910 ();
 FILLCELL_X2 FILLER_14_921 ();
 FILLCELL_X16 FILLER_14_936 ();
 FILLCELL_X8 FILLER_14_952 ();
 FILLCELL_X2 FILLER_14_960 ();
 FILLCELL_X1 FILLER_14_962 ();
 FILLCELL_X8 FILLER_14_983 ();
 FILLCELL_X4 FILLER_14_991 ();
 FILLCELL_X2 FILLER_14_995 ();
 FILLCELL_X32 FILLER_14_1014 ();
 FILLCELL_X4 FILLER_14_1046 ();
 FILLCELL_X2 FILLER_14_1050 ();
 FILLCELL_X1 FILLER_14_1052 ();
 FILLCELL_X32 FILLER_14_1062 ();
 FILLCELL_X32 FILLER_14_1094 ();
 FILLCELL_X32 FILLER_14_1126 ();
 FILLCELL_X32 FILLER_14_1158 ();
 FILLCELL_X32 FILLER_14_1190 ();
 FILLCELL_X16 FILLER_14_1222 ();
 FILLCELL_X2 FILLER_14_1238 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X1 FILLER_15_673 ();
 FILLCELL_X1 FILLER_15_705 ();
 FILLCELL_X16 FILLER_15_723 ();
 FILLCELL_X8 FILLER_15_739 ();
 FILLCELL_X4 FILLER_15_747 ();
 FILLCELL_X4 FILLER_15_761 ();
 FILLCELL_X2 FILLER_15_765 ();
 FILLCELL_X16 FILLER_15_772 ();
 FILLCELL_X8 FILLER_15_788 ();
 FILLCELL_X4 FILLER_15_796 ();
 FILLCELL_X4 FILLER_15_837 ();
 FILLCELL_X32 FILLER_15_860 ();
 FILLCELL_X8 FILLER_15_892 ();
 FILLCELL_X4 FILLER_15_900 ();
 FILLCELL_X2 FILLER_15_904 ();
 FILLCELL_X8 FILLER_15_911 ();
 FILLCELL_X1 FILLER_15_919 ();
 FILLCELL_X16 FILLER_15_927 ();
 FILLCELL_X4 FILLER_15_943 ();
 FILLCELL_X2 FILLER_15_947 ();
 FILLCELL_X16 FILLER_15_963 ();
 FILLCELL_X8 FILLER_15_979 ();
 FILLCELL_X4 FILLER_15_987 ();
 FILLCELL_X2 FILLER_15_991 ();
 FILLCELL_X1 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1016 ();
 FILLCELL_X16 FILLER_15_1048 ();
 FILLCELL_X8 FILLER_15_1064 ();
 FILLCELL_X4 FILLER_15_1072 ();
 FILLCELL_X2 FILLER_15_1076 ();
 FILLCELL_X1 FILLER_15_1078 ();
 FILLCELL_X8 FILLER_15_1086 ();
 FILLCELL_X1 FILLER_15_1094 ();
 FILLCELL_X32 FILLER_15_1119 ();
 FILLCELL_X32 FILLER_15_1151 ();
 FILLCELL_X32 FILLER_15_1183 ();
 FILLCELL_X16 FILLER_15_1215 ();
 FILLCELL_X8 FILLER_15_1231 ();
 FILLCELL_X1 FILLER_15_1239 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X16 FILLER_16_664 ();
 FILLCELL_X8 FILLER_16_687 ();
 FILLCELL_X1 FILLER_16_695 ();
 FILLCELL_X1 FILLER_16_698 ();
 FILLCELL_X1 FILLER_16_706 ();
 FILLCELL_X4 FILLER_16_714 ();
 FILLCELL_X1 FILLER_16_718 ();
 FILLCELL_X8 FILLER_16_729 ();
 FILLCELL_X4 FILLER_16_737 ();
 FILLCELL_X2 FILLER_16_741 ();
 FILLCELL_X4 FILLER_16_773 ();
 FILLCELL_X1 FILLER_16_777 ();
 FILLCELL_X1 FILLER_16_780 ();
 FILLCELL_X8 FILLER_16_801 ();
 FILLCELL_X2 FILLER_16_809 ();
 FILLCELL_X1 FILLER_16_811 ();
 FILLCELL_X4 FILLER_16_819 ();
 FILLCELL_X2 FILLER_16_823 ();
 FILLCELL_X8 FILLER_16_868 ();
 FILLCELL_X4 FILLER_16_876 ();
 FILLCELL_X16 FILLER_16_897 ();
 FILLCELL_X16 FILLER_16_930 ();
 FILLCELL_X4 FILLER_16_946 ();
 FILLCELL_X2 FILLER_16_950 ();
 FILLCELL_X16 FILLER_16_976 ();
 FILLCELL_X4 FILLER_16_1037 ();
 FILLCELL_X2 FILLER_16_1041 ();
 FILLCELL_X1 FILLER_16_1043 ();
 FILLCELL_X8 FILLER_16_1051 ();
 FILLCELL_X2 FILLER_16_1059 ();
 FILLCELL_X1 FILLER_16_1061 ();
 FILLCELL_X32 FILLER_16_1100 ();
 FILLCELL_X32 FILLER_16_1132 ();
 FILLCELL_X32 FILLER_16_1164 ();
 FILLCELL_X32 FILLER_16_1196 ();
 FILLCELL_X8 FILLER_16_1228 ();
 FILLCELL_X4 FILLER_16_1236 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X8 FILLER_17_735 ();
 FILLCELL_X2 FILLER_17_743 ();
 FILLCELL_X8 FILLER_17_752 ();
 FILLCELL_X2 FILLER_17_760 ();
 FILLCELL_X1 FILLER_17_776 ();
 FILLCELL_X16 FILLER_17_807 ();
 FILLCELL_X4 FILLER_17_823 ();
 FILLCELL_X2 FILLER_17_827 ();
 FILLCELL_X1 FILLER_17_829 ();
 FILLCELL_X4 FILLER_17_837 ();
 FILLCELL_X2 FILLER_17_856 ();
 FILLCELL_X2 FILLER_17_865 ();
 FILLCELL_X1 FILLER_17_874 ();
 FILLCELL_X4 FILLER_17_889 ();
 FILLCELL_X1 FILLER_17_893 ();
 FILLCELL_X8 FILLER_17_918 ();
 FILLCELL_X2 FILLER_17_933 ();
 FILLCELL_X8 FILLER_17_942 ();
 FILLCELL_X2 FILLER_17_967 ();
 FILLCELL_X2 FILLER_17_993 ();
 FILLCELL_X1 FILLER_17_995 ();
 FILLCELL_X2 FILLER_17_1016 ();
 FILLCELL_X1 FILLER_17_1018 ();
 FILLCELL_X2 FILLER_17_1033 ();
 FILLCELL_X1 FILLER_17_1035 ();
 FILLCELL_X1 FILLER_17_1043 ();
 FILLCELL_X1 FILLER_17_1061 ();
 FILLCELL_X1 FILLER_17_1069 ();
 FILLCELL_X1 FILLER_17_1087 ();
 FILLCELL_X1 FILLER_17_1112 ();
 FILLCELL_X4 FILLER_17_1130 ();
 FILLCELL_X2 FILLER_17_1134 ();
 FILLCELL_X1 FILLER_17_1136 ();
 FILLCELL_X32 FILLER_17_1154 ();
 FILLCELL_X32 FILLER_17_1186 ();
 FILLCELL_X16 FILLER_17_1218 ();
 FILLCELL_X4 FILLER_17_1234 ();
 FILLCELL_X2 FILLER_17_1238 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X4 FILLER_18_664 ();
 FILLCELL_X1 FILLER_18_668 ();
 FILLCELL_X4 FILLER_18_686 ();
 FILLCELL_X8 FILLER_18_697 ();
 FILLCELL_X4 FILLER_18_705 ();
 FILLCELL_X2 FILLER_18_711 ();
 FILLCELL_X4 FILLER_18_720 ();
 FILLCELL_X2 FILLER_18_724 ();
 FILLCELL_X1 FILLER_18_726 ();
 FILLCELL_X4 FILLER_18_775 ();
 FILLCELL_X16 FILLER_18_800 ();
 FILLCELL_X2 FILLER_18_816 ();
 FILLCELL_X16 FILLER_18_823 ();
 FILLCELL_X2 FILLER_18_839 ();
 FILLCELL_X1 FILLER_18_992 ();
 FILLCELL_X2 FILLER_18_1041 ();
 FILLCELL_X1 FILLER_18_1043 ();
 FILLCELL_X16 FILLER_18_1061 ();
 FILLCELL_X8 FILLER_18_1077 ();
 FILLCELL_X2 FILLER_18_1085 ();
 FILLCELL_X16 FILLER_18_1096 ();
 FILLCELL_X2 FILLER_18_1112 ();
 FILLCELL_X16 FILLER_18_1121 ();
 FILLCELL_X2 FILLER_18_1137 ();
 FILLCELL_X16 FILLER_18_1156 ();
 FILLCELL_X4 FILLER_18_1172 ();
 FILLCELL_X1 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1194 ();
 FILLCELL_X8 FILLER_18_1226 ();
 FILLCELL_X4 FILLER_18_1234 ();
 FILLCELL_X2 FILLER_18_1238 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X16 FILLER_19_641 ();
 FILLCELL_X8 FILLER_19_657 ();
 FILLCELL_X4 FILLER_19_665 ();
 FILLCELL_X1 FILLER_19_669 ();
 FILLCELL_X2 FILLER_19_694 ();
 FILLCELL_X1 FILLER_19_696 ();
 FILLCELL_X2 FILLER_19_761 ();
 FILLCELL_X1 FILLER_19_763 ();
 FILLCELL_X8 FILLER_19_766 ();
 FILLCELL_X2 FILLER_19_774 ();
 FILLCELL_X1 FILLER_19_776 ();
 FILLCELL_X4 FILLER_19_801 ();
 FILLCELL_X4 FILLER_19_829 ();
 FILLCELL_X16 FILLER_19_840 ();
 FILLCELL_X8 FILLER_19_856 ();
 FILLCELL_X4 FILLER_19_864 ();
 FILLCELL_X2 FILLER_19_868 ();
 FILLCELL_X1 FILLER_19_870 ();
 FILLCELL_X4 FILLER_19_878 ();
 FILLCELL_X2 FILLER_19_882 ();
 FILLCELL_X1 FILLER_19_884 ();
 FILLCELL_X1 FILLER_19_910 ();
 FILLCELL_X1 FILLER_19_918 ();
 FILLCELL_X1 FILLER_19_970 ();
 FILLCELL_X4 FILLER_19_1013 ();
 FILLCELL_X16 FILLER_19_1035 ();
 FILLCELL_X8 FILLER_19_1051 ();
 FILLCELL_X4 FILLER_19_1100 ();
 FILLCELL_X1 FILLER_19_1142 ();
 FILLCELL_X8 FILLER_19_1157 ();
 FILLCELL_X1 FILLER_19_1173 ();
 FILLCELL_X2 FILLER_19_1181 ();
 FILLCELL_X1 FILLER_19_1183 ();
 FILLCELL_X32 FILLER_19_1191 ();
 FILLCELL_X16 FILLER_19_1223 ();
 FILLCELL_X1 FILLER_19_1239 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X16 FILLER_20_632 ();
 FILLCELL_X4 FILLER_20_648 ();
 FILLCELL_X4 FILLER_20_676 ();
 FILLCELL_X1 FILLER_20_680 ();
 FILLCELL_X1 FILLER_20_688 ();
 FILLCELL_X1 FILLER_20_696 ();
 FILLCELL_X1 FILLER_20_704 ();
 FILLCELL_X2 FILLER_20_722 ();
 FILLCELL_X1 FILLER_20_724 ();
 FILLCELL_X8 FILLER_20_733 ();
 FILLCELL_X2 FILLER_20_741 ();
 FILLCELL_X8 FILLER_20_750 ();
 FILLCELL_X4 FILLER_20_758 ();
 FILLCELL_X1 FILLER_20_762 ();
 FILLCELL_X2 FILLER_20_770 ();
 FILLCELL_X4 FILLER_20_775 ();
 FILLCELL_X1 FILLER_20_779 ();
 FILLCELL_X8 FILLER_20_787 ();
 FILLCELL_X4 FILLER_20_795 ();
 FILLCELL_X1 FILLER_20_799 ();
 FILLCELL_X32 FILLER_20_843 ();
 FILLCELL_X2 FILLER_20_875 ();
 FILLCELL_X1 FILLER_20_877 ();
 FILLCELL_X16 FILLER_20_880 ();
 FILLCELL_X2 FILLER_20_896 ();
 FILLCELL_X8 FILLER_20_905 ();
 FILLCELL_X4 FILLER_20_913 ();
 FILLCELL_X1 FILLER_20_917 ();
 FILLCELL_X4 FILLER_20_925 ();
 FILLCELL_X2 FILLER_20_929 ();
 FILLCELL_X1 FILLER_20_931 ();
 FILLCELL_X1 FILLER_20_993 ();
 FILLCELL_X16 FILLER_20_1043 ();
 FILLCELL_X4 FILLER_20_1059 ();
 FILLCELL_X2 FILLER_20_1063 ();
 FILLCELL_X32 FILLER_20_1079 ();
 FILLCELL_X32 FILLER_20_1121 ();
 FILLCELL_X16 FILLER_20_1153 ();
 FILLCELL_X8 FILLER_20_1169 ();
 FILLCELL_X1 FILLER_20_1177 ();
 FILLCELL_X32 FILLER_20_1202 ();
 FILLCELL_X4 FILLER_20_1234 ();
 FILLCELL_X2 FILLER_20_1238 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X4 FILLER_21_641 ();
 FILLCELL_X8 FILLER_21_686 ();
 FILLCELL_X4 FILLER_21_694 ();
 FILLCELL_X16 FILLER_21_712 ();
 FILLCELL_X8 FILLER_21_742 ();
 FILLCELL_X1 FILLER_21_750 ();
 FILLCELL_X4 FILLER_21_758 ();
 FILLCELL_X1 FILLER_21_762 ();
 FILLCELL_X8 FILLER_21_793 ();
 FILLCELL_X4 FILLER_21_801 ();
 FILLCELL_X4 FILLER_21_836 ();
 FILLCELL_X2 FILLER_21_857 ();
 FILLCELL_X4 FILLER_21_864 ();
 FILLCELL_X1 FILLER_21_868 ();
 FILLCELL_X8 FILLER_21_898 ();
 FILLCELL_X1 FILLER_21_906 ();
 FILLCELL_X32 FILLER_21_914 ();
 FILLCELL_X2 FILLER_21_946 ();
 FILLCELL_X1 FILLER_21_948 ();
 FILLCELL_X2 FILLER_21_956 ();
 FILLCELL_X1 FILLER_21_958 ();
 FILLCELL_X4 FILLER_21_962 ();
 FILLCELL_X2 FILLER_21_966 ();
 FILLCELL_X4 FILLER_21_977 ();
 FILLCELL_X1 FILLER_21_981 ();
 FILLCELL_X1 FILLER_21_994 ();
 FILLCELL_X4 FILLER_21_1012 ();
 FILLCELL_X1 FILLER_21_1016 ();
 FILLCELL_X8 FILLER_21_1033 ();
 FILLCELL_X4 FILLER_21_1041 ();
 FILLCELL_X2 FILLER_21_1045 ();
 FILLCELL_X16 FILLER_21_1052 ();
 FILLCELL_X8 FILLER_21_1068 ();
 FILLCELL_X4 FILLER_21_1076 ();
 FILLCELL_X2 FILLER_21_1080 ();
 FILLCELL_X4 FILLER_21_1099 ();
 FILLCELL_X2 FILLER_21_1103 ();
 FILLCELL_X2 FILLER_21_1129 ();
 FILLCELL_X8 FILLER_21_1135 ();
 FILLCELL_X2 FILLER_21_1143 ();
 FILLCELL_X1 FILLER_21_1145 ();
 FILLCELL_X8 FILLER_21_1150 ();
 FILLCELL_X32 FILLER_21_1186 ();
 FILLCELL_X2 FILLER_21_1218 ();
 FILLCELL_X2 FILLER_21_1237 ();
 FILLCELL_X1 FILLER_21_1239 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X16 FILLER_22_385 ();
 FILLCELL_X8 FILLER_22_401 ();
 FILLCELL_X2 FILLER_22_409 ();
 FILLCELL_X32 FILLER_22_415 ();
 FILLCELL_X32 FILLER_22_447 ();
 FILLCELL_X32 FILLER_22_479 ();
 FILLCELL_X32 FILLER_22_511 ();
 FILLCELL_X32 FILLER_22_543 ();
 FILLCELL_X32 FILLER_22_575 ();
 FILLCELL_X16 FILLER_22_607 ();
 FILLCELL_X8 FILLER_22_623 ();
 FILLCELL_X8 FILLER_22_632 ();
 FILLCELL_X1 FILLER_22_640 ();
 FILLCELL_X16 FILLER_22_686 ();
 FILLCELL_X8 FILLER_22_702 ();
 FILLCELL_X4 FILLER_22_710 ();
 FILLCELL_X1 FILLER_22_714 ();
 FILLCELL_X16 FILLER_22_756 ();
 FILLCELL_X8 FILLER_22_772 ();
 FILLCELL_X2 FILLER_22_780 ();
 FILLCELL_X1 FILLER_22_782 ();
 FILLCELL_X16 FILLER_22_790 ();
 FILLCELL_X1 FILLER_22_806 ();
 FILLCELL_X1 FILLER_22_814 ();
 FILLCELL_X2 FILLER_22_822 ();
 FILLCELL_X1 FILLER_22_824 ();
 FILLCELL_X16 FILLER_22_872 ();
 FILLCELL_X2 FILLER_22_888 ();
 FILLCELL_X8 FILLER_22_907 ();
 FILLCELL_X4 FILLER_22_915 ();
 FILLCELL_X1 FILLER_22_919 ();
 FILLCELL_X8 FILLER_22_944 ();
 FILLCELL_X1 FILLER_22_952 ();
 FILLCELL_X4 FILLER_22_987 ();
 FILLCELL_X1 FILLER_22_991 ();
 FILLCELL_X1 FILLER_22_1009 ();
 FILLCELL_X4 FILLER_22_1017 ();
 FILLCELL_X2 FILLER_22_1021 ();
 FILLCELL_X2 FILLER_22_1040 ();
 FILLCELL_X1 FILLER_22_1042 ();
 FILLCELL_X8 FILLER_22_1060 ();
 FILLCELL_X4 FILLER_22_1068 ();
 FILLCELL_X2 FILLER_22_1079 ();
 FILLCELL_X4 FILLER_22_1124 ();
 FILLCELL_X4 FILLER_22_1162 ();
 FILLCELL_X4 FILLER_22_1194 ();
 FILLCELL_X2 FILLER_22_1215 ();
 FILLCELL_X16 FILLER_22_1224 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X8 FILLER_23_673 ();
 FILLCELL_X4 FILLER_23_681 ();
 FILLCELL_X2 FILLER_23_685 ();
 FILLCELL_X8 FILLER_23_696 ();
 FILLCELL_X4 FILLER_23_704 ();
 FILLCELL_X2 FILLER_23_708 ();
 FILLCELL_X8 FILLER_23_727 ();
 FILLCELL_X4 FILLER_23_735 ();
 FILLCELL_X4 FILLER_23_746 ();
 FILLCELL_X2 FILLER_23_764 ();
 FILLCELL_X1 FILLER_23_766 ();
 FILLCELL_X1 FILLER_23_798 ();
 FILLCELL_X4 FILLER_23_823 ();
 FILLCELL_X1 FILLER_23_827 ();
 FILLCELL_X8 FILLER_23_855 ();
 FILLCELL_X1 FILLER_23_870 ();
 FILLCELL_X2 FILLER_23_878 ();
 FILLCELL_X2 FILLER_23_887 ();
 FILLCELL_X1 FILLER_23_889 ();
 FILLCELL_X1 FILLER_23_931 ();
 FILLCELL_X4 FILLER_23_954 ();
 FILLCELL_X2 FILLER_23_958 ();
 FILLCELL_X1 FILLER_23_960 ();
 FILLCELL_X8 FILLER_23_975 ();
 FILLCELL_X2 FILLER_23_983 ();
 FILLCELL_X4 FILLER_23_1034 ();
 FILLCELL_X2 FILLER_23_1038 ();
 FILLCELL_X4 FILLER_23_1064 ();
 FILLCELL_X4 FILLER_23_1085 ();
 FILLCELL_X4 FILLER_23_1096 ();
 FILLCELL_X8 FILLER_23_1124 ();
 FILLCELL_X2 FILLER_23_1132 ();
 FILLCELL_X1 FILLER_23_1134 ();
 FILLCELL_X4 FILLER_23_1149 ();
 FILLCELL_X2 FILLER_23_1153 ();
 FILLCELL_X8 FILLER_23_1162 ();
 FILLCELL_X1 FILLER_23_1177 ();
 FILLCELL_X1 FILLER_23_1191 ();
 FILLCELL_X1 FILLER_23_1199 ();
 FILLCELL_X2 FILLER_23_1217 ();
 FILLCELL_X4 FILLER_23_1236 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X4 FILLER_24_17 ();
 FILLCELL_X1 FILLER_24_21 ();
 FILLCELL_X32 FILLER_24_26 ();
 FILLCELL_X32 FILLER_24_58 ();
 FILLCELL_X32 FILLER_24_90 ();
 FILLCELL_X32 FILLER_24_122 ();
 FILLCELL_X32 FILLER_24_154 ();
 FILLCELL_X32 FILLER_24_186 ();
 FILLCELL_X32 FILLER_24_218 ();
 FILLCELL_X32 FILLER_24_250 ();
 FILLCELL_X32 FILLER_24_282 ();
 FILLCELL_X32 FILLER_24_314 ();
 FILLCELL_X32 FILLER_24_346 ();
 FILLCELL_X32 FILLER_24_378 ();
 FILLCELL_X32 FILLER_24_410 ();
 FILLCELL_X32 FILLER_24_442 ();
 FILLCELL_X32 FILLER_24_474 ();
 FILLCELL_X32 FILLER_24_506 ();
 FILLCELL_X32 FILLER_24_538 ();
 FILLCELL_X32 FILLER_24_570 ();
 FILLCELL_X16 FILLER_24_602 ();
 FILLCELL_X8 FILLER_24_618 ();
 FILLCELL_X4 FILLER_24_626 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X8 FILLER_24_664 ();
 FILLCELL_X2 FILLER_24_672 ();
 FILLCELL_X16 FILLER_24_698 ();
 FILLCELL_X2 FILLER_24_714 ();
 FILLCELL_X1 FILLER_24_716 ();
 FILLCELL_X1 FILLER_24_731 ();
 FILLCELL_X16 FILLER_24_773 ();
 FILLCELL_X4 FILLER_24_789 ();
 FILLCELL_X1 FILLER_24_855 ();
 FILLCELL_X4 FILLER_24_861 ();
 FILLCELL_X2 FILLER_24_865 ();
 FILLCELL_X4 FILLER_24_887 ();
 FILLCELL_X1 FILLER_24_898 ();
 FILLCELL_X4 FILLER_24_906 ();
 FILLCELL_X1 FILLER_24_910 ();
 FILLCELL_X1 FILLER_24_918 ();
 FILLCELL_X2 FILLER_24_962 ();
 FILLCELL_X8 FILLER_24_976 ();
 FILLCELL_X4 FILLER_24_984 ();
 FILLCELL_X16 FILLER_24_1009 ();
 FILLCELL_X2 FILLER_24_1025 ();
 FILLCELL_X2 FILLER_24_1034 ();
 FILLCELL_X1 FILLER_24_1036 ();
 FILLCELL_X4 FILLER_24_1051 ();
 FILLCELL_X2 FILLER_24_1055 ();
 FILLCELL_X8 FILLER_24_1064 ();
 FILLCELL_X4 FILLER_24_1072 ();
 FILLCELL_X2 FILLER_24_1076 ();
 FILLCELL_X8 FILLER_24_1109 ();
 FILLCELL_X8 FILLER_24_1130 ();
 FILLCELL_X2 FILLER_24_1138 ();
 FILLCELL_X4 FILLER_24_1153 ();
 FILLCELL_X16 FILLER_24_1162 ();
 FILLCELL_X8 FILLER_24_1178 ();
 FILLCELL_X4 FILLER_24_1213 ();
 FILLCELL_X1 FILLER_24_1217 ();
 FILLCELL_X8 FILLER_24_1232 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_9 ();
 FILLCELL_X1 FILLER_25_11 ();
 FILLCELL_X32 FILLER_25_16 ();
 FILLCELL_X32 FILLER_25_48 ();
 FILLCELL_X32 FILLER_25_80 ();
 FILLCELL_X32 FILLER_25_112 ();
 FILLCELL_X32 FILLER_25_144 ();
 FILLCELL_X32 FILLER_25_176 ();
 FILLCELL_X32 FILLER_25_208 ();
 FILLCELL_X32 FILLER_25_240 ();
 FILLCELL_X32 FILLER_25_272 ();
 FILLCELL_X32 FILLER_25_304 ();
 FILLCELL_X32 FILLER_25_336 ();
 FILLCELL_X32 FILLER_25_368 ();
 FILLCELL_X32 FILLER_25_400 ();
 FILLCELL_X32 FILLER_25_432 ();
 FILLCELL_X32 FILLER_25_464 ();
 FILLCELL_X32 FILLER_25_496 ();
 FILLCELL_X32 FILLER_25_528 ();
 FILLCELL_X32 FILLER_25_560 ();
 FILLCELL_X32 FILLER_25_592 ();
 FILLCELL_X16 FILLER_25_624 ();
 FILLCELL_X8 FILLER_25_640 ();
 FILLCELL_X2 FILLER_25_648 ();
 FILLCELL_X8 FILLER_25_686 ();
 FILLCELL_X2 FILLER_25_694 ();
 FILLCELL_X4 FILLER_25_703 ();
 FILLCELL_X16 FILLER_25_715 ();
 FILLCELL_X2 FILLER_25_731 ();
 FILLCELL_X1 FILLER_25_733 ();
 FILLCELL_X16 FILLER_25_737 ();
 FILLCELL_X8 FILLER_25_753 ();
 FILLCELL_X2 FILLER_25_761 ();
 FILLCELL_X1 FILLER_25_763 ();
 FILLCELL_X8 FILLER_25_771 ();
 FILLCELL_X1 FILLER_25_779 ();
 FILLCELL_X4 FILLER_25_815 ();
 FILLCELL_X1 FILLER_25_819 ();
 FILLCELL_X1 FILLER_25_837 ();
 FILLCELL_X16 FILLER_25_869 ();
 FILLCELL_X4 FILLER_25_885 ();
 FILLCELL_X2 FILLER_25_889 ();
 FILLCELL_X16 FILLER_25_908 ();
 FILLCELL_X2 FILLER_25_924 ();
 FILLCELL_X1 FILLER_25_926 ();
 FILLCELL_X2 FILLER_25_929 ();
 FILLCELL_X4 FILLER_25_938 ();
 FILLCELL_X1 FILLER_25_942 ();
 FILLCELL_X4 FILLER_25_957 ();
 FILLCELL_X2 FILLER_25_961 ();
 FILLCELL_X1 FILLER_25_963 ();
 FILLCELL_X32 FILLER_25_971 ();
 FILLCELL_X16 FILLER_25_1003 ();
 FILLCELL_X4 FILLER_25_1019 ();
 FILLCELL_X1 FILLER_25_1023 ();
 FILLCELL_X16 FILLER_25_1048 ();
 FILLCELL_X8 FILLER_25_1064 ();
 FILLCELL_X4 FILLER_25_1072 ();
 FILLCELL_X2 FILLER_25_1076 ();
 FILLCELL_X1 FILLER_25_1078 ();
 FILLCELL_X32 FILLER_25_1084 ();
 FILLCELL_X32 FILLER_25_1116 ();
 FILLCELL_X1 FILLER_25_1148 ();
 FILLCELL_X8 FILLER_25_1170 ();
 FILLCELL_X4 FILLER_25_1178 ();
 FILLCELL_X2 FILLER_25_1182 ();
 FILLCELL_X4 FILLER_25_1204 ();
 FILLCELL_X1 FILLER_25_1208 ();
 FILLCELL_X4 FILLER_25_1212 ();
 FILLCELL_X16 FILLER_25_1224 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X8 FILLER_26_97 ();
 FILLCELL_X4 FILLER_26_105 ();
 FILLCELL_X2 FILLER_26_109 ();
 FILLCELL_X1 FILLER_26_111 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X4 FILLER_26_664 ();
 FILLCELL_X1 FILLER_26_699 ();
 FILLCELL_X8 FILLER_26_720 ();
 FILLCELL_X2 FILLER_26_728 ();
 FILLCELL_X16 FILLER_26_777 ();
 FILLCELL_X8 FILLER_26_793 ();
 FILLCELL_X2 FILLER_26_801 ();
 FILLCELL_X1 FILLER_26_803 ();
 FILLCELL_X1 FILLER_26_821 ();
 FILLCELL_X2 FILLER_26_829 ();
 FILLCELL_X1 FILLER_26_831 ();
 FILLCELL_X8 FILLER_26_869 ();
 FILLCELL_X2 FILLER_26_877 ();
 FILLCELL_X1 FILLER_26_879 ();
 FILLCELL_X8 FILLER_26_889 ();
 FILLCELL_X4 FILLER_26_897 ();
 FILLCELL_X2 FILLER_26_901 ();
 FILLCELL_X1 FILLER_26_903 ();
 FILLCELL_X8 FILLER_26_909 ();
 FILLCELL_X1 FILLER_26_917 ();
 FILLCELL_X4 FILLER_26_921 ();
 FILLCELL_X16 FILLER_26_932 ();
 FILLCELL_X1 FILLER_26_948 ();
 FILLCELL_X2 FILLER_26_962 ();
 FILLCELL_X2 FILLER_26_998 ();
 FILLCELL_X32 FILLER_26_1008 ();
 FILLCELL_X16 FILLER_26_1040 ();
 FILLCELL_X1 FILLER_26_1056 ();
 FILLCELL_X4 FILLER_26_1061 ();
 FILLCELL_X2 FILLER_26_1065 ();
 FILLCELL_X1 FILLER_26_1067 ();
 FILLCELL_X8 FILLER_26_1073 ();
 FILLCELL_X4 FILLER_26_1081 ();
 FILLCELL_X2 FILLER_26_1085 ();
 FILLCELL_X16 FILLER_26_1104 ();
 FILLCELL_X8 FILLER_26_1120 ();
 FILLCELL_X8 FILLER_26_1179 ();
 FILLCELL_X4 FILLER_26_1204 ();
 FILLCELL_X2 FILLER_26_1208 ();
 FILLCELL_X4 FILLER_26_1234 ();
 FILLCELL_X2 FILLER_26_1238 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_97 ();
 FILLCELL_X8 FILLER_27_113 ();
 FILLCELL_X4 FILLER_27_121 ();
 FILLCELL_X1 FILLER_27_125 ();
 FILLCELL_X32 FILLER_27_157 ();
 FILLCELL_X32 FILLER_27_189 ();
 FILLCELL_X32 FILLER_27_221 ();
 FILLCELL_X32 FILLER_27_253 ();
 FILLCELL_X32 FILLER_27_285 ();
 FILLCELL_X32 FILLER_27_317 ();
 FILLCELL_X32 FILLER_27_349 ();
 FILLCELL_X32 FILLER_27_381 ();
 FILLCELL_X32 FILLER_27_413 ();
 FILLCELL_X32 FILLER_27_445 ();
 FILLCELL_X32 FILLER_27_477 ();
 FILLCELL_X32 FILLER_27_509 ();
 FILLCELL_X32 FILLER_27_541 ();
 FILLCELL_X32 FILLER_27_573 ();
 FILLCELL_X32 FILLER_27_605 ();
 FILLCELL_X16 FILLER_27_637 ();
 FILLCELL_X4 FILLER_27_653 ();
 FILLCELL_X2 FILLER_27_657 ();
 FILLCELL_X8 FILLER_27_676 ();
 FILLCELL_X1 FILLER_27_701 ();
 FILLCELL_X1 FILLER_27_704 ();
 FILLCELL_X1 FILLER_27_722 ();
 FILLCELL_X2 FILLER_27_730 ();
 FILLCELL_X8 FILLER_27_739 ();
 FILLCELL_X4 FILLER_27_747 ();
 FILLCELL_X1 FILLER_27_751 ();
 FILLCELL_X4 FILLER_27_759 ();
 FILLCELL_X1 FILLER_27_763 ();
 FILLCELL_X4 FILLER_27_767 ();
 FILLCELL_X2 FILLER_27_771 ();
 FILLCELL_X16 FILLER_27_780 ();
 FILLCELL_X4 FILLER_27_796 ();
 FILLCELL_X1 FILLER_27_800 ();
 FILLCELL_X16 FILLER_27_811 ();
 FILLCELL_X1 FILLER_27_827 ();
 FILLCELL_X4 FILLER_27_883 ();
 FILLCELL_X2 FILLER_27_887 ();
 FILLCELL_X1 FILLER_27_896 ();
 FILLCELL_X4 FILLER_27_914 ();
 FILLCELL_X2 FILLER_27_918 ();
 FILLCELL_X4 FILLER_27_937 ();
 FILLCELL_X1 FILLER_27_941 ();
 FILLCELL_X4 FILLER_27_959 ();
 FILLCELL_X1 FILLER_27_963 ();
 FILLCELL_X4 FILLER_27_981 ();
 FILLCELL_X8 FILLER_27_992 ();
 FILLCELL_X1 FILLER_27_1000 ();
 FILLCELL_X8 FILLER_27_1008 ();
 FILLCELL_X2 FILLER_27_1016 ();
 FILLCELL_X1 FILLER_27_1018 ();
 FILLCELL_X4 FILLER_27_1067 ();
 FILLCELL_X8 FILLER_27_1100 ();
 FILLCELL_X2 FILLER_27_1108 ();
 FILLCELL_X8 FILLER_27_1169 ();
 FILLCELL_X2 FILLER_27_1177 ();
 FILLCELL_X1 FILLER_27_1179 ();
 FILLCELL_X4 FILLER_27_1198 ();
 FILLCELL_X16 FILLER_27_1216 ();
 FILLCELL_X8 FILLER_27_1232 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X16 FILLER_28_65 ();
 FILLCELL_X4 FILLER_28_81 ();
 FILLCELL_X1 FILLER_28_85 ();
 FILLCELL_X8 FILLER_28_103 ();
 FILLCELL_X1 FILLER_28_111 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X1 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_179 ();
 FILLCELL_X8 FILLER_28_211 ();
 FILLCELL_X1 FILLER_28_219 ();
 FILLCELL_X4 FILLER_28_237 ();
 FILLCELL_X2 FILLER_28_241 ();
 FILLCELL_X1 FILLER_28_243 ();
 FILLCELL_X32 FILLER_28_261 ();
 FILLCELL_X32 FILLER_28_293 ();
 FILLCELL_X32 FILLER_28_325 ();
 FILLCELL_X1 FILLER_28_357 ();
 FILLCELL_X32 FILLER_28_361 ();
 FILLCELL_X32 FILLER_28_393 ();
 FILLCELL_X32 FILLER_28_425 ();
 FILLCELL_X32 FILLER_28_457 ();
 FILLCELL_X32 FILLER_28_489 ();
 FILLCELL_X32 FILLER_28_521 ();
 FILLCELL_X32 FILLER_28_553 ();
 FILLCELL_X32 FILLER_28_585 ();
 FILLCELL_X8 FILLER_28_617 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X8 FILLER_28_664 ();
 FILLCELL_X16 FILLER_28_703 ();
 FILLCELL_X4 FILLER_28_719 ();
 FILLCELL_X2 FILLER_28_723 ();
 FILLCELL_X1 FILLER_28_725 ();
 FILLCELL_X4 FILLER_28_733 ();
 FILLCELL_X1 FILLER_28_737 ();
 FILLCELL_X2 FILLER_28_740 ();
 FILLCELL_X1 FILLER_28_742 ();
 FILLCELL_X2 FILLER_28_759 ();
 FILLCELL_X1 FILLER_28_761 ();
 FILLCELL_X8 FILLER_28_786 ();
 FILLCELL_X16 FILLER_28_828 ();
 FILLCELL_X8 FILLER_28_844 ();
 FILLCELL_X4 FILLER_28_852 ();
 FILLCELL_X2 FILLER_28_873 ();
 FILLCELL_X1 FILLER_28_882 ();
 FILLCELL_X2 FILLER_28_900 ();
 FILLCELL_X4 FILLER_28_909 ();
 FILLCELL_X1 FILLER_28_913 ();
 FILLCELL_X32 FILLER_28_938 ();
 FILLCELL_X2 FILLER_28_970 ();
 FILLCELL_X1 FILLER_28_972 ();
 FILLCELL_X8 FILLER_28_980 ();
 FILLCELL_X2 FILLER_28_988 ();
 FILLCELL_X2 FILLER_28_997 ();
 FILLCELL_X2 FILLER_28_1016 ();
 FILLCELL_X2 FILLER_28_1083 ();
 FILLCELL_X2 FILLER_28_1109 ();
 FILLCELL_X1 FILLER_28_1111 ();
 FILLCELL_X4 FILLER_28_1119 ();
 FILLCELL_X4 FILLER_28_1130 ();
 FILLCELL_X16 FILLER_28_1158 ();
 FILLCELL_X1 FILLER_28_1174 ();
 FILLCELL_X16 FILLER_28_1188 ();
 FILLCELL_X1 FILLER_28_1204 ();
 FILLCELL_X8 FILLER_28_1232 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X16 FILLER_29_65 ();
 FILLCELL_X8 FILLER_29_81 ();
 FILLCELL_X4 FILLER_29_106 ();
 FILLCELL_X1 FILLER_29_128 ();
 FILLCELL_X2 FILLER_29_136 ();
 FILLCELL_X2 FILLER_29_145 ();
 FILLCELL_X2 FILLER_29_164 ();
 FILLCELL_X8 FILLER_29_173 ();
 FILLCELL_X1 FILLER_29_181 ();
 FILLCELL_X2 FILLER_29_185 ();
 FILLCELL_X1 FILLER_29_187 ();
 FILLCELL_X8 FILLER_29_205 ();
 FILLCELL_X2 FILLER_29_213 ();
 FILLCELL_X4 FILLER_29_239 ();
 FILLCELL_X2 FILLER_29_243 ();
 FILLCELL_X32 FILLER_29_269 ();
 FILLCELL_X32 FILLER_29_301 ();
 FILLCELL_X32 FILLER_29_333 ();
 FILLCELL_X4 FILLER_29_365 ();
 FILLCELL_X2 FILLER_29_369 ();
 FILLCELL_X1 FILLER_29_371 ();
 FILLCELL_X8 FILLER_29_389 ();
 FILLCELL_X4 FILLER_29_397 ();
 FILLCELL_X32 FILLER_29_404 ();
 FILLCELL_X32 FILLER_29_436 ();
 FILLCELL_X32 FILLER_29_468 ();
 FILLCELL_X32 FILLER_29_500 ();
 FILLCELL_X32 FILLER_29_532 ();
 FILLCELL_X32 FILLER_29_564 ();
 FILLCELL_X32 FILLER_29_596 ();
 FILLCELL_X16 FILLER_29_628 ();
 FILLCELL_X4 FILLER_29_644 ();
 FILLCELL_X8 FILLER_29_672 ();
 FILLCELL_X1 FILLER_29_680 ();
 FILLCELL_X8 FILLER_29_705 ();
 FILLCELL_X4 FILLER_29_713 ();
 FILLCELL_X2 FILLER_29_717 ();
 FILLCELL_X4 FILLER_29_744 ();
 FILLCELL_X2 FILLER_29_748 ();
 FILLCELL_X2 FILLER_29_767 ();
 FILLCELL_X1 FILLER_29_769 ();
 FILLCELL_X4 FILLER_29_787 ();
 FILLCELL_X1 FILLER_29_791 ();
 FILLCELL_X2 FILLER_29_809 ();
 FILLCELL_X2 FILLER_29_818 ();
 FILLCELL_X1 FILLER_29_820 ();
 FILLCELL_X2 FILLER_29_828 ();
 FILLCELL_X1 FILLER_29_830 ();
 FILLCELL_X1 FILLER_29_838 ();
 FILLCELL_X1 FILLER_29_848 ();
 FILLCELL_X2 FILLER_29_862 ();
 FILLCELL_X2 FILLER_29_871 ();
 FILLCELL_X4 FILLER_29_886 ();
 FILLCELL_X4 FILLER_29_897 ();
 FILLCELL_X2 FILLER_29_914 ();
 FILLCELL_X1 FILLER_29_916 ();
 FILLCELL_X8 FILLER_29_937 ();
 FILLCELL_X4 FILLER_29_945 ();
 FILLCELL_X2 FILLER_29_949 ();
 FILLCELL_X1 FILLER_29_951 ();
 FILLCELL_X8 FILLER_29_969 ();
 FILLCELL_X4 FILLER_29_977 ();
 FILLCELL_X4 FILLER_29_988 ();
 FILLCELL_X2 FILLER_29_1016 ();
 FILLCELL_X1 FILLER_29_1018 ();
 FILLCELL_X1 FILLER_29_1040 ();
 FILLCELL_X32 FILLER_29_1098 ();
 FILLCELL_X8 FILLER_29_1130 ();
 FILLCELL_X2 FILLER_29_1138 ();
 FILLCELL_X1 FILLER_29_1140 ();
 FILLCELL_X16 FILLER_29_1154 ();
 FILLCELL_X8 FILLER_29_1170 ();
 FILLCELL_X2 FILLER_29_1195 ();
 FILLCELL_X8 FILLER_29_1231 ();
 FILLCELL_X1 FILLER_29_1239 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X16 FILLER_30_65 ();
 FILLCELL_X4 FILLER_30_102 ();
 FILLCELL_X2 FILLER_30_106 ();
 FILLCELL_X1 FILLER_30_108 ();
 FILLCELL_X2 FILLER_30_116 ();
 FILLCELL_X1 FILLER_30_135 ();
 FILLCELL_X1 FILLER_30_143 ();
 FILLCELL_X1 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_169 ();
 FILLCELL_X2 FILLER_30_180 ();
 FILLCELL_X2 FILLER_30_194 ();
 FILLCELL_X1 FILLER_30_196 ();
 FILLCELL_X4 FILLER_30_214 ();
 FILLCELL_X2 FILLER_30_218 ();
 FILLCELL_X1 FILLER_30_220 ();
 FILLCELL_X4 FILLER_30_228 ();
 FILLCELL_X2 FILLER_30_232 ();
 FILLCELL_X1 FILLER_30_234 ();
 FILLCELL_X8 FILLER_30_242 ();
 FILLCELL_X2 FILLER_30_250 ();
 FILLCELL_X8 FILLER_30_274 ();
 FILLCELL_X1 FILLER_30_282 ();
 FILLCELL_X8 FILLER_30_286 ();
 FILLCELL_X4 FILLER_30_294 ();
 FILLCELL_X2 FILLER_30_298 ();
 FILLCELL_X1 FILLER_30_300 ();
 FILLCELL_X32 FILLER_30_318 ();
 FILLCELL_X16 FILLER_30_350 ();
 FILLCELL_X4 FILLER_30_366 ();
 FILLCELL_X8 FILLER_30_401 ();
 FILLCELL_X1 FILLER_30_409 ();
 FILLCELL_X16 FILLER_30_427 ();
 FILLCELL_X32 FILLER_30_484 ();
 FILLCELL_X32 FILLER_30_516 ();
 FILLCELL_X32 FILLER_30_548 ();
 FILLCELL_X32 FILLER_30_580 ();
 FILLCELL_X16 FILLER_30_612 ();
 FILLCELL_X2 FILLER_30_628 ();
 FILLCELL_X1 FILLER_30_630 ();
 FILLCELL_X8 FILLER_30_632 ();
 FILLCELL_X4 FILLER_30_640 ();
 FILLCELL_X2 FILLER_30_644 ();
 FILLCELL_X4 FILLER_30_701 ();
 FILLCELL_X2 FILLER_30_705 ();
 FILLCELL_X16 FILLER_30_712 ();
 FILLCELL_X2 FILLER_30_728 ();
 FILLCELL_X16 FILLER_30_788 ();
 FILLCELL_X4 FILLER_30_804 ();
 FILLCELL_X1 FILLER_30_808 ();
 FILLCELL_X32 FILLER_30_826 ();
 FILLCELL_X32 FILLER_30_858 ();
 FILLCELL_X32 FILLER_30_890 ();
 FILLCELL_X4 FILLER_30_922 ();
 FILLCELL_X2 FILLER_30_926 ();
 FILLCELL_X2 FILLER_30_952 ();
 FILLCELL_X16 FILLER_30_968 ();
 FILLCELL_X8 FILLER_30_984 ();
 FILLCELL_X4 FILLER_30_992 ();
 FILLCELL_X2 FILLER_30_996 ();
 FILLCELL_X4 FILLER_30_1015 ();
 FILLCELL_X2 FILLER_30_1019 ();
 FILLCELL_X1 FILLER_30_1021 ();
 FILLCELL_X4 FILLER_30_1039 ();
 FILLCELL_X2 FILLER_30_1043 ();
 FILLCELL_X1 FILLER_30_1045 ();
 FILLCELL_X4 FILLER_30_1064 ();
 FILLCELL_X16 FILLER_30_1075 ();
 FILLCELL_X1 FILLER_30_1091 ();
 FILLCELL_X4 FILLER_30_1106 ();
 FILLCELL_X2 FILLER_30_1110 ();
 FILLCELL_X1 FILLER_30_1112 ();
 FILLCELL_X8 FILLER_30_1118 ();
 FILLCELL_X4 FILLER_30_1126 ();
 FILLCELL_X16 FILLER_30_1147 ();
 FILLCELL_X1 FILLER_30_1163 ();
 FILLCELL_X2 FILLER_30_1207 ();
 FILLCELL_X1 FILLER_30_1209 ();
 FILLCELL_X16 FILLER_30_1224 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X4 FILLER_31_33 ();
 FILLCELL_X1 FILLER_31_37 ();
 FILLCELL_X8 FILLER_31_55 ();
 FILLCELL_X2 FILLER_31_63 ();
 FILLCELL_X1 FILLER_31_65 ();
 FILLCELL_X4 FILLER_31_90 ();
 FILLCELL_X2 FILLER_31_94 ();
 FILLCELL_X8 FILLER_31_100 ();
 FILLCELL_X4 FILLER_31_125 ();
 FILLCELL_X2 FILLER_31_129 ();
 FILLCELL_X1 FILLER_31_162 ();
 FILLCELL_X8 FILLER_31_170 ();
 FILLCELL_X2 FILLER_31_178 ();
 FILLCELL_X1 FILLER_31_180 ();
 FILLCELL_X16 FILLER_31_226 ();
 FILLCELL_X8 FILLER_31_242 ();
 FILLCELL_X4 FILLER_31_250 ();
 FILLCELL_X16 FILLER_31_278 ();
 FILLCELL_X8 FILLER_31_294 ();
 FILLCELL_X2 FILLER_31_302 ();
 FILLCELL_X2 FILLER_31_328 ();
 FILLCELL_X16 FILLER_31_354 ();
 FILLCELL_X2 FILLER_31_370 ();
 FILLCELL_X8 FILLER_31_403 ();
 FILLCELL_X2 FILLER_31_411 ();
 FILLCELL_X16 FILLER_31_420 ();
 FILLCELL_X4 FILLER_31_436 ();
 FILLCELL_X2 FILLER_31_478 ();
 FILLCELL_X1 FILLER_31_480 ();
 FILLCELL_X32 FILLER_31_498 ();
 FILLCELL_X32 FILLER_31_530 ();
 FILLCELL_X32 FILLER_31_562 ();
 FILLCELL_X32 FILLER_31_594 ();
 FILLCELL_X8 FILLER_31_626 ();
 FILLCELL_X2 FILLER_31_634 ();
 FILLCELL_X16 FILLER_31_674 ();
 FILLCELL_X4 FILLER_31_690 ();
 FILLCELL_X2 FILLER_31_694 ();
 FILLCELL_X1 FILLER_31_696 ();
 FILLCELL_X4 FILLER_31_704 ();
 FILLCELL_X2 FILLER_31_708 ();
 FILLCELL_X1 FILLER_31_710 ();
 FILLCELL_X1 FILLER_31_720 ();
 FILLCELL_X16 FILLER_31_737 ();
 FILLCELL_X8 FILLER_31_753 ();
 FILLCELL_X4 FILLER_31_761 ();
 FILLCELL_X1 FILLER_31_765 ();
 FILLCELL_X4 FILLER_31_773 ();
 FILLCELL_X2 FILLER_31_777 ();
 FILLCELL_X16 FILLER_31_788 ();
 FILLCELL_X4 FILLER_31_804 ();
 FILLCELL_X1 FILLER_31_808 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X8 FILLER_31_865 ();
 FILLCELL_X4 FILLER_31_873 ();
 FILLCELL_X16 FILLER_31_884 ();
 FILLCELL_X4 FILLER_31_900 ();
 FILLCELL_X1 FILLER_31_904 ();
 FILLCELL_X16 FILLER_31_929 ();
 FILLCELL_X2 FILLER_31_945 ();
 FILLCELL_X1 FILLER_31_947 ();
 FILLCELL_X2 FILLER_31_955 ();
 FILLCELL_X4 FILLER_31_973 ();
 FILLCELL_X8 FILLER_31_1008 ();
 FILLCELL_X4 FILLER_31_1016 ();
 FILLCELL_X16 FILLER_31_1037 ();
 FILLCELL_X2 FILLER_31_1053 ();
 FILLCELL_X8 FILLER_31_1079 ();
 FILLCELL_X2 FILLER_31_1087 ();
 FILLCELL_X8 FILLER_31_1113 ();
 FILLCELL_X4 FILLER_31_1121 ();
 FILLCELL_X1 FILLER_31_1125 ();
 FILLCELL_X32 FILLER_31_1133 ();
 FILLCELL_X8 FILLER_31_1165 ();
 FILLCELL_X4 FILLER_31_1173 ();
 FILLCELL_X2 FILLER_31_1177 ();
 FILLCELL_X16 FILLER_31_1196 ();
 FILLCELL_X1 FILLER_31_1212 ();
 FILLCELL_X4 FILLER_31_1220 ();
 FILLCELL_X2 FILLER_31_1224 ();
 FILLCELL_X1 FILLER_31_1226 ();
 FILLCELL_X4 FILLER_31_1230 ();
 FILLCELL_X2 FILLER_31_1234 ();
 FILLCELL_X1 FILLER_31_1239 ();
 FILLCELL_X16 FILLER_32_1 ();
 FILLCELL_X8 FILLER_32_17 ();
 FILLCELL_X2 FILLER_32_25 ();
 FILLCELL_X8 FILLER_32_34 ();
 FILLCELL_X1 FILLER_32_42 ();
 FILLCELL_X8 FILLER_32_50 ();
 FILLCELL_X2 FILLER_32_65 ();
 FILLCELL_X4 FILLER_32_98 ();
 FILLCELL_X2 FILLER_32_102 ();
 FILLCELL_X4 FILLER_32_111 ();
 FILLCELL_X1 FILLER_32_115 ();
 FILLCELL_X2 FILLER_32_123 ();
 FILLCELL_X1 FILLER_32_125 ();
 FILLCELL_X2 FILLER_32_138 ();
 FILLCELL_X1 FILLER_32_140 ();
 FILLCELL_X32 FILLER_32_148 ();
 FILLCELL_X4 FILLER_32_180 ();
 FILLCELL_X1 FILLER_32_205 ();
 FILLCELL_X4 FILLER_32_213 ();
 FILLCELL_X4 FILLER_32_248 ();
 FILLCELL_X2 FILLER_32_252 ();
 FILLCELL_X8 FILLER_32_316 ();
 FILLCELL_X2 FILLER_32_355 ();
 FILLCELL_X2 FILLER_32_365 ();
 FILLCELL_X2 FILLER_32_398 ();
 FILLCELL_X1 FILLER_32_400 ();
 FILLCELL_X2 FILLER_32_456 ();
 FILLCELL_X32 FILLER_32_473 ();
 FILLCELL_X32 FILLER_32_505 ();
 FILLCELL_X32 FILLER_32_537 ();
 FILLCELL_X32 FILLER_32_569 ();
 FILLCELL_X16 FILLER_32_601 ();
 FILLCELL_X8 FILLER_32_617 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X4 FILLER_32_632 ();
 FILLCELL_X2 FILLER_32_636 ();
 FILLCELL_X2 FILLER_32_655 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X4 FILLER_32_696 ();
 FILLCELL_X2 FILLER_32_700 ();
 FILLCELL_X16 FILLER_32_714 ();
 FILLCELL_X2 FILLER_32_730 ();
 FILLCELL_X32 FILLER_32_739 ();
 FILLCELL_X32 FILLER_32_771 ();
 FILLCELL_X16 FILLER_32_803 ();
 FILLCELL_X8 FILLER_32_819 ();
 FILLCELL_X4 FILLER_32_827 ();
 FILLCELL_X8 FILLER_32_855 ();
 FILLCELL_X4 FILLER_32_863 ();
 FILLCELL_X8 FILLER_32_898 ();
 FILLCELL_X2 FILLER_32_906 ();
 FILLCELL_X16 FILLER_32_925 ();
 FILLCELL_X2 FILLER_32_941 ();
 FILLCELL_X1 FILLER_32_943 ();
 FILLCELL_X1 FILLER_32_974 ();
 FILLCELL_X8 FILLER_32_1006 ();
 FILLCELL_X2 FILLER_32_1028 ();
 FILLCELL_X1 FILLER_32_1030 ();
 FILLCELL_X16 FILLER_32_1045 ();
 FILLCELL_X1 FILLER_32_1061 ();
 FILLCELL_X8 FILLER_32_1066 ();
 FILLCELL_X4 FILLER_32_1074 ();
 FILLCELL_X1 FILLER_32_1078 ();
 FILLCELL_X8 FILLER_32_1083 ();
 FILLCELL_X2 FILLER_32_1091 ();
 FILLCELL_X1 FILLER_32_1100 ();
 FILLCELL_X2 FILLER_32_1156 ();
 FILLCELL_X4 FILLER_32_1175 ();
 FILLCELL_X1 FILLER_32_1186 ();
 FILLCELL_X2 FILLER_32_1204 ();
 FILLCELL_X2 FILLER_32_1223 ();
 FILLCELL_X2 FILLER_32_1232 ();
 FILLCELL_X2 FILLER_32_1237 ();
 FILLCELL_X1 FILLER_32_1239 ();
 FILLCELL_X8 FILLER_33_1 ();
 FILLCELL_X4 FILLER_33_9 ();
 FILLCELL_X2 FILLER_33_13 ();
 FILLCELL_X1 FILLER_33_15 ();
 FILLCELL_X4 FILLER_33_44 ();
 FILLCELL_X8 FILLER_33_55 ();
 FILLCELL_X1 FILLER_33_63 ();
 FILLCELL_X4 FILLER_33_71 ();
 FILLCELL_X1 FILLER_33_75 ();
 FILLCELL_X2 FILLER_33_100 ();
 FILLCELL_X1 FILLER_33_102 ();
 FILLCELL_X2 FILLER_33_110 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X8 FILLER_33_161 ();
 FILLCELL_X2 FILLER_33_169 ();
 FILLCELL_X8 FILLER_33_188 ();
 FILLCELL_X16 FILLER_33_203 ();
 FILLCELL_X4 FILLER_33_219 ();
 FILLCELL_X2 FILLER_33_223 ();
 FILLCELL_X2 FILLER_33_239 ();
 FILLCELL_X4 FILLER_33_248 ();
 FILLCELL_X2 FILLER_33_252 ();
 FILLCELL_X1 FILLER_33_254 ();
 FILLCELL_X4 FILLER_33_262 ();
 FILLCELL_X2 FILLER_33_266 ();
 FILLCELL_X16 FILLER_33_275 ();
 FILLCELL_X2 FILLER_33_291 ();
 FILLCELL_X8 FILLER_33_317 ();
 FILLCELL_X4 FILLER_33_325 ();
 FILLCELL_X2 FILLER_33_329 ();
 FILLCELL_X1 FILLER_33_331 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X8 FILLER_33_385 ();
 FILLCELL_X4 FILLER_33_393 ();
 FILLCELL_X2 FILLER_33_397 ();
 FILLCELL_X4 FILLER_33_406 ();
 FILLCELL_X2 FILLER_33_410 ();
 FILLCELL_X1 FILLER_33_412 ();
 FILLCELL_X4 FILLER_33_427 ();
 FILLCELL_X1 FILLER_33_431 ();
 FILLCELL_X16 FILLER_33_439 ();
 FILLCELL_X2 FILLER_33_455 ();
 FILLCELL_X1 FILLER_33_457 ();
 FILLCELL_X32 FILLER_33_469 ();
 FILLCELL_X32 FILLER_33_501 ();
 FILLCELL_X32 FILLER_33_533 ();
 FILLCELL_X32 FILLER_33_565 ();
 FILLCELL_X32 FILLER_33_597 ();
 FILLCELL_X32 FILLER_33_629 ();
 FILLCELL_X16 FILLER_33_661 ();
 FILLCELL_X8 FILLER_33_677 ();
 FILLCELL_X4 FILLER_33_702 ();
 FILLCELL_X2 FILLER_33_706 ();
 FILLCELL_X8 FILLER_33_738 ();
 FILLCELL_X16 FILLER_33_770 ();
 FILLCELL_X4 FILLER_33_786 ();
 FILLCELL_X1 FILLER_33_790 ();
 FILLCELL_X8 FILLER_33_820 ();
 FILLCELL_X2 FILLER_33_828 ();
 FILLCELL_X4 FILLER_33_854 ();
 FILLCELL_X1 FILLER_33_858 ();
 FILLCELL_X2 FILLER_33_900 ();
 FILLCELL_X1 FILLER_33_902 ();
 FILLCELL_X1 FILLER_33_917 ();
 FILLCELL_X4 FILLER_33_949 ();
 FILLCELL_X1 FILLER_33_977 ();
 FILLCELL_X8 FILLER_33_1009 ();
 FILLCELL_X2 FILLER_33_1017 ();
 FILLCELL_X1 FILLER_33_1019 ();
 FILLCELL_X8 FILLER_33_1044 ();
 FILLCELL_X2 FILLER_33_1059 ();
 FILLCELL_X1 FILLER_33_1061 ();
 FILLCELL_X1 FILLER_33_1075 ();
 FILLCELL_X1 FILLER_33_1089 ();
 FILLCELL_X1 FILLER_33_1097 ();
 FILLCELL_X2 FILLER_33_1115 ();
 FILLCELL_X4 FILLER_33_1124 ();
 FILLCELL_X2 FILLER_33_1128 ();
 FILLCELL_X1 FILLER_33_1130 ();
 FILLCELL_X1 FILLER_33_1155 ();
 FILLCELL_X1 FILLER_33_1163 ();
 FILLCELL_X2 FILLER_33_1188 ();
 FILLCELL_X1 FILLER_33_1190 ();
 FILLCELL_X1 FILLER_33_1198 ();
 FILLCELL_X2 FILLER_33_1206 ();
 FILLCELL_X2 FILLER_33_1235 ();
 FILLCELL_X16 FILLER_34_1 ();
 FILLCELL_X8 FILLER_34_17 ();
 FILLCELL_X2 FILLER_34_25 ();
 FILLCELL_X1 FILLER_34_27 ();
 FILLCELL_X1 FILLER_34_45 ();
 FILLCELL_X2 FILLER_34_63 ();
 FILLCELL_X1 FILLER_34_72 ();
 FILLCELL_X2 FILLER_34_97 ();
 FILLCELL_X4 FILLER_34_123 ();
 FILLCELL_X1 FILLER_34_127 ();
 FILLCELL_X32 FILLER_34_149 ();
 FILLCELL_X4 FILLER_34_181 ();
 FILLCELL_X2 FILLER_34_185 ();
 FILLCELL_X1 FILLER_34_187 ();
 FILLCELL_X16 FILLER_34_195 ();
 FILLCELL_X8 FILLER_34_211 ();
 FILLCELL_X4 FILLER_34_219 ();
 FILLCELL_X1 FILLER_34_223 ();
 FILLCELL_X8 FILLER_34_250 ();
 FILLCELL_X16 FILLER_34_267 ();
 FILLCELL_X4 FILLER_34_283 ();
 FILLCELL_X2 FILLER_34_287 ();
 FILLCELL_X1 FILLER_34_289 ();
 FILLCELL_X8 FILLER_34_321 ();
 FILLCELL_X4 FILLER_34_329 ();
 FILLCELL_X8 FILLER_34_357 ();
 FILLCELL_X4 FILLER_34_365 ();
 FILLCELL_X2 FILLER_34_369 ();
 FILLCELL_X1 FILLER_34_371 ();
 FILLCELL_X32 FILLER_34_379 ();
 FILLCELL_X2 FILLER_34_411 ();
 FILLCELL_X8 FILLER_34_437 ();
 FILLCELL_X1 FILLER_34_445 ();
 FILLCELL_X1 FILLER_34_449 ();
 FILLCELL_X8 FILLER_34_457 ();
 FILLCELL_X2 FILLER_34_465 ();
 FILLCELL_X32 FILLER_34_491 ();
 FILLCELL_X32 FILLER_34_523 ();
 FILLCELL_X32 FILLER_34_555 ();
 FILLCELL_X32 FILLER_34_587 ();
 FILLCELL_X8 FILLER_34_619 ();
 FILLCELL_X4 FILLER_34_627 ();
 FILLCELL_X16 FILLER_34_632 ();
 FILLCELL_X4 FILLER_34_648 ();
 FILLCELL_X1 FILLER_34_652 ();
 FILLCELL_X16 FILLER_34_660 ();
 FILLCELL_X4 FILLER_34_676 ();
 FILLCELL_X1 FILLER_34_680 ();
 FILLCELL_X4 FILLER_34_705 ();
 FILLCELL_X2 FILLER_34_709 ();
 FILLCELL_X8 FILLER_34_766 ();
 FILLCELL_X4 FILLER_34_774 ();
 FILLCELL_X2 FILLER_34_778 ();
 FILLCELL_X2 FILLER_34_804 ();
 FILLCELL_X1 FILLER_34_826 ();
 FILLCELL_X4 FILLER_34_844 ();
 FILLCELL_X4 FILLER_34_855 ();
 FILLCELL_X8 FILLER_34_897 ();
 FILLCELL_X4 FILLER_34_905 ();
 FILLCELL_X2 FILLER_34_926 ();
 FILLCELL_X1 FILLER_34_928 ();
 FILLCELL_X4 FILLER_34_938 ();
 FILLCELL_X2 FILLER_34_942 ();
 FILLCELL_X16 FILLER_34_961 ();
 FILLCELL_X1 FILLER_34_977 ();
 FILLCELL_X16 FILLER_34_1002 ();
 FILLCELL_X8 FILLER_34_1018 ();
 FILLCELL_X1 FILLER_34_1026 ();
 FILLCELL_X4 FILLER_34_1048 ();
 FILLCELL_X2 FILLER_34_1052 ();
 FILLCELL_X1 FILLER_34_1071 ();
 FILLCELL_X16 FILLER_34_1079 ();
 FILLCELL_X16 FILLER_34_1102 ();
 FILLCELL_X1 FILLER_34_1118 ();
 FILLCELL_X8 FILLER_34_1136 ();
 FILLCELL_X4 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1155 ();
 FILLCELL_X16 FILLER_34_1187 ();
 FILLCELL_X1 FILLER_34_1203 ();
 FILLCELL_X1 FILLER_34_1235 ();
 FILLCELL_X1 FILLER_34_1239 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X8 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_48 ();
 FILLCELL_X16 FILLER_35_80 ();
 FILLCELL_X8 FILLER_35_96 ();
 FILLCELL_X4 FILLER_35_104 ();
 FILLCELL_X1 FILLER_35_125 ();
 FILLCELL_X4 FILLER_35_160 ();
 FILLCELL_X8 FILLER_35_171 ();
 FILLCELL_X4 FILLER_35_179 ();
 FILLCELL_X2 FILLER_35_183 ();
 FILLCELL_X1 FILLER_35_185 ();
 FILLCELL_X16 FILLER_35_220 ();
 FILLCELL_X8 FILLER_35_236 ();
 FILLCELL_X2 FILLER_35_244 ();
 FILLCELL_X16 FILLER_35_265 ();
 FILLCELL_X8 FILLER_35_281 ();
 FILLCELL_X4 FILLER_35_289 ();
 FILLCELL_X2 FILLER_35_293 ();
 FILLCELL_X1 FILLER_35_295 ();
 FILLCELL_X1 FILLER_35_310 ();
 FILLCELL_X8 FILLER_35_313 ();
 FILLCELL_X4 FILLER_35_321 ();
 FILLCELL_X2 FILLER_35_325 ();
 FILLCELL_X1 FILLER_35_327 ();
 FILLCELL_X32 FILLER_35_332 ();
 FILLCELL_X4 FILLER_35_364 ();
 FILLCELL_X32 FILLER_35_407 ();
 FILLCELL_X2 FILLER_35_439 ();
 FILLCELL_X4 FILLER_35_463 ();
 FILLCELL_X32 FILLER_35_498 ();
 FILLCELL_X32 FILLER_35_530 ();
 FILLCELL_X32 FILLER_35_562 ();
 FILLCELL_X32 FILLER_35_594 ();
 FILLCELL_X16 FILLER_35_626 ();
 FILLCELL_X4 FILLER_35_642 ();
 FILLCELL_X2 FILLER_35_646 ();
 FILLCELL_X1 FILLER_35_648 ();
 FILLCELL_X16 FILLER_35_666 ();
 FILLCELL_X2 FILLER_35_682 ();
 FILLCELL_X4 FILLER_35_691 ();
 FILLCELL_X2 FILLER_35_695 ();
 FILLCELL_X1 FILLER_35_697 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X16 FILLER_35_737 ();
 FILLCELL_X4 FILLER_35_753 ();
 FILLCELL_X2 FILLER_35_757 ();
 FILLCELL_X16 FILLER_35_766 ();
 FILLCELL_X4 FILLER_35_782 ();
 FILLCELL_X2 FILLER_35_786 ();
 FILLCELL_X8 FILLER_35_819 ();
 FILLCELL_X1 FILLER_35_827 ();
 FILLCELL_X32 FILLER_35_852 ();
 FILLCELL_X32 FILLER_35_884 ();
 FILLCELL_X16 FILLER_35_916 ();
 FILLCELL_X8 FILLER_35_932 ();
 FILLCELL_X8 FILLER_35_971 ();
 FILLCELL_X1 FILLER_35_986 ();
 FILLCELL_X16 FILLER_35_1001 ();
 FILLCELL_X8 FILLER_35_1017 ();
 FILLCELL_X1 FILLER_35_1025 ();
 FILLCELL_X8 FILLER_35_1044 ();
 FILLCELL_X1 FILLER_35_1052 ();
 FILLCELL_X1 FILLER_35_1089 ();
 FILLCELL_X2 FILLER_35_1097 ();
 FILLCELL_X8 FILLER_35_1106 ();
 FILLCELL_X4 FILLER_35_1114 ();
 FILLCELL_X2 FILLER_35_1118 ();
 FILLCELL_X1 FILLER_35_1127 ();
 FILLCELL_X32 FILLER_35_1145 ();
 FILLCELL_X8 FILLER_35_1228 ();
 FILLCELL_X4 FILLER_35_1236 ();
 FILLCELL_X16 FILLER_36_1 ();
 FILLCELL_X1 FILLER_36_17 ();
 FILLCELL_X8 FILLER_36_22 ();
 FILLCELL_X4 FILLER_36_30 ();
 FILLCELL_X32 FILLER_36_48 ();
 FILLCELL_X16 FILLER_36_80 ();
 FILLCELL_X8 FILLER_36_96 ();
 FILLCELL_X4 FILLER_36_104 ();
 FILLCELL_X1 FILLER_36_108 ();
 FILLCELL_X4 FILLER_36_116 ();
 FILLCELL_X2 FILLER_36_120 ();
 FILLCELL_X8 FILLER_36_129 ();
 FILLCELL_X4 FILLER_36_144 ();
 FILLCELL_X8 FILLER_36_155 ();
 FILLCELL_X1 FILLER_36_180 ();
 FILLCELL_X4 FILLER_36_195 ();
 FILLCELL_X2 FILLER_36_199 ();
 FILLCELL_X8 FILLER_36_208 ();
 FILLCELL_X1 FILLER_36_216 ();
 FILLCELL_X8 FILLER_36_234 ();
 FILLCELL_X2 FILLER_36_249 ();
 FILLCELL_X16 FILLER_36_277 ();
 FILLCELL_X8 FILLER_36_293 ();
 FILLCELL_X2 FILLER_36_301 ();
 FILLCELL_X8 FILLER_36_325 ();
 FILLCELL_X4 FILLER_36_333 ();
 FILLCELL_X2 FILLER_36_337 ();
 FILLCELL_X1 FILLER_36_339 ();
 FILLCELL_X4 FILLER_36_364 ();
 FILLCELL_X1 FILLER_36_368 ();
 FILLCELL_X8 FILLER_36_373 ();
 FILLCELL_X1 FILLER_36_381 ();
 FILLCELL_X1 FILLER_36_413 ();
 FILLCELL_X8 FILLER_36_431 ();
 FILLCELL_X32 FILLER_36_463 ();
 FILLCELL_X16 FILLER_36_495 ();
 FILLCELL_X8 FILLER_36_511 ();
 FILLCELL_X32 FILLER_36_543 ();
 FILLCELL_X32 FILLER_36_575 ();
 FILLCELL_X16 FILLER_36_607 ();
 FILLCELL_X8 FILLER_36_623 ();
 FILLCELL_X8 FILLER_36_675 ();
 FILLCELL_X16 FILLER_36_703 ();
 FILLCELL_X4 FILLER_36_719 ();
 FILLCELL_X1 FILLER_36_723 ();
 FILLCELL_X2 FILLER_36_741 ();
 FILLCELL_X4 FILLER_36_748 ();
 FILLCELL_X2 FILLER_36_752 ();
 FILLCELL_X2 FILLER_36_761 ();
 FILLCELL_X1 FILLER_36_763 ();
 FILLCELL_X16 FILLER_36_771 ();
 FILLCELL_X4 FILLER_36_787 ();
 FILLCELL_X1 FILLER_36_791 ();
 FILLCELL_X2 FILLER_36_799 ();
 FILLCELL_X16 FILLER_36_808 ();
 FILLCELL_X4 FILLER_36_824 ();
 FILLCELL_X2 FILLER_36_828 ();
 FILLCELL_X4 FILLER_36_837 ();
 FILLCELL_X2 FILLER_36_841 ();
 FILLCELL_X1 FILLER_36_843 ();
 FILLCELL_X32 FILLER_36_851 ();
 FILLCELL_X16 FILLER_36_883 ();
 FILLCELL_X4 FILLER_36_899 ();
 FILLCELL_X1 FILLER_36_903 ();
 FILLCELL_X16 FILLER_36_922 ();
 FILLCELL_X4 FILLER_36_938 ();
 FILLCELL_X2 FILLER_36_942 ();
 FILLCELL_X4 FILLER_36_951 ();
 FILLCELL_X32 FILLER_36_962 ();
 FILLCELL_X1 FILLER_36_994 ();
 FILLCELL_X16 FILLER_36_1002 ();
 FILLCELL_X1 FILLER_36_1018 ();
 FILLCELL_X8 FILLER_36_1045 ();
 FILLCELL_X4 FILLER_36_1053 ();
 FILLCELL_X1 FILLER_36_1057 ();
 FILLCELL_X2 FILLER_36_1061 ();
 FILLCELL_X2 FILLER_36_1100 ();
 FILLCELL_X1 FILLER_36_1102 ();
 FILLCELL_X4 FILLER_36_1127 ();
 FILLCELL_X2 FILLER_36_1131 ();
 FILLCELL_X16 FILLER_36_1147 ();
 FILLCELL_X2 FILLER_36_1163 ();
 FILLCELL_X1 FILLER_36_1165 ();
 FILLCELL_X8 FILLER_36_1174 ();
 FILLCELL_X2 FILLER_36_1182 ();
 FILLCELL_X1 FILLER_36_1184 ();
 FILLCELL_X2 FILLER_36_1216 ();
 FILLCELL_X8 FILLER_36_1227 ();
 FILLCELL_X4 FILLER_36_1235 ();
 FILLCELL_X1 FILLER_36_1239 ();
 FILLCELL_X16 FILLER_37_1 ();
 FILLCELL_X8 FILLER_37_17 ();
 FILLCELL_X4 FILLER_37_25 ();
 FILLCELL_X2 FILLER_37_53 ();
 FILLCELL_X16 FILLER_37_94 ();
 FILLCELL_X2 FILLER_37_110 ();
 FILLCELL_X32 FILLER_37_116 ();
 FILLCELL_X2 FILLER_37_148 ();
 FILLCELL_X1 FILLER_37_150 ();
 FILLCELL_X16 FILLER_37_168 ();
 FILLCELL_X4 FILLER_37_184 ();
 FILLCELL_X1 FILLER_37_188 ();
 FILLCELL_X8 FILLER_37_211 ();
 FILLCELL_X4 FILLER_37_236 ();
 FILLCELL_X1 FILLER_37_240 ();
 FILLCELL_X16 FILLER_37_282 ();
 FILLCELL_X4 FILLER_37_298 ();
 FILLCELL_X1 FILLER_37_302 ();
 FILLCELL_X16 FILLER_37_324 ();
 FILLCELL_X2 FILLER_37_340 ();
 FILLCELL_X1 FILLER_37_342 ();
 FILLCELL_X2 FILLER_37_388 ();
 FILLCELL_X1 FILLER_37_390 ();
 FILLCELL_X1 FILLER_37_398 ();
 FILLCELL_X4 FILLER_37_416 ();
 FILLCELL_X1 FILLER_37_420 ();
 FILLCELL_X4 FILLER_37_438 ();
 FILLCELL_X1 FILLER_37_442 ();
 FILLCELL_X2 FILLER_37_450 ();
 FILLCELL_X1 FILLER_37_452 ();
 FILLCELL_X16 FILLER_37_470 ();
 FILLCELL_X8 FILLER_37_486 ();
 FILLCELL_X2 FILLER_37_494 ();
 FILLCELL_X8 FILLER_37_527 ();
 FILLCELL_X32 FILLER_37_552 ();
 FILLCELL_X32 FILLER_37_584 ();
 FILLCELL_X4 FILLER_37_616 ();
 FILLCELL_X2 FILLER_37_620 ();
 FILLCELL_X1 FILLER_37_622 ();
 FILLCELL_X4 FILLER_37_640 ();
 FILLCELL_X2 FILLER_37_644 ();
 FILLCELL_X1 FILLER_37_646 ();
 FILLCELL_X2 FILLER_37_654 ();
 FILLCELL_X1 FILLER_37_656 ();
 FILLCELL_X8 FILLER_37_664 ();
 FILLCELL_X2 FILLER_37_672 ();
 FILLCELL_X2 FILLER_37_705 ();
 FILLCELL_X2 FILLER_37_724 ();
 FILLCELL_X1 FILLER_37_726 ();
 FILLCELL_X1 FILLER_37_734 ();
 FILLCELL_X2 FILLER_37_742 ();
 FILLCELL_X1 FILLER_37_744 ();
 FILLCELL_X2 FILLER_37_762 ();
 FILLCELL_X1 FILLER_37_764 ();
 FILLCELL_X8 FILLER_37_782 ();
 FILLCELL_X2 FILLER_37_790 ();
 FILLCELL_X1 FILLER_37_792 ();
 FILLCELL_X16 FILLER_37_800 ();
 FILLCELL_X8 FILLER_37_816 ();
 FILLCELL_X4 FILLER_37_824 ();
 FILLCELL_X2 FILLER_37_828 ();
 FILLCELL_X1 FILLER_37_830 ();
 FILLCELL_X2 FILLER_37_842 ();
 FILLCELL_X1 FILLER_37_848 ();
 FILLCELL_X1 FILLER_37_856 ();
 FILLCELL_X8 FILLER_37_864 ();
 FILLCELL_X2 FILLER_37_872 ();
 FILLCELL_X2 FILLER_37_898 ();
 FILLCELL_X1 FILLER_37_900 ();
 FILLCELL_X2 FILLER_37_931 ();
 FILLCELL_X1 FILLER_37_938 ();
 FILLCELL_X16 FILLER_37_956 ();
 FILLCELL_X4 FILLER_37_972 ();
 FILLCELL_X1 FILLER_37_976 ();
 FILLCELL_X8 FILLER_37_1001 ();
 FILLCELL_X2 FILLER_37_1009 ();
 FILLCELL_X1 FILLER_37_1011 ();
 FILLCELL_X8 FILLER_37_1053 ();
 FILLCELL_X4 FILLER_37_1061 ();
 FILLCELL_X2 FILLER_37_1065 ();
 FILLCELL_X4 FILLER_37_1101 ();
 FILLCELL_X8 FILLER_37_1156 ();
 FILLCELL_X1 FILLER_37_1164 ();
 FILLCELL_X1 FILLER_37_1189 ();
 FILLCELL_X8 FILLER_37_1199 ();
 FILLCELL_X2 FILLER_37_1219 ();
 FILLCELL_X2 FILLER_37_1228 ();
 FILLCELL_X1 FILLER_37_1230 ();
 FILLCELL_X2 FILLER_37_1234 ();
 FILLCELL_X1 FILLER_37_1236 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X8 FILLER_38_17 ();
 FILLCELL_X4 FILLER_38_25 ();
 FILLCELL_X2 FILLER_38_29 ();
 FILLCELL_X1 FILLER_38_31 ();
 FILLCELL_X8 FILLER_38_56 ();
 FILLCELL_X4 FILLER_38_64 ();
 FILLCELL_X1 FILLER_38_68 ();
 FILLCELL_X4 FILLER_38_100 ();
 FILLCELL_X1 FILLER_38_104 ();
 FILLCELL_X32 FILLER_38_146 ();
 FILLCELL_X32 FILLER_38_178 ();
 FILLCELL_X2 FILLER_38_210 ();
 FILLCELL_X1 FILLER_38_212 ();
 FILLCELL_X8 FILLER_38_234 ();
 FILLCELL_X2 FILLER_38_242 ();
 FILLCELL_X1 FILLER_38_244 ();
 FILLCELL_X8 FILLER_38_292 ();
 FILLCELL_X4 FILLER_38_300 ();
 FILLCELL_X2 FILLER_38_304 ();
 FILLCELL_X4 FILLER_38_323 ();
 FILLCELL_X2 FILLER_38_327 ();
 FILLCELL_X2 FILLER_38_377 ();
 FILLCELL_X16 FILLER_38_386 ();
 FILLCELL_X4 FILLER_38_402 ();
 FILLCELL_X8 FILLER_38_420 ();
 FILLCELL_X4 FILLER_38_428 ();
 FILLCELL_X1 FILLER_38_432 ();
 FILLCELL_X16 FILLER_38_471 ();
 FILLCELL_X4 FILLER_38_494 ();
 FILLCELL_X2 FILLER_38_498 ();
 FILLCELL_X1 FILLER_38_500 ();
 FILLCELL_X2 FILLER_38_515 ();
 FILLCELL_X1 FILLER_38_517 ();
 FILLCELL_X4 FILLER_38_532 ();
 FILLCELL_X1 FILLER_38_536 ();
 FILLCELL_X32 FILLER_38_554 ();
 FILLCELL_X32 FILLER_38_586 ();
 FILLCELL_X8 FILLER_38_618 ();
 FILLCELL_X4 FILLER_38_626 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X8 FILLER_38_632 ();
 FILLCELL_X4 FILLER_38_640 ();
 FILLCELL_X1 FILLER_38_644 ();
 FILLCELL_X1 FILLER_38_662 ();
 FILLCELL_X4 FILLER_38_692 ();
 FILLCELL_X2 FILLER_38_696 ();
 FILLCELL_X1 FILLER_38_707 ();
 FILLCELL_X4 FILLER_38_730 ();
 FILLCELL_X1 FILLER_38_741 ();
 FILLCELL_X8 FILLER_38_747 ();
 FILLCELL_X2 FILLER_38_755 ();
 FILLCELL_X1 FILLER_38_762 ();
 FILLCELL_X4 FILLER_38_783 ();
 FILLCELL_X2 FILLER_38_787 ();
 FILLCELL_X8 FILLER_38_813 ();
 FILLCELL_X4 FILLER_38_821 ();
 FILLCELL_X4 FILLER_38_851 ();
 FILLCELL_X2 FILLER_38_872 ();
 FILLCELL_X1 FILLER_38_891 ();
 FILLCELL_X8 FILLER_38_899 ();
 FILLCELL_X4 FILLER_38_921 ();
 FILLCELL_X4 FILLER_38_932 ();
 FILLCELL_X1 FILLER_38_960 ();
 FILLCELL_X2 FILLER_38_978 ();
 FILLCELL_X1 FILLER_38_987 ();
 FILLCELL_X1 FILLER_38_1005 ();
 FILLCELL_X1 FILLER_38_1023 ();
 FILLCELL_X1 FILLER_38_1031 ();
 FILLCELL_X1 FILLER_38_1046 ();
 FILLCELL_X8 FILLER_38_1051 ();
 FILLCELL_X4 FILLER_38_1059 ();
 FILLCELL_X4 FILLER_38_1070 ();
 FILLCELL_X2 FILLER_38_1074 ();
 FILLCELL_X16 FILLER_38_1103 ();
 FILLCELL_X1 FILLER_38_1119 ();
 FILLCELL_X16 FILLER_38_1129 ();
 FILLCELL_X8 FILLER_38_1145 ();
 FILLCELL_X2 FILLER_38_1153 ();
 FILLCELL_X1 FILLER_38_1155 ();
 FILLCELL_X8 FILLER_38_1173 ();
 FILLCELL_X2 FILLER_38_1181 ();
 FILLCELL_X16 FILLER_38_1190 ();
 FILLCELL_X1 FILLER_38_1206 ();
 FILLCELL_X2 FILLER_38_1237 ();
 FILLCELL_X1 FILLER_38_1239 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X8 FILLER_39_17 ();
 FILLCELL_X4 FILLER_39_25 ();
 FILLCELL_X2 FILLER_39_29 ();
 FILLCELL_X16 FILLER_39_48 ();
 FILLCELL_X4 FILLER_39_64 ();
 FILLCELL_X8 FILLER_39_85 ();
 FILLCELL_X8 FILLER_39_104 ();
 FILLCELL_X2 FILLER_39_112 ();
 FILLCELL_X1 FILLER_39_165 ();
 FILLCELL_X8 FILLER_39_173 ();
 FILLCELL_X2 FILLER_39_181 ();
 FILLCELL_X1 FILLER_39_183 ();
 FILLCELL_X32 FILLER_39_201 ();
 FILLCELL_X32 FILLER_39_233 ();
 FILLCELL_X16 FILLER_39_265 ();
 FILLCELL_X8 FILLER_39_281 ();
 FILLCELL_X2 FILLER_39_289 ();
 FILLCELL_X1 FILLER_39_291 ();
 FILLCELL_X1 FILLER_39_309 ();
 FILLCELL_X4 FILLER_39_324 ();
 FILLCELL_X2 FILLER_39_328 ();
 FILLCELL_X1 FILLER_39_330 ();
 FILLCELL_X1 FILLER_39_379 ();
 FILLCELL_X16 FILLER_39_387 ();
 FILLCELL_X8 FILLER_39_403 ();
 FILLCELL_X4 FILLER_39_411 ();
 FILLCELL_X1 FILLER_39_415 ();
 FILLCELL_X2 FILLER_39_425 ();
 FILLCELL_X16 FILLER_39_436 ();
 FILLCELL_X4 FILLER_39_452 ();
 FILLCELL_X1 FILLER_39_456 ();
 FILLCELL_X2 FILLER_39_464 ();
 FILLCELL_X1 FILLER_39_466 ();
 FILLCELL_X8 FILLER_39_471 ();
 FILLCELL_X4 FILLER_39_479 ();
 FILLCELL_X2 FILLER_39_483 ();
 FILLCELL_X8 FILLER_39_519 ();
 FILLCELL_X4 FILLER_39_527 ();
 FILLCELL_X2 FILLER_39_531 ();
 FILLCELL_X1 FILLER_39_533 ();
 FILLCELL_X32 FILLER_39_555 ();
 FILLCELL_X32 FILLER_39_587 ();
 FILLCELL_X16 FILLER_39_619 ();
 FILLCELL_X1 FILLER_39_635 ();
 FILLCELL_X2 FILLER_39_660 ();
 FILLCELL_X8 FILLER_39_693 ();
 FILLCELL_X2 FILLER_39_734 ();
 FILLCELL_X1 FILLER_39_736 ();
 FILLCELL_X1 FILLER_39_777 ();
 FILLCELL_X4 FILLER_39_819 ();
 FILLCELL_X4 FILLER_39_840 ();
 FILLCELL_X1 FILLER_39_844 ();
 FILLCELL_X1 FILLER_39_869 ();
 FILLCELL_X8 FILLER_39_877 ();
 FILLCELL_X4 FILLER_39_885 ();
 FILLCELL_X4 FILLER_39_896 ();
 FILLCELL_X2 FILLER_39_900 ();
 FILLCELL_X1 FILLER_39_943 ();
 FILLCELL_X1 FILLER_39_958 ();
 FILLCELL_X2 FILLER_39_966 ();
 FILLCELL_X2 FILLER_39_985 ();
 FILLCELL_X8 FILLER_39_999 ();
 FILLCELL_X1 FILLER_39_1007 ();
 FILLCELL_X4 FILLER_39_1022 ();
 FILLCELL_X2 FILLER_39_1026 ();
 FILLCELL_X4 FILLER_39_1041 ();
 FILLCELL_X1 FILLER_39_1045 ();
 FILLCELL_X16 FILLER_39_1103 ();
 FILLCELL_X4 FILLER_39_1119 ();
 FILLCELL_X2 FILLER_39_1123 ();
 FILLCELL_X1 FILLER_39_1125 ();
 FILLCELL_X16 FILLER_39_1139 ();
 FILLCELL_X4 FILLER_39_1155 ();
 FILLCELL_X1 FILLER_39_1173 ();
 FILLCELL_X2 FILLER_39_1181 ();
 FILLCELL_X4 FILLER_39_1200 ();
 FILLCELL_X4 FILLER_39_1211 ();
 FILLCELL_X2 FILLER_39_1215 ();
 FILLCELL_X4 FILLER_39_1234 ();
 FILLCELL_X2 FILLER_39_1238 ();
 FILLCELL_X8 FILLER_40_1 ();
 FILLCELL_X4 FILLER_40_9 ();
 FILLCELL_X8 FILLER_40_17 ();
 FILLCELL_X2 FILLER_40_25 ();
 FILLCELL_X4 FILLER_40_34 ();
 FILLCELL_X4 FILLER_40_45 ();
 FILLCELL_X2 FILLER_40_49 ();
 FILLCELL_X8 FILLER_40_58 ();
 FILLCELL_X1 FILLER_40_66 ();
 FILLCELL_X1 FILLER_40_98 ();
 FILLCELL_X2 FILLER_40_123 ();
 FILLCELL_X1 FILLER_40_125 ();
 FILLCELL_X2 FILLER_40_138 ();
 FILLCELL_X1 FILLER_40_147 ();
 FILLCELL_X4 FILLER_40_155 ();
 FILLCELL_X4 FILLER_40_166 ();
 FILLCELL_X2 FILLER_40_170 ();
 FILLCELL_X4 FILLER_40_196 ();
 FILLCELL_X2 FILLER_40_200 ();
 FILLCELL_X16 FILLER_40_209 ();
 FILLCELL_X4 FILLER_40_225 ();
 FILLCELL_X2 FILLER_40_229 ();
 FILLCELL_X1 FILLER_40_231 ();
 FILLCELL_X32 FILLER_40_239 ();
 FILLCELL_X8 FILLER_40_271 ();
 FILLCELL_X1 FILLER_40_279 ();
 FILLCELL_X32 FILLER_40_311 ();
 FILLCELL_X4 FILLER_40_343 ();
 FILLCELL_X1 FILLER_40_356 ();
 FILLCELL_X4 FILLER_40_369 ();
 FILLCELL_X2 FILLER_40_373 ();
 FILLCELL_X1 FILLER_40_375 ();
 FILLCELL_X16 FILLER_40_383 ();
 FILLCELL_X4 FILLER_40_399 ();
 FILLCELL_X1 FILLER_40_403 ();
 FILLCELL_X2 FILLER_40_411 ();
 FILLCELL_X1 FILLER_40_413 ();
 FILLCELL_X4 FILLER_40_423 ();
 FILLCELL_X16 FILLER_40_445 ();
 FILLCELL_X4 FILLER_40_461 ();
 FILLCELL_X2 FILLER_40_465 ();
 FILLCELL_X16 FILLER_40_479 ();
 FILLCELL_X32 FILLER_40_502 ();
 FILLCELL_X32 FILLER_40_534 ();
 FILLCELL_X32 FILLER_40_566 ();
 FILLCELL_X32 FILLER_40_598 ();
 FILLCELL_X1 FILLER_40_630 ();
 FILLCELL_X4 FILLER_40_632 ();
 FILLCELL_X2 FILLER_40_636 ();
 FILLCELL_X32 FILLER_40_662 ();
 FILLCELL_X8 FILLER_40_694 ();
 FILLCELL_X4 FILLER_40_702 ();
 FILLCELL_X2 FILLER_40_706 ();
 FILLCELL_X1 FILLER_40_708 ();
 FILLCELL_X1 FILLER_40_711 ();
 FILLCELL_X4 FILLER_40_715 ();
 FILLCELL_X8 FILLER_40_729 ();
 FILLCELL_X2 FILLER_40_737 ();
 FILLCELL_X16 FILLER_40_744 ();
 FILLCELL_X1 FILLER_40_760 ();
 FILLCELL_X2 FILLER_40_764 ();
 FILLCELL_X1 FILLER_40_766 ();
 FILLCELL_X1 FILLER_40_815 ();
 FILLCELL_X16 FILLER_40_840 ();
 FILLCELL_X8 FILLER_40_856 ();
 FILLCELL_X4 FILLER_40_864 ();
 FILLCELL_X16 FILLER_40_875 ();
 FILLCELL_X4 FILLER_40_891 ();
 FILLCELL_X1 FILLER_40_895 ();
 FILLCELL_X16 FILLER_40_920 ();
 FILLCELL_X4 FILLER_40_936 ();
 FILLCELL_X1 FILLER_40_940 ();
 FILLCELL_X4 FILLER_40_958 ();
 FILLCELL_X2 FILLER_40_969 ();
 FILLCELL_X1 FILLER_40_971 ();
 FILLCELL_X1 FILLER_40_979 ();
 FILLCELL_X1 FILLER_40_983 ();
 FILLCELL_X8 FILLER_40_991 ();
 FILLCELL_X2 FILLER_40_999 ();
 FILLCELL_X1 FILLER_40_1001 ();
 FILLCELL_X16 FILLER_40_1016 ();
 FILLCELL_X4 FILLER_40_1032 ();
 FILLCELL_X2 FILLER_40_1036 ();
 FILLCELL_X2 FILLER_40_1045 ();
 FILLCELL_X1 FILLER_40_1064 ();
 FILLCELL_X2 FILLER_40_1082 ();
 FILLCELL_X16 FILLER_40_1106 ();
 FILLCELL_X8 FILLER_40_1122 ();
 FILLCELL_X1 FILLER_40_1130 ();
 FILLCELL_X4 FILLER_40_1148 ();
 FILLCELL_X2 FILLER_40_1152 ();
 FILLCELL_X4 FILLER_40_1187 ();
 FILLCELL_X2 FILLER_40_1191 ();
 FILLCELL_X2 FILLER_40_1217 ();
 FILLCELL_X4 FILLER_40_1226 ();
 FILLCELL_X4 FILLER_40_1233 ();
 FILLCELL_X2 FILLER_40_1237 ();
 FILLCELL_X1 FILLER_40_1239 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X4 FILLER_41_33 ();
 FILLCELL_X1 FILLER_41_37 ();
 FILLCELL_X32 FILLER_41_55 ();
 FILLCELL_X2 FILLER_41_87 ();
 FILLCELL_X32 FILLER_41_96 ();
 FILLCELL_X16 FILLER_41_128 ();
 FILLCELL_X8 FILLER_41_144 ();
 FILLCELL_X4 FILLER_41_152 ();
 FILLCELL_X2 FILLER_41_156 ();
 FILLCELL_X1 FILLER_41_158 ();
 FILLCELL_X4 FILLER_41_176 ();
 FILLCELL_X4 FILLER_41_187 ();
 FILLCELL_X2 FILLER_41_191 ();
 FILLCELL_X1 FILLER_41_193 ();
 FILLCELL_X2 FILLER_41_201 ();
 FILLCELL_X1 FILLER_41_203 ();
 FILLCELL_X32 FILLER_41_249 ();
 FILLCELL_X32 FILLER_41_281 ();
 FILLCELL_X2 FILLER_41_313 ();
 FILLCELL_X32 FILLER_41_318 ();
 FILLCELL_X4 FILLER_41_350 ();
 FILLCELL_X2 FILLER_41_354 ();
 FILLCELL_X1 FILLER_41_356 ();
 FILLCELL_X4 FILLER_41_386 ();
 FILLCELL_X2 FILLER_41_397 ();
 FILLCELL_X2 FILLER_41_416 ();
 FILLCELL_X1 FILLER_41_418 ();
 FILLCELL_X2 FILLER_41_428 ();
 FILLCELL_X1 FILLER_41_430 ();
 FILLCELL_X8 FILLER_41_448 ();
 FILLCELL_X2 FILLER_41_456 ();
 FILLCELL_X1 FILLER_41_458 ();
 FILLCELL_X4 FILLER_41_476 ();
 FILLCELL_X8 FILLER_41_487 ();
 FILLCELL_X4 FILLER_41_536 ();
 FILLCELL_X2 FILLER_41_540 ();
 FILLCELL_X32 FILLER_41_559 ();
 FILLCELL_X32 FILLER_41_591 ();
 FILLCELL_X16 FILLER_41_623 ();
 FILLCELL_X4 FILLER_41_639 ();
 FILLCELL_X32 FILLER_41_650 ();
 FILLCELL_X8 FILLER_41_689 ();
 FILLCELL_X4 FILLER_41_697 ();
 FILLCELL_X2 FILLER_41_701 ();
 FILLCELL_X1 FILLER_41_703 ();
 FILLCELL_X32 FILLER_41_734 ();
 FILLCELL_X16 FILLER_41_766 ();
 FILLCELL_X4 FILLER_41_782 ();
 FILLCELL_X4 FILLER_41_793 ();
 FILLCELL_X2 FILLER_41_797 ();
 FILLCELL_X8 FILLER_41_814 ();
 FILLCELL_X2 FILLER_41_822 ();
 FILLCELL_X32 FILLER_41_850 ();
 FILLCELL_X16 FILLER_41_882 ();
 FILLCELL_X8 FILLER_41_898 ();
 FILLCELL_X4 FILLER_41_906 ();
 FILLCELL_X2 FILLER_41_910 ();
 FILLCELL_X32 FILLER_41_923 ();
 FILLCELL_X32 FILLER_41_955 ();
 FILLCELL_X16 FILLER_41_987 ();
 FILLCELL_X2 FILLER_41_1003 ();
 FILLCELL_X1 FILLER_41_1005 ();
 FILLCELL_X8 FILLER_41_1018 ();
 FILLCELL_X1 FILLER_41_1033 ();
 FILLCELL_X8 FILLER_41_1058 ();
 FILLCELL_X2 FILLER_41_1066 ();
 FILLCELL_X1 FILLER_41_1068 ();
 FILLCELL_X2 FILLER_41_1090 ();
 FILLCELL_X4 FILLER_41_1123 ();
 FILLCELL_X2 FILLER_41_1127 ();
 FILLCELL_X32 FILLER_41_1146 ();
 FILLCELL_X16 FILLER_41_1178 ();
 FILLCELL_X8 FILLER_41_1194 ();
 FILLCELL_X2 FILLER_41_1202 ();
 FILLCELL_X1 FILLER_41_1233 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X8 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_48 ();
 FILLCELL_X8 FILLER_42_80 ();
 FILLCELL_X4 FILLER_42_88 ();
 FILLCELL_X2 FILLER_42_92 ();
 FILLCELL_X1 FILLER_42_94 ();
 FILLCELL_X1 FILLER_42_119 ();
 FILLCELL_X4 FILLER_42_127 ();
 FILLCELL_X1 FILLER_42_131 ();
 FILLCELL_X8 FILLER_42_139 ();
 FILLCELL_X16 FILLER_42_154 ();
 FILLCELL_X8 FILLER_42_170 ();
 FILLCELL_X4 FILLER_42_178 ();
 FILLCELL_X1 FILLER_42_231 ();
 FILLCELL_X2 FILLER_42_239 ();
 FILLCELL_X2 FILLER_42_250 ();
 FILLCELL_X2 FILLER_42_259 ();
 FILLCELL_X2 FILLER_42_268 ();
 FILLCELL_X16 FILLER_42_292 ();
 FILLCELL_X2 FILLER_42_308 ();
 FILLCELL_X8 FILLER_42_317 ();
 FILLCELL_X2 FILLER_42_325 ();
 FILLCELL_X1 FILLER_42_327 ();
 FILLCELL_X16 FILLER_42_345 ();
 FILLCELL_X1 FILLER_42_361 ();
 FILLCELL_X1 FILLER_42_427 ();
 FILLCELL_X2 FILLER_42_435 ();
 FILLCELL_X1 FILLER_42_437 ();
 FILLCELL_X2 FILLER_42_445 ();
 FILLCELL_X1 FILLER_42_447 ();
 FILLCELL_X1 FILLER_42_479 ();
 FILLCELL_X2 FILLER_42_497 ();
 FILLCELL_X2 FILLER_42_516 ();
 FILLCELL_X2 FILLER_42_535 ();
 FILLCELL_X1 FILLER_42_537 ();
 FILLCELL_X32 FILLER_42_562 ();
 FILLCELL_X32 FILLER_42_594 ();
 FILLCELL_X4 FILLER_42_626 ();
 FILLCELL_X1 FILLER_42_630 ();
 FILLCELL_X4 FILLER_42_632 ();
 FILLCELL_X8 FILLER_42_660 ();
 FILLCELL_X4 FILLER_42_668 ();
 FILLCELL_X2 FILLER_42_672 ();
 FILLCELL_X1 FILLER_42_674 ();
 FILLCELL_X4 FILLER_42_692 ();
 FILLCELL_X1 FILLER_42_696 ();
 FILLCELL_X4 FILLER_42_739 ();
 FILLCELL_X16 FILLER_42_763 ();
 FILLCELL_X1 FILLER_42_779 ();
 FILLCELL_X4 FILLER_42_804 ();
 FILLCELL_X2 FILLER_42_808 ();
 FILLCELL_X1 FILLER_42_810 ();
 FILLCELL_X16 FILLER_42_820 ();
 FILLCELL_X8 FILLER_42_836 ();
 FILLCELL_X4 FILLER_42_844 ();
 FILLCELL_X2 FILLER_42_848 ();
 FILLCELL_X1 FILLER_42_850 ();
 FILLCELL_X4 FILLER_42_875 ();
 FILLCELL_X4 FILLER_42_886 ();
 FILLCELL_X8 FILLER_42_897 ();
 FILLCELL_X4 FILLER_42_918 ();
 FILLCELL_X1 FILLER_42_926 ();
 FILLCELL_X2 FILLER_42_941 ();
 FILLCELL_X1 FILLER_42_943 ();
 FILLCELL_X1 FILLER_42_950 ();
 FILLCELL_X4 FILLER_42_965 ();
 FILLCELL_X2 FILLER_42_969 ();
 FILLCELL_X1 FILLER_42_981 ();
 FILLCELL_X2 FILLER_42_1013 ();
 FILLCELL_X1 FILLER_42_1015 ();
 FILLCELL_X4 FILLER_42_1033 ();
 FILLCELL_X2 FILLER_42_1037 ();
 FILLCELL_X1 FILLER_42_1039 ();
 FILLCELL_X4 FILLER_42_1054 ();
 FILLCELL_X4 FILLER_42_1062 ();
 FILLCELL_X16 FILLER_42_1074 ();
 FILLCELL_X1 FILLER_42_1090 ();
 FILLCELL_X1 FILLER_42_1131 ();
 FILLCELL_X16 FILLER_42_1150 ();
 FILLCELL_X8 FILLER_42_1166 ();
 FILLCELL_X1 FILLER_42_1174 ();
 FILLCELL_X16 FILLER_42_1189 ();
 FILLCELL_X4 FILLER_42_1205 ();
 FILLCELL_X1 FILLER_42_1216 ();
 FILLCELL_X4 FILLER_42_1234 ();
 FILLCELL_X2 FILLER_42_1238 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X2 FILLER_43_33 ();
 FILLCELL_X1 FILLER_43_35 ();
 FILLCELL_X4 FILLER_43_84 ();
 FILLCELL_X1 FILLER_43_100 ();
 FILLCELL_X2 FILLER_43_108 ();
 FILLCELL_X1 FILLER_43_110 ();
 FILLCELL_X2 FILLER_43_145 ();
 FILLCELL_X1 FILLER_43_164 ();
 FILLCELL_X8 FILLER_43_172 ();
 FILLCELL_X2 FILLER_43_180 ();
 FILLCELL_X32 FILLER_43_198 ();
 FILLCELL_X16 FILLER_43_230 ();
 FILLCELL_X2 FILLER_43_246 ();
 FILLCELL_X2 FILLER_43_323 ();
 FILLCELL_X1 FILLER_43_325 ();
 FILLCELL_X32 FILLER_43_357 ();
 FILLCELL_X4 FILLER_43_389 ();
 FILLCELL_X2 FILLER_43_393 ();
 FILLCELL_X1 FILLER_43_402 ();
 FILLCELL_X8 FILLER_43_417 ();
 FILLCELL_X1 FILLER_43_425 ();
 FILLCELL_X4 FILLER_43_467 ();
 FILLCELL_X2 FILLER_43_471 ();
 FILLCELL_X2 FILLER_43_480 ();
 FILLCELL_X1 FILLER_43_482 ();
 FILLCELL_X1 FILLER_43_490 ();
 FILLCELL_X1 FILLER_43_505 ();
 FILLCELL_X2 FILLER_43_514 ();
 FILLCELL_X2 FILLER_43_523 ();
 FILLCELL_X16 FILLER_43_532 ();
 FILLCELL_X2 FILLER_43_548 ();
 FILLCELL_X1 FILLER_43_550 ();
 FILLCELL_X32 FILLER_43_558 ();
 FILLCELL_X32 FILLER_43_590 ();
 FILLCELL_X16 FILLER_43_622 ();
 FILLCELL_X2 FILLER_43_638 ();
 FILLCELL_X1 FILLER_43_640 ();
 FILLCELL_X2 FILLER_43_703 ();
 FILLCELL_X1 FILLER_43_707 ();
 FILLCELL_X1 FILLER_43_711 ();
 FILLCELL_X2 FILLER_43_732 ();
 FILLCELL_X8 FILLER_43_770 ();
 FILLCELL_X1 FILLER_43_778 ();
 FILLCELL_X2 FILLER_43_796 ();
 FILLCELL_X1 FILLER_43_798 ();
 FILLCELL_X16 FILLER_43_806 ();
 FILLCELL_X8 FILLER_43_822 ();
 FILLCELL_X2 FILLER_43_830 ();
 FILLCELL_X2 FILLER_43_847 ();
 FILLCELL_X2 FILLER_43_914 ();
 FILLCELL_X1 FILLER_43_916 ();
 FILLCELL_X4 FILLER_43_936 ();
 FILLCELL_X2 FILLER_43_940 ();
 FILLCELL_X1 FILLER_43_942 ();
 FILLCELL_X4 FILLER_43_958 ();
 FILLCELL_X1 FILLER_43_962 ();
 FILLCELL_X2 FILLER_43_980 ();
 FILLCELL_X1 FILLER_43_982 ();
 FILLCELL_X1 FILLER_43_1036 ();
 FILLCELL_X2 FILLER_43_1079 ();
 FILLCELL_X1 FILLER_43_1081 ();
 FILLCELL_X4 FILLER_43_1089 ();
 FILLCELL_X4 FILLER_43_1100 ();
 FILLCELL_X1 FILLER_43_1104 ();
 FILLCELL_X4 FILLER_43_1109 ();
 FILLCELL_X1 FILLER_43_1113 ();
 FILLCELL_X1 FILLER_43_1121 ();
 FILLCELL_X1 FILLER_43_1129 ();
 FILLCELL_X2 FILLER_43_1137 ();
 FILLCELL_X2 FILLER_43_1156 ();
 FILLCELL_X2 FILLER_43_1175 ();
 FILLCELL_X1 FILLER_43_1177 ();
 FILLCELL_X1 FILLER_43_1185 ();
 FILLCELL_X2 FILLER_43_1193 ();
 FILLCELL_X1 FILLER_43_1195 ();
 FILLCELL_X4 FILLER_43_1203 ();
 FILLCELL_X2 FILLER_43_1207 ();
 FILLCELL_X4 FILLER_43_1223 ();
 FILLCELL_X16 FILLER_44_1 ();
 FILLCELL_X8 FILLER_44_17 ();
 FILLCELL_X4 FILLER_44_62 ();
 FILLCELL_X8 FILLER_44_90 ();
 FILLCELL_X4 FILLER_44_98 ();
 FILLCELL_X1 FILLER_44_102 ();
 FILLCELL_X4 FILLER_44_124 ();
 FILLCELL_X2 FILLER_44_128 ();
 FILLCELL_X1 FILLER_44_130 ();
 FILLCELL_X8 FILLER_44_145 ();
 FILLCELL_X1 FILLER_44_153 ();
 FILLCELL_X2 FILLER_44_178 ();
 FILLCELL_X1 FILLER_44_180 ();
 FILLCELL_X16 FILLER_44_212 ();
 FILLCELL_X4 FILLER_44_228 ();
 FILLCELL_X2 FILLER_44_232 ();
 FILLCELL_X8 FILLER_44_272 ();
 FILLCELL_X1 FILLER_44_290 ();
 FILLCELL_X8 FILLER_44_305 ();
 FILLCELL_X2 FILLER_44_313 ();
 FILLCELL_X16 FILLER_44_319 ();
 FILLCELL_X1 FILLER_44_335 ();
 FILLCELL_X32 FILLER_44_350 ();
 FILLCELL_X16 FILLER_44_382 ();
 FILLCELL_X8 FILLER_44_398 ();
 FILLCELL_X4 FILLER_44_406 ();
 FILLCELL_X2 FILLER_44_410 ();
 FILLCELL_X32 FILLER_44_415 ();
 FILLCELL_X2 FILLER_44_455 ();
 FILLCELL_X1 FILLER_44_457 ();
 FILLCELL_X16 FILLER_44_465 ();
 FILLCELL_X8 FILLER_44_481 ();
 FILLCELL_X4 FILLER_44_489 ();
 FILLCELL_X16 FILLER_44_500 ();
 FILLCELL_X8 FILLER_44_516 ();
 FILLCELL_X2 FILLER_44_524 ();
 FILLCELL_X1 FILLER_44_526 ();
 FILLCELL_X32 FILLER_44_551 ();
 FILLCELL_X32 FILLER_44_583 ();
 FILLCELL_X16 FILLER_44_615 ();
 FILLCELL_X8 FILLER_44_632 ();
 FILLCELL_X2 FILLER_44_640 ();
 FILLCELL_X4 FILLER_44_649 ();
 FILLCELL_X1 FILLER_44_653 ();
 FILLCELL_X2 FILLER_44_721 ();
 FILLCELL_X4 FILLER_44_733 ();
 FILLCELL_X2 FILLER_44_747 ();
 FILLCELL_X2 FILLER_44_767 ();
 FILLCELL_X4 FILLER_44_779 ();
 FILLCELL_X1 FILLER_44_807 ();
 FILLCELL_X4 FILLER_44_822 ();
 FILLCELL_X8 FILLER_44_847 ();
 FILLCELL_X2 FILLER_44_855 ();
 FILLCELL_X1 FILLER_44_857 ();
 FILLCELL_X1 FILLER_44_865 ();
 FILLCELL_X1 FILLER_44_891 ();
 FILLCELL_X1 FILLER_44_909 ();
 FILLCELL_X4 FILLER_44_916 ();
 FILLCELL_X8 FILLER_44_923 ();
 FILLCELL_X4 FILLER_44_931 ();
 FILLCELL_X2 FILLER_44_969 ();
 FILLCELL_X1 FILLER_44_971 ();
 FILLCELL_X4 FILLER_44_998 ();
 FILLCELL_X1 FILLER_44_1002 ();
 FILLCELL_X4 FILLER_44_1016 ();
 FILLCELL_X4 FILLER_44_1034 ();
 FILLCELL_X2 FILLER_44_1038 ();
 FILLCELL_X1 FILLER_44_1040 ();
 FILLCELL_X2 FILLER_44_1054 ();
 FILLCELL_X1 FILLER_44_1063 ();
 FILLCELL_X2 FILLER_44_1071 ();
 FILLCELL_X8 FILLER_44_1080 ();
 FILLCELL_X4 FILLER_44_1088 ();
 FILLCELL_X2 FILLER_44_1092 ();
 FILLCELL_X1 FILLER_44_1094 ();
 FILLCELL_X2 FILLER_44_1102 ();
 FILLCELL_X1 FILLER_44_1104 ();
 FILLCELL_X1 FILLER_44_1125 ();
 FILLCELL_X16 FILLER_44_1157 ();
 FILLCELL_X1 FILLER_44_1190 ();
 FILLCELL_X2 FILLER_44_1208 ();
 FILLCELL_X1 FILLER_44_1227 ();
 FILLCELL_X2 FILLER_44_1235 ();
 FILLCELL_X4 FILLER_45_1 ();
 FILLCELL_X2 FILLER_45_30 ();
 FILLCELL_X1 FILLER_45_51 ();
 FILLCELL_X4 FILLER_45_59 ();
 FILLCELL_X2 FILLER_45_63 ();
 FILLCELL_X1 FILLER_45_65 ();
 FILLCELL_X8 FILLER_45_73 ();
 FILLCELL_X1 FILLER_45_81 ();
 FILLCELL_X32 FILLER_45_89 ();
 FILLCELL_X16 FILLER_45_121 ();
 FILLCELL_X4 FILLER_45_137 ();
 FILLCELL_X2 FILLER_45_141 ();
 FILLCELL_X8 FILLER_45_151 ();
 FILLCELL_X4 FILLER_45_159 ();
 FILLCELL_X2 FILLER_45_163 ();
 FILLCELL_X8 FILLER_45_182 ();
 FILLCELL_X1 FILLER_45_190 ();
 FILLCELL_X8 FILLER_45_203 ();
 FILLCELL_X4 FILLER_45_211 ();
 FILLCELL_X2 FILLER_45_215 ();
 FILLCELL_X4 FILLER_45_234 ();
 FILLCELL_X2 FILLER_45_238 ();
 FILLCELL_X1 FILLER_45_240 ();
 FILLCELL_X16 FILLER_45_265 ();
 FILLCELL_X4 FILLER_45_281 ();
 FILLCELL_X1 FILLER_45_285 ();
 FILLCELL_X16 FILLER_45_303 ();
 FILLCELL_X8 FILLER_45_319 ();
 FILLCELL_X4 FILLER_45_327 ();
 FILLCELL_X2 FILLER_45_331 ();
 FILLCELL_X32 FILLER_45_350 ();
 FILLCELL_X32 FILLER_45_382 ();
 FILLCELL_X16 FILLER_45_421 ();
 FILLCELL_X2 FILLER_45_437 ();
 FILLCELL_X1 FILLER_45_439 ();
 FILLCELL_X8 FILLER_45_468 ();
 FILLCELL_X1 FILLER_45_476 ();
 FILLCELL_X16 FILLER_45_484 ();
 FILLCELL_X4 FILLER_45_500 ();
 FILLCELL_X4 FILLER_45_528 ();
 FILLCELL_X1 FILLER_45_532 ();
 FILLCELL_X16 FILLER_45_557 ();
 FILLCELL_X1 FILLER_45_573 ();
 FILLCELL_X32 FILLER_45_581 ();
 FILLCELL_X16 FILLER_45_613 ();
 FILLCELL_X2 FILLER_45_629 ();
 FILLCELL_X1 FILLER_45_631 ();
 FILLCELL_X2 FILLER_45_656 ();
 FILLCELL_X1 FILLER_45_658 ();
 FILLCELL_X2 FILLER_45_666 ();
 FILLCELL_X1 FILLER_45_668 ();
 FILLCELL_X4 FILLER_45_676 ();
 FILLCELL_X1 FILLER_45_680 ();
 FILLCELL_X4 FILLER_45_698 ();
 FILLCELL_X1 FILLER_45_702 ();
 FILLCELL_X2 FILLER_45_706 ();
 FILLCELL_X4 FILLER_45_715 ();
 FILLCELL_X2 FILLER_45_719 ();
 FILLCELL_X8 FILLER_45_767 ();
 FILLCELL_X1 FILLER_45_844 ();
 FILLCELL_X8 FILLER_45_852 ();
 FILLCELL_X4 FILLER_45_860 ();
 FILLCELL_X2 FILLER_45_864 ();
 FILLCELL_X8 FILLER_45_888 ();
 FILLCELL_X4 FILLER_45_917 ();
 FILLCELL_X2 FILLER_45_952 ();
 FILLCELL_X1 FILLER_45_954 ();
 FILLCELL_X4 FILLER_45_962 ();
 FILLCELL_X2 FILLER_45_966 ();
 FILLCELL_X1 FILLER_45_968 ();
 FILLCELL_X1 FILLER_45_976 ();
 FILLCELL_X1 FILLER_45_990 ();
 FILLCELL_X8 FILLER_45_1008 ();
 FILLCELL_X8 FILLER_45_1033 ();
 FILLCELL_X4 FILLER_45_1041 ();
 FILLCELL_X2 FILLER_45_1045 ();
 FILLCELL_X1 FILLER_45_1054 ();
 FILLCELL_X4 FILLER_45_1062 ();
 FILLCELL_X1 FILLER_45_1073 ();
 FILLCELL_X1 FILLER_45_1091 ();
 FILLCELL_X4 FILLER_45_1112 ();
 FILLCELL_X2 FILLER_45_1116 ();
 FILLCELL_X2 FILLER_45_1135 ();
 FILLCELL_X16 FILLER_45_1150 ();
 FILLCELL_X8 FILLER_45_1166 ();
 FILLCELL_X1 FILLER_45_1174 ();
 FILLCELL_X8 FILLER_45_1199 ();
 FILLCELL_X2 FILLER_45_1207 ();
 FILLCELL_X1 FILLER_45_1209 ();
 FILLCELL_X4 FILLER_46_4 ();
 FILLCELL_X8 FILLER_46_11 ();
 FILLCELL_X32 FILLER_46_52 ();
 FILLCELL_X1 FILLER_46_84 ();
 FILLCELL_X2 FILLER_46_135 ();
 FILLCELL_X1 FILLER_46_137 ();
 FILLCELL_X8 FILLER_46_162 ();
 FILLCELL_X4 FILLER_46_170 ();
 FILLCELL_X1 FILLER_46_174 ();
 FILLCELL_X16 FILLER_46_199 ();
 FILLCELL_X4 FILLER_46_215 ();
 FILLCELL_X1 FILLER_46_219 ();
 FILLCELL_X2 FILLER_46_227 ();
 FILLCELL_X1 FILLER_46_229 ();
 FILLCELL_X2 FILLER_46_254 ();
 FILLCELL_X16 FILLER_46_263 ();
 FILLCELL_X2 FILLER_46_279 ();
 FILLCELL_X1 FILLER_46_281 ();
 FILLCELL_X8 FILLER_46_289 ();
 FILLCELL_X8 FILLER_46_304 ();
 FILLCELL_X1 FILLER_46_312 ();
 FILLCELL_X8 FILLER_46_330 ();
 FILLCELL_X4 FILLER_46_338 ();
 FILLCELL_X8 FILLER_46_349 ();
 FILLCELL_X1 FILLER_46_357 ();
 FILLCELL_X8 FILLER_46_389 ();
 FILLCELL_X1 FILLER_46_402 ();
 FILLCELL_X8 FILLER_46_427 ();
 FILLCELL_X4 FILLER_46_435 ();
 FILLCELL_X2 FILLER_46_439 ();
 FILLCELL_X1 FILLER_46_441 ();
 FILLCELL_X2 FILLER_46_466 ();
 FILLCELL_X4 FILLER_46_475 ();
 FILLCELL_X8 FILLER_46_499 ();
 FILLCELL_X4 FILLER_46_507 ();
 FILLCELL_X1 FILLER_46_511 ();
 FILLCELL_X32 FILLER_46_558 ();
 FILLCELL_X32 FILLER_46_590 ();
 FILLCELL_X8 FILLER_46_622 ();
 FILLCELL_X1 FILLER_46_630 ();
 FILLCELL_X8 FILLER_46_632 ();
 FILLCELL_X4 FILLER_46_640 ();
 FILLCELL_X2 FILLER_46_644 ();
 FILLCELL_X32 FILLER_46_663 ();
 FILLCELL_X4 FILLER_46_695 ();
 FILLCELL_X2 FILLER_46_699 ();
 FILLCELL_X16 FILLER_46_724 ();
 FILLCELL_X1 FILLER_46_740 ();
 FILLCELL_X4 FILLER_46_773 ();
 FILLCELL_X4 FILLER_46_784 ();
 FILLCELL_X2 FILLER_46_788 ();
 FILLCELL_X1 FILLER_46_790 ();
 FILLCELL_X1 FILLER_46_800 ();
 FILLCELL_X16 FILLER_46_821 ();
 FILLCELL_X4 FILLER_46_837 ();
 FILLCELL_X2 FILLER_46_841 ();
 FILLCELL_X1 FILLER_46_843 ();
 FILLCELL_X4 FILLER_46_868 ();
 FILLCELL_X1 FILLER_46_872 ();
 FILLCELL_X2 FILLER_46_876 ();
 FILLCELL_X1 FILLER_46_878 ();
 FILLCELL_X16 FILLER_46_886 ();
 FILLCELL_X4 FILLER_46_902 ();
 FILLCELL_X2 FILLER_46_906 ();
 FILLCELL_X16 FILLER_46_914 ();
 FILLCELL_X4 FILLER_46_930 ();
 FILLCELL_X1 FILLER_46_934 ();
 FILLCELL_X32 FILLER_46_938 ();
 FILLCELL_X16 FILLER_46_970 ();
 FILLCELL_X2 FILLER_46_986 ();
 FILLCELL_X1 FILLER_46_1005 ();
 FILLCELL_X16 FILLER_46_1019 ();
 FILLCELL_X8 FILLER_46_1035 ();
 FILLCELL_X8 FILLER_46_1090 ();
 FILLCELL_X1 FILLER_46_1098 ();
 FILLCELL_X8 FILLER_46_1123 ();
 FILLCELL_X2 FILLER_46_1131 ();
 FILLCELL_X1 FILLER_46_1133 ();
 FILLCELL_X4 FILLER_46_1151 ();
 FILLCELL_X1 FILLER_46_1155 ();
 FILLCELL_X16 FILLER_46_1161 ();
 FILLCELL_X4 FILLER_46_1177 ();
 FILLCELL_X2 FILLER_46_1181 ();
 FILLCELL_X1 FILLER_46_1183 ();
 FILLCELL_X16 FILLER_46_1193 ();
 FILLCELL_X4 FILLER_46_1209 ();
 FILLCELL_X1 FILLER_46_1213 ();
 FILLCELL_X4 FILLER_46_1236 ();
 FILLCELL_X1 FILLER_47_1 ();
 FILLCELL_X16 FILLER_47_5 ();
 FILLCELL_X8 FILLER_47_21 ();
 FILLCELL_X4 FILLER_47_29 ();
 FILLCELL_X2 FILLER_47_33 ();
 FILLCELL_X1 FILLER_47_35 ();
 FILLCELL_X4 FILLER_47_53 ();
 FILLCELL_X1 FILLER_47_57 ();
 FILLCELL_X16 FILLER_47_75 ();
 FILLCELL_X2 FILLER_47_91 ();
 FILLCELL_X1 FILLER_47_93 ();
 FILLCELL_X2 FILLER_47_111 ();
 FILLCELL_X1 FILLER_47_113 ();
 FILLCELL_X1 FILLER_47_121 ();
 FILLCELL_X16 FILLER_47_139 ();
 FILLCELL_X4 FILLER_47_155 ();
 FILLCELL_X1 FILLER_47_159 ();
 FILLCELL_X2 FILLER_47_167 ();
 FILLCELL_X4 FILLER_47_176 ();
 FILLCELL_X8 FILLER_47_194 ();
 FILLCELL_X2 FILLER_47_202 ();
 FILLCELL_X4 FILLER_47_221 ();
 FILLCELL_X2 FILLER_47_225 ();
 FILLCELL_X1 FILLER_47_227 ();
 FILLCELL_X4 FILLER_47_235 ();
 FILLCELL_X8 FILLER_47_247 ();
 FILLCELL_X4 FILLER_47_255 ();
 FILLCELL_X1 FILLER_47_259 ();
 FILLCELL_X2 FILLER_47_269 ();
 FILLCELL_X1 FILLER_47_271 ();
 FILLCELL_X8 FILLER_47_296 ();
 FILLCELL_X2 FILLER_47_304 ();
 FILLCELL_X1 FILLER_47_306 ();
 FILLCELL_X2 FILLER_47_314 ();
 FILLCELL_X4 FILLER_47_335 ();
 FILLCELL_X1 FILLER_47_339 ();
 FILLCELL_X2 FILLER_47_354 ();
 FILLCELL_X1 FILLER_47_356 ();
 FILLCELL_X1 FILLER_47_381 ();
 FILLCELL_X4 FILLER_47_399 ();
 FILLCELL_X2 FILLER_47_427 ();
 FILLCELL_X1 FILLER_47_429 ();
 FILLCELL_X4 FILLER_47_437 ();
 FILLCELL_X1 FILLER_47_441 ();
 FILLCELL_X4 FILLER_47_449 ();
 FILLCELL_X1 FILLER_47_453 ();
 FILLCELL_X4 FILLER_47_461 ();
 FILLCELL_X2 FILLER_47_465 ();
 FILLCELL_X1 FILLER_47_467 ();
 FILLCELL_X2 FILLER_47_492 ();
 FILLCELL_X1 FILLER_47_494 ();
 FILLCELL_X8 FILLER_47_505 ();
 FILLCELL_X1 FILLER_47_513 ();
 FILLCELL_X1 FILLER_47_518 ();
 FILLCELL_X32 FILLER_47_549 ();
 FILLCELL_X32 FILLER_47_581 ();
 FILLCELL_X32 FILLER_47_613 ();
 FILLCELL_X32 FILLER_47_645 ();
 FILLCELL_X32 FILLER_47_677 ();
 FILLCELL_X8 FILLER_47_709 ();
 FILLCELL_X16 FILLER_47_724 ();
 FILLCELL_X8 FILLER_47_740 ();
 FILLCELL_X4 FILLER_47_748 ();
 FILLCELL_X16 FILLER_47_762 ();
 FILLCELL_X2 FILLER_47_781 ();
 FILLCELL_X1 FILLER_47_783 ();
 FILLCELL_X2 FILLER_47_787 ();
 FILLCELL_X1 FILLER_47_789 ();
 FILLCELL_X4 FILLER_47_793 ();
 FILLCELL_X32 FILLER_47_802 ();
 FILLCELL_X8 FILLER_47_834 ();
 FILLCELL_X1 FILLER_47_866 ();
 FILLCELL_X16 FILLER_47_895 ();
 FILLCELL_X8 FILLER_47_911 ();
 FILLCELL_X4 FILLER_47_919 ();
 FILLCELL_X1 FILLER_47_923 ();
 FILLCELL_X4 FILLER_47_948 ();
 FILLCELL_X8 FILLER_47_959 ();
 FILLCELL_X2 FILLER_47_967 ();
 FILLCELL_X2 FILLER_47_976 ();
 FILLCELL_X1 FILLER_47_978 ();
 FILLCELL_X1 FILLER_47_1004 ();
 FILLCELL_X32 FILLER_47_1012 ();
 FILLCELL_X32 FILLER_47_1044 ();
 FILLCELL_X32 FILLER_47_1076 ();
 FILLCELL_X16 FILLER_47_1108 ();
 FILLCELL_X4 FILLER_47_1124 ();
 FILLCELL_X2 FILLER_47_1128 ();
 FILLCELL_X1 FILLER_47_1130 ();
 FILLCELL_X2 FILLER_47_1155 ();
 FILLCELL_X1 FILLER_47_1157 ();
 FILLCELL_X16 FILLER_47_1175 ();
 FILLCELL_X4 FILLER_47_1191 ();
 FILLCELL_X1 FILLER_47_1195 ();
 FILLCELL_X16 FILLER_47_1199 ();
 FILLCELL_X1 FILLER_47_1215 ();
 FILLCELL_X8 FILLER_47_1225 ();
 FILLCELL_X4 FILLER_47_1233 ();
 FILLCELL_X4 FILLER_48_1 ();
 FILLCELL_X2 FILLER_48_5 ();
 FILLCELL_X8 FILLER_48_24 ();
 FILLCELL_X4 FILLER_48_32 ();
 FILLCELL_X2 FILLER_48_36 ();
 FILLCELL_X2 FILLER_48_55 ();
 FILLCELL_X1 FILLER_48_57 ();
 FILLCELL_X2 FILLER_48_65 ();
 FILLCELL_X2 FILLER_48_91 ();
 FILLCELL_X2 FILLER_48_107 ();
 FILLCELL_X8 FILLER_48_116 ();
 FILLCELL_X2 FILLER_48_124 ();
 FILLCELL_X1 FILLER_48_126 ();
 FILLCELL_X16 FILLER_48_134 ();
 FILLCELL_X2 FILLER_48_150 ();
 FILLCELL_X16 FILLER_48_169 ();
 FILLCELL_X1 FILLER_48_185 ();
 FILLCELL_X8 FILLER_48_193 ();
 FILLCELL_X2 FILLER_48_201 ();
 FILLCELL_X1 FILLER_48_203 ();
 FILLCELL_X4 FILLER_48_225 ();
 FILLCELL_X1 FILLER_48_229 ();
 FILLCELL_X4 FILLER_48_247 ();
 FILLCELL_X2 FILLER_48_251 ();
 FILLCELL_X8 FILLER_48_270 ();
 FILLCELL_X2 FILLER_48_285 ();
 FILLCELL_X1 FILLER_48_287 ();
 FILLCELL_X4 FILLER_48_305 ();
 FILLCELL_X4 FILLER_48_326 ();
 FILLCELL_X1 FILLER_48_330 ();
 FILLCELL_X2 FILLER_48_348 ();
 FILLCELL_X1 FILLER_48_350 ();
 FILLCELL_X16 FILLER_48_382 ();
 FILLCELL_X2 FILLER_48_398 ();
 FILLCELL_X1 FILLER_48_400 ();
 FILLCELL_X2 FILLER_48_432 ();
 FILLCELL_X1 FILLER_48_434 ();
 FILLCELL_X2 FILLER_48_452 ();
 FILLCELL_X2 FILLER_48_461 ();
 FILLCELL_X2 FILLER_48_466 ();
 FILLCELL_X1 FILLER_48_468 ();
 FILLCELL_X8 FILLER_48_472 ();
 FILLCELL_X4 FILLER_48_480 ();
 FILLCELL_X1 FILLER_48_484 ();
 FILLCELL_X8 FILLER_48_503 ();
 FILLCELL_X1 FILLER_48_511 ();
 FILLCELL_X8 FILLER_48_516 ();
 FILLCELL_X32 FILLER_48_561 ();
 FILLCELL_X32 FILLER_48_593 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X4 FILLER_48_632 ();
 FILLCELL_X2 FILLER_48_636 ();
 FILLCELL_X1 FILLER_48_638 ();
 FILLCELL_X4 FILLER_48_656 ();
 FILLCELL_X1 FILLER_48_660 ();
 FILLCELL_X16 FILLER_48_678 ();
 FILLCELL_X8 FILLER_48_694 ();
 FILLCELL_X4 FILLER_48_702 ();
 FILLCELL_X1 FILLER_48_706 ();
 FILLCELL_X32 FILLER_48_724 ();
 FILLCELL_X8 FILLER_48_756 ();
 FILLCELL_X4 FILLER_48_764 ();
 FILLCELL_X1 FILLER_48_768 ();
 FILLCELL_X16 FILLER_48_789 ();
 FILLCELL_X4 FILLER_48_805 ();
 FILLCELL_X2 FILLER_48_809 ();
 FILLCELL_X1 FILLER_48_811 ();
 FILLCELL_X4 FILLER_48_815 ();
 FILLCELL_X4 FILLER_48_822 ();
 FILLCELL_X4 FILLER_48_829 ();
 FILLCELL_X2 FILLER_48_833 ();
 FILLCELL_X1 FILLER_48_835 ();
 FILLCELL_X1 FILLER_48_839 ();
 FILLCELL_X4 FILLER_48_860 ();
 FILLCELL_X2 FILLER_48_868 ();
 FILLCELL_X1 FILLER_48_870 ();
 FILLCELL_X8 FILLER_48_905 ();
 FILLCELL_X2 FILLER_48_916 ();
 FILLCELL_X2 FILLER_48_1056 ();
 FILLCELL_X8 FILLER_48_1075 ();
 FILLCELL_X1 FILLER_48_1083 ();
 FILLCELL_X4 FILLER_48_1118 ();
 FILLCELL_X1 FILLER_48_1122 ();
 FILLCELL_X16 FILLER_48_1176 ();
 FILLCELL_X4 FILLER_48_1192 ();
 FILLCELL_X2 FILLER_48_1196 ();
 FILLCELL_X8 FILLER_48_1201 ();
 FILLCELL_X2 FILLER_48_1209 ();
 FILLCELL_X1 FILLER_48_1211 ();
 FILLCELL_X4 FILLER_48_1215 ();
 FILLCELL_X2 FILLER_48_1219 ();
 FILLCELL_X8 FILLER_48_1228 ();
 FILLCELL_X4 FILLER_48_1236 ();
 FILLCELL_X2 FILLER_49_16 ();
 FILLCELL_X1 FILLER_49_18 ();
 FILLCELL_X4 FILLER_49_45 ();
 FILLCELL_X1 FILLER_49_49 ();
 FILLCELL_X8 FILLER_49_64 ();
 FILLCELL_X1 FILLER_49_72 ();
 FILLCELL_X16 FILLER_49_80 ();
 FILLCELL_X8 FILLER_49_96 ();
 FILLCELL_X4 FILLER_49_104 ();
 FILLCELL_X2 FILLER_49_108 ();
 FILLCELL_X1 FILLER_49_110 ();
 FILLCELL_X4 FILLER_49_135 ();
 FILLCELL_X1 FILLER_49_144 ();
 FILLCELL_X16 FILLER_49_162 ();
 FILLCELL_X8 FILLER_49_178 ();
 FILLCELL_X1 FILLER_49_186 ();
 FILLCELL_X2 FILLER_49_194 ();
 FILLCELL_X1 FILLER_49_196 ();
 FILLCELL_X8 FILLER_49_203 ();
 FILLCELL_X4 FILLER_49_211 ();
 FILLCELL_X16 FILLER_49_222 ();
 FILLCELL_X8 FILLER_49_238 ();
 FILLCELL_X2 FILLER_49_246 ();
 FILLCELL_X16 FILLER_49_272 ();
 FILLCELL_X8 FILLER_49_288 ();
 FILLCELL_X2 FILLER_49_310 ();
 FILLCELL_X4 FILLER_49_319 ();
 FILLCELL_X2 FILLER_49_323 ();
 FILLCELL_X8 FILLER_49_342 ();
 FILLCELL_X4 FILLER_49_350 ();
 FILLCELL_X1 FILLER_49_354 ();
 FILLCELL_X16 FILLER_49_376 ();
 FILLCELL_X8 FILLER_49_392 ();
 FILLCELL_X4 FILLER_49_400 ();
 FILLCELL_X1 FILLER_49_404 ();
 FILLCELL_X4 FILLER_49_408 ();
 FILLCELL_X1 FILLER_49_412 ();
 FILLCELL_X2 FILLER_49_430 ();
 FILLCELL_X1 FILLER_49_449 ();
 FILLCELL_X2 FILLER_49_475 ();
 FILLCELL_X8 FILLER_49_484 ();
 FILLCELL_X4 FILLER_49_492 ();
 FILLCELL_X2 FILLER_49_496 ();
 FILLCELL_X1 FILLER_49_498 ();
 FILLCELL_X16 FILLER_49_506 ();
 FILLCELL_X8 FILLER_49_522 ();
 FILLCELL_X2 FILLER_49_530 ();
 FILLCELL_X2 FILLER_49_553 ();
 FILLCELL_X1 FILLER_49_555 ();
 FILLCELL_X2 FILLER_49_560 ();
 FILLCELL_X1 FILLER_49_562 ();
 FILLCELL_X32 FILLER_49_587 ();
 FILLCELL_X16 FILLER_49_619 ();
 FILLCELL_X2 FILLER_49_642 ();
 FILLCELL_X1 FILLER_49_644 ();
 FILLCELL_X4 FILLER_49_652 ();
 FILLCELL_X2 FILLER_49_656 ();
 FILLCELL_X4 FILLER_49_665 ();
 FILLCELL_X2 FILLER_49_669 ();
 FILLCELL_X4 FILLER_49_688 ();
 FILLCELL_X1 FILLER_49_692 ();
 FILLCELL_X4 FILLER_49_700 ();
 FILLCELL_X1 FILLER_49_704 ();
 FILLCELL_X8 FILLER_49_712 ();
 FILLCELL_X2 FILLER_49_720 ();
 FILLCELL_X1 FILLER_49_722 ();
 FILLCELL_X4 FILLER_49_730 ();
 FILLCELL_X1 FILLER_49_734 ();
 FILLCELL_X4 FILLER_49_759 ();
 FILLCELL_X8 FILLER_49_793 ();
 FILLCELL_X1 FILLER_49_801 ();
 FILLCELL_X1 FILLER_49_822 ();
 FILLCELL_X2 FILLER_49_830 ();
 FILLCELL_X1 FILLER_49_835 ();
 FILLCELL_X4 FILLER_49_839 ();
 FILLCELL_X2 FILLER_49_843 ();
 FILLCELL_X1 FILLER_49_845 ();
 FILLCELL_X2 FILLER_49_849 ();
 FILLCELL_X1 FILLER_49_851 ();
 FILLCELL_X8 FILLER_49_855 ();
 FILLCELL_X4 FILLER_49_863 ();
 FILLCELL_X4 FILLER_49_874 ();
 FILLCELL_X2 FILLER_49_878 ();
 FILLCELL_X4 FILLER_49_883 ();
 FILLCELL_X1 FILLER_49_924 ();
 FILLCELL_X1 FILLER_49_942 ();
 FILLCELL_X2 FILLER_49_950 ();
 FILLCELL_X1 FILLER_49_952 ();
 FILLCELL_X2 FILLER_49_1012 ();
 FILLCELL_X1 FILLER_49_1014 ();
 FILLCELL_X4 FILLER_49_1032 ();
 FILLCELL_X2 FILLER_49_1036 ();
 FILLCELL_X1 FILLER_49_1038 ();
 FILLCELL_X2 FILLER_49_1107 ();
 FILLCELL_X8 FILLER_49_1116 ();
 FILLCELL_X4 FILLER_49_1124 ();
 FILLCELL_X2 FILLER_49_1128 ();
 FILLCELL_X1 FILLER_49_1170 ();
 FILLCELL_X8 FILLER_49_1188 ();
 FILLCELL_X4 FILLER_49_1196 ();
 FILLCELL_X2 FILLER_49_1200 ();
 FILLCELL_X1 FILLER_49_1236 ();
 FILLCELL_X2 FILLER_50_1 ();
 FILLCELL_X1 FILLER_50_3 ();
 FILLCELL_X2 FILLER_50_14 ();
 FILLCELL_X1 FILLER_50_16 ();
 FILLCELL_X16 FILLER_50_21 ();
 FILLCELL_X4 FILLER_50_37 ();
 FILLCELL_X1 FILLER_50_41 ();
 FILLCELL_X4 FILLER_50_66 ();
 FILLCELL_X2 FILLER_50_70 ();
 FILLCELL_X4 FILLER_50_86 ();
 FILLCELL_X2 FILLER_50_90 ();
 FILLCELL_X2 FILLER_50_127 ();
 FILLCELL_X1 FILLER_50_129 ();
 FILLCELL_X4 FILLER_50_137 ();
 FILLCELL_X2 FILLER_50_141 ();
 FILLCELL_X4 FILLER_50_150 ();
 FILLCELL_X2 FILLER_50_154 ();
 FILLCELL_X4 FILLER_50_163 ();
 FILLCELL_X2 FILLER_50_174 ();
 FILLCELL_X8 FILLER_50_207 ();
 FILLCELL_X2 FILLER_50_215 ();
 FILLCELL_X4 FILLER_50_237 ();
 FILLCELL_X2 FILLER_50_241 ();
 FILLCELL_X2 FILLER_50_250 ();
 FILLCELL_X32 FILLER_50_266 ();
 FILLCELL_X8 FILLER_50_298 ();
 FILLCELL_X2 FILLER_50_306 ();
 FILLCELL_X1 FILLER_50_308 ();
 FILLCELL_X4 FILLER_50_312 ();
 FILLCELL_X2 FILLER_50_316 ();
 FILLCELL_X1 FILLER_50_318 ();
 FILLCELL_X2 FILLER_50_329 ();
 FILLCELL_X1 FILLER_50_331 ();
 FILLCELL_X4 FILLER_50_349 ();
 FILLCELL_X2 FILLER_50_353 ();
 FILLCELL_X16 FILLER_50_368 ();
 FILLCELL_X4 FILLER_50_384 ();
 FILLCELL_X2 FILLER_50_388 ();
 FILLCELL_X1 FILLER_50_390 ();
 FILLCELL_X16 FILLER_50_398 ();
 FILLCELL_X2 FILLER_50_414 ();
 FILLCELL_X8 FILLER_50_421 ();
 FILLCELL_X2 FILLER_50_429 ();
 FILLCELL_X4 FILLER_50_436 ();
 FILLCELL_X1 FILLER_50_440 ();
 FILLCELL_X8 FILLER_50_455 ();
 FILLCELL_X1 FILLER_50_477 ();
 FILLCELL_X1 FILLER_50_495 ();
 FILLCELL_X16 FILLER_50_516 ();
 FILLCELL_X8 FILLER_50_532 ();
 FILLCELL_X2 FILLER_50_540 ();
 FILLCELL_X32 FILLER_50_559 ();
 FILLCELL_X32 FILLER_50_591 ();
 FILLCELL_X8 FILLER_50_623 ();
 FILLCELL_X8 FILLER_50_632 ();
 FILLCELL_X1 FILLER_50_640 ();
 FILLCELL_X8 FILLER_50_679 ();
 FILLCELL_X2 FILLER_50_687 ();
 FILLCELL_X4 FILLER_50_713 ();
 FILLCELL_X2 FILLER_50_717 ();
 FILLCELL_X1 FILLER_50_719 ();
 FILLCELL_X8 FILLER_50_744 ();
 FILLCELL_X4 FILLER_50_752 ();
 FILLCELL_X2 FILLER_50_756 ();
 FILLCELL_X1 FILLER_50_758 ();
 FILLCELL_X16 FILLER_50_786 ();
 FILLCELL_X1 FILLER_50_802 ();
 FILLCELL_X2 FILLER_50_820 ();
 FILLCELL_X1 FILLER_50_857 ();
 FILLCELL_X4 FILLER_50_874 ();
 FILLCELL_X4 FILLER_50_929 ();
 FILLCELL_X1 FILLER_50_933 ();
 FILLCELL_X8 FILLER_50_948 ();
 FILLCELL_X2 FILLER_50_1033 ();
 FILLCELL_X4 FILLER_50_1078 ();
 FILLCELL_X16 FILLER_50_1101 ();
 FILLCELL_X1 FILLER_50_1117 ();
 FILLCELL_X16 FILLER_50_1149 ();
 FILLCELL_X2 FILLER_50_1165 ();
 FILLCELL_X8 FILLER_50_1172 ();
 FILLCELL_X2 FILLER_50_1180 ();
 FILLCELL_X4 FILLER_50_1202 ();
 FILLCELL_X4 FILLER_51_32 ();
 FILLCELL_X2 FILLER_51_36 ();
 FILLCELL_X1 FILLER_51_38 ();
 FILLCELL_X2 FILLER_51_46 ();
 FILLCELL_X4 FILLER_51_51 ();
 FILLCELL_X2 FILLER_51_55 ();
 FILLCELL_X4 FILLER_51_81 ();
 FILLCELL_X2 FILLER_51_85 ();
 FILLCELL_X1 FILLER_51_104 ();
 FILLCELL_X4 FILLER_51_119 ();
 FILLCELL_X1 FILLER_51_123 ();
 FILLCELL_X1 FILLER_51_139 ();
 FILLCELL_X8 FILLER_51_147 ();
 FILLCELL_X8 FILLER_51_172 ();
 FILLCELL_X4 FILLER_51_180 ();
 FILLCELL_X1 FILLER_51_184 ();
 FILLCELL_X16 FILLER_51_209 ();
 FILLCELL_X8 FILLER_51_225 ();
 FILLCELL_X4 FILLER_51_233 ();
 FILLCELL_X1 FILLER_51_237 ();
 FILLCELL_X16 FILLER_51_269 ();
 FILLCELL_X1 FILLER_51_285 ();
 FILLCELL_X16 FILLER_51_310 ();
 FILLCELL_X1 FILLER_51_340 ();
 FILLCELL_X16 FILLER_51_348 ();
 FILLCELL_X2 FILLER_51_364 ();
 FILLCELL_X1 FILLER_51_366 ();
 FILLCELL_X8 FILLER_51_384 ();
 FILLCELL_X1 FILLER_51_392 ();
 FILLCELL_X4 FILLER_51_407 ();
 FILLCELL_X1 FILLER_51_411 ();
 FILLCELL_X2 FILLER_51_429 ();
 FILLCELL_X1 FILLER_51_431 ();
 FILLCELL_X8 FILLER_51_456 ();
 FILLCELL_X4 FILLER_51_464 ();
 FILLCELL_X4 FILLER_51_472 ();
 FILLCELL_X2 FILLER_51_476 ();
 FILLCELL_X1 FILLER_51_478 ();
 FILLCELL_X1 FILLER_51_496 ();
 FILLCELL_X4 FILLER_51_509 ();
 FILLCELL_X1 FILLER_51_520 ();
 FILLCELL_X32 FILLER_51_528 ();
 FILLCELL_X32 FILLER_51_560 ();
 FILLCELL_X32 FILLER_51_592 ();
 FILLCELL_X32 FILLER_51_624 ();
 FILLCELL_X16 FILLER_51_656 ();
 FILLCELL_X8 FILLER_51_672 ();
 FILLCELL_X4 FILLER_51_680 ();
 FILLCELL_X1 FILLER_51_684 ();
 FILLCELL_X16 FILLER_51_692 ();
 FILLCELL_X8 FILLER_51_708 ();
 FILLCELL_X4 FILLER_51_716 ();
 FILLCELL_X1 FILLER_51_720 ();
 FILLCELL_X1 FILLER_51_738 ();
 FILLCELL_X4 FILLER_51_756 ();
 FILLCELL_X2 FILLER_51_760 ();
 FILLCELL_X1 FILLER_51_762 ();
 FILLCELL_X8 FILLER_51_781 ();
 FILLCELL_X4 FILLER_51_789 ();
 FILLCELL_X2 FILLER_51_793 ();
 FILLCELL_X1 FILLER_51_795 ();
 FILLCELL_X4 FILLER_51_799 ();
 FILLCELL_X2 FILLER_51_803 ();
 FILLCELL_X2 FILLER_51_812 ();
 FILLCELL_X2 FILLER_51_824 ();
 FILLCELL_X2 FILLER_51_829 ();
 FILLCELL_X2 FILLER_51_834 ();
 FILLCELL_X2 FILLER_51_843 ();
 FILLCELL_X8 FILLER_51_848 ();
 FILLCELL_X4 FILLER_51_873 ();
 FILLCELL_X2 FILLER_51_877 ();
 FILLCELL_X1 FILLER_51_879 ();
 FILLCELL_X1 FILLER_51_886 ();
 FILLCELL_X2 FILLER_51_900 ();
 FILLCELL_X1 FILLER_51_902 ();
 FILLCELL_X1 FILLER_51_919 ();
 FILLCELL_X2 FILLER_51_923 ();
 FILLCELL_X8 FILLER_51_932 ();
 FILLCELL_X32 FILLER_51_949 ();
 FILLCELL_X16 FILLER_51_981 ();
 FILLCELL_X8 FILLER_51_997 ();
 FILLCELL_X4 FILLER_51_1005 ();
 FILLCELL_X16 FILLER_51_1013 ();
 FILLCELL_X4 FILLER_51_1029 ();
 FILLCELL_X2 FILLER_51_1033 ();
 FILLCELL_X1 FILLER_51_1035 ();
 FILLCELL_X16 FILLER_51_1040 ();
 FILLCELL_X4 FILLER_51_1056 ();
 FILLCELL_X2 FILLER_51_1060 ();
 FILLCELL_X4 FILLER_51_1086 ();
 FILLCELL_X1 FILLER_51_1090 ();
 FILLCELL_X8 FILLER_51_1098 ();
 FILLCELL_X4 FILLER_51_1106 ();
 FILLCELL_X2 FILLER_51_1238 ();
 FILLCELL_X1 FILLER_52_4 ();
 FILLCELL_X2 FILLER_52_57 ();
 FILLCELL_X32 FILLER_52_83 ();
 FILLCELL_X8 FILLER_52_115 ();
 FILLCELL_X4 FILLER_52_123 ();
 FILLCELL_X2 FILLER_52_127 ();
 FILLCELL_X1 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_147 ();
 FILLCELL_X4 FILLER_52_179 ();
 FILLCELL_X1 FILLER_52_183 ();
 FILLCELL_X1 FILLER_52_194 ();
 FILLCELL_X8 FILLER_52_205 ();
 FILLCELL_X4 FILLER_52_230 ();
 FILLCELL_X2 FILLER_52_234 ();
 FILLCELL_X2 FILLER_52_267 ();
 FILLCELL_X8 FILLER_52_280 ();
 FILLCELL_X4 FILLER_52_288 ();
 FILLCELL_X4 FILLER_52_299 ();
 FILLCELL_X8 FILLER_52_320 ();
 FILLCELL_X4 FILLER_52_328 ();
 FILLCELL_X8 FILLER_52_349 ();
 FILLCELL_X4 FILLER_52_357 ();
 FILLCELL_X2 FILLER_52_361 ();
 FILLCELL_X1 FILLER_52_363 ();
 FILLCELL_X2 FILLER_52_371 ();
 FILLCELL_X2 FILLER_52_380 ();
 FILLCELL_X4 FILLER_52_399 ();
 FILLCELL_X2 FILLER_52_403 ();
 FILLCELL_X2 FILLER_52_422 ();
 FILLCELL_X1 FILLER_52_424 ();
 FILLCELL_X4 FILLER_52_432 ();
 FILLCELL_X2 FILLER_52_436 ();
 FILLCELL_X2 FILLER_52_462 ();
 FILLCELL_X4 FILLER_52_495 ();
 FILLCELL_X1 FILLER_52_499 ();
 FILLCELL_X1 FILLER_52_514 ();
 FILLCELL_X32 FILLER_52_532 ();
 FILLCELL_X32 FILLER_52_564 ();
 FILLCELL_X1 FILLER_52_596 ();
 FILLCELL_X16 FILLER_52_602 ();
 FILLCELL_X8 FILLER_52_618 ();
 FILLCELL_X4 FILLER_52_626 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X2 FILLER_52_632 ();
 FILLCELL_X1 FILLER_52_634 ();
 FILLCELL_X4 FILLER_52_652 ();
 FILLCELL_X2 FILLER_52_656 ();
 FILLCELL_X1 FILLER_52_665 ();
 FILLCELL_X2 FILLER_52_675 ();
 FILLCELL_X1 FILLER_52_677 ();
 FILLCELL_X2 FILLER_52_749 ();
 FILLCELL_X16 FILLER_52_761 ();
 FILLCELL_X2 FILLER_52_777 ();
 FILLCELL_X2 FILLER_52_813 ();
 FILLCELL_X1 FILLER_52_815 ();
 FILLCELL_X2 FILLER_52_819 ();
 FILLCELL_X16 FILLER_52_828 ();
 FILLCELL_X8 FILLER_52_844 ();
 FILLCELL_X4 FILLER_52_852 ();
 FILLCELL_X2 FILLER_52_856 ();
 FILLCELL_X1 FILLER_52_858 ();
 FILLCELL_X16 FILLER_52_862 ();
 FILLCELL_X4 FILLER_52_878 ();
 FILLCELL_X2 FILLER_52_882 ();
 FILLCELL_X2 FILLER_52_892 ();
 FILLCELL_X8 FILLER_52_904 ();
 FILLCELL_X16 FILLER_52_920 ();
 FILLCELL_X4 FILLER_52_936 ();
 FILLCELL_X2 FILLER_52_940 ();
 FILLCELL_X1 FILLER_52_942 ();
 FILLCELL_X4 FILLER_52_953 ();
 FILLCELL_X1 FILLER_52_957 ();
 FILLCELL_X8 FILLER_52_970 ();
 FILLCELL_X4 FILLER_52_978 ();
 FILLCELL_X2 FILLER_52_982 ();
 FILLCELL_X1 FILLER_52_984 ();
 FILLCELL_X8 FILLER_52_1014 ();
 FILLCELL_X4 FILLER_52_1022 ();
 FILLCELL_X1 FILLER_52_1026 ();
 FILLCELL_X4 FILLER_52_1040 ();
 FILLCELL_X2 FILLER_52_1044 ();
 FILLCELL_X2 FILLER_52_1063 ();
 FILLCELL_X4 FILLER_52_1069 ();
 FILLCELL_X4 FILLER_52_1090 ();
 FILLCELL_X2 FILLER_52_1094 ();
 FILLCELL_X1 FILLER_52_1096 ();
 FILLCELL_X8 FILLER_52_1111 ();
 FILLCELL_X4 FILLER_52_1119 ();
 FILLCELL_X1 FILLER_52_1123 ();
 FILLCELL_X8 FILLER_52_1148 ();
 FILLCELL_X2 FILLER_52_1156 ();
 FILLCELL_X1 FILLER_52_1158 ();
 FILLCELL_X4 FILLER_52_1202 ();
 FILLCELL_X1 FILLER_52_1209 ();
 FILLCELL_X1 FILLER_52_1217 ();
 FILLCELL_X2 FILLER_52_1231 ();
 FILLCELL_X1 FILLER_52_1233 ();
 FILLCELL_X2 FILLER_52_1237 ();
 FILLCELL_X1 FILLER_52_1239 ();
 FILLCELL_X8 FILLER_53_1 ();
 FILLCELL_X2 FILLER_53_9 ();
 FILLCELL_X1 FILLER_53_11 ();
 FILLCELL_X4 FILLER_53_33 ();
 FILLCELL_X2 FILLER_53_37 ();
 FILLCELL_X2 FILLER_53_46 ();
 FILLCELL_X4 FILLER_53_55 ();
 FILLCELL_X2 FILLER_53_59 ();
 FILLCELL_X1 FILLER_53_61 ();
 FILLCELL_X32 FILLER_53_76 ();
 FILLCELL_X32 FILLER_53_108 ();
 FILLCELL_X1 FILLER_53_140 ();
 FILLCELL_X8 FILLER_53_165 ();
 FILLCELL_X4 FILLER_53_202 ();
 FILLCELL_X2 FILLER_53_206 ();
 FILLCELL_X4 FILLER_53_246 ();
 FILLCELL_X2 FILLER_53_250 ();
 FILLCELL_X1 FILLER_53_252 ();
 FILLCELL_X16 FILLER_53_266 ();
 FILLCELL_X8 FILLER_53_282 ();
 FILLCELL_X4 FILLER_53_290 ();
 FILLCELL_X4 FILLER_53_308 ();
 FILLCELL_X4 FILLER_53_319 ();
 FILLCELL_X4 FILLER_53_327 ();
 FILLCELL_X1 FILLER_53_331 ();
 FILLCELL_X2 FILLER_53_339 ();
 FILLCELL_X1 FILLER_53_341 ();
 FILLCELL_X2 FILLER_53_373 ();
 FILLCELL_X1 FILLER_53_375 ();
 FILLCELL_X16 FILLER_53_383 ();
 FILLCELL_X8 FILLER_53_399 ();
 FILLCELL_X2 FILLER_53_407 ();
 FILLCELL_X1 FILLER_53_423 ();
 FILLCELL_X16 FILLER_53_431 ();
 FILLCELL_X4 FILLER_53_447 ();
 FILLCELL_X1 FILLER_53_451 ();
 FILLCELL_X8 FILLER_53_476 ();
 FILLCELL_X1 FILLER_53_484 ();
 FILLCELL_X4 FILLER_53_492 ();
 FILLCELL_X1 FILLER_53_496 ();
 FILLCELL_X8 FILLER_53_521 ();
 FILLCELL_X2 FILLER_53_529 ();
 FILLCELL_X4 FILLER_53_538 ();
 FILLCELL_X2 FILLER_53_542 ();
 FILLCELL_X1 FILLER_53_544 ();
 FILLCELL_X32 FILLER_53_562 ();
 FILLCELL_X32 FILLER_53_594 ();
 FILLCELL_X4 FILLER_53_626 ();
 FILLCELL_X2 FILLER_53_630 ();
 FILLCELL_X1 FILLER_53_632 ();
 FILLCELL_X4 FILLER_53_650 ();
 FILLCELL_X1 FILLER_53_661 ();
 FILLCELL_X4 FILLER_53_669 ();
 FILLCELL_X2 FILLER_53_673 ();
 FILLCELL_X1 FILLER_53_712 ();
 FILLCELL_X4 FILLER_53_726 ();
 FILLCELL_X1 FILLER_53_730 ();
 FILLCELL_X1 FILLER_53_738 ();
 FILLCELL_X1 FILLER_53_752 ();
 FILLCELL_X1 FILLER_53_757 ();
 FILLCELL_X2 FILLER_53_768 ();
 FILLCELL_X1 FILLER_53_770 ();
 FILLCELL_X8 FILLER_53_774 ();
 FILLCELL_X4 FILLER_53_782 ();
 FILLCELL_X1 FILLER_53_786 ();
 FILLCELL_X8 FILLER_53_790 ();
 FILLCELL_X2 FILLER_53_805 ();
 FILLCELL_X1 FILLER_53_807 ();
 FILLCELL_X8 FILLER_53_811 ();
 FILLCELL_X2 FILLER_53_825 ();
 FILLCELL_X1 FILLER_53_827 ();
 FILLCELL_X2 FILLER_53_831 ();
 FILLCELL_X1 FILLER_53_833 ();
 FILLCELL_X8 FILLER_53_842 ();
 FILLCELL_X4 FILLER_53_850 ();
 FILLCELL_X1 FILLER_53_854 ();
 FILLCELL_X4 FILLER_53_866 ();
 FILLCELL_X1 FILLER_53_873 ();
 FILLCELL_X1 FILLER_53_896 ();
 FILLCELL_X2 FILLER_53_906 ();
 FILLCELL_X1 FILLER_53_913 ();
 FILLCELL_X2 FILLER_53_919 ();
 FILLCELL_X8 FILLER_53_930 ();
 FILLCELL_X2 FILLER_53_938 ();
 FILLCELL_X16 FILLER_53_945 ();
 FILLCELL_X1 FILLER_53_961 ();
 FILLCELL_X2 FILLER_53_972 ();
 FILLCELL_X1 FILLER_53_974 ();
 FILLCELL_X1 FILLER_53_978 ();
 FILLCELL_X16 FILLER_53_1027 ();
 FILLCELL_X4 FILLER_53_1043 ();
 FILLCELL_X2 FILLER_53_1047 ();
 FILLCELL_X4 FILLER_53_1063 ();
 FILLCELL_X2 FILLER_53_1067 ();
 FILLCELL_X4 FILLER_53_1117 ();
 FILLCELL_X1 FILLER_53_1121 ();
 FILLCELL_X16 FILLER_53_1146 ();
 FILLCELL_X4 FILLER_53_1162 ();
 FILLCELL_X8 FILLER_53_1180 ();
 FILLCELL_X2 FILLER_53_1188 ();
 FILLCELL_X8 FILLER_53_1194 ();
 FILLCELL_X4 FILLER_53_1202 ();
 FILLCELL_X2 FILLER_53_1206 ();
 FILLCELL_X16 FILLER_54_1 ();
 FILLCELL_X8 FILLER_54_17 ();
 FILLCELL_X4 FILLER_54_25 ();
 FILLCELL_X32 FILLER_54_46 ();
 FILLCELL_X8 FILLER_54_78 ();
 FILLCELL_X2 FILLER_54_86 ();
 FILLCELL_X1 FILLER_54_88 ();
 FILLCELL_X4 FILLER_54_106 ();
 FILLCELL_X2 FILLER_54_127 ();
 FILLCELL_X2 FILLER_54_136 ();
 FILLCELL_X1 FILLER_54_138 ();
 FILLCELL_X1 FILLER_54_146 ();
 FILLCELL_X2 FILLER_54_164 ();
 FILLCELL_X1 FILLER_54_166 ();
 FILLCELL_X2 FILLER_54_181 ();
 FILLCELL_X1 FILLER_54_183 ();
 FILLCELL_X1 FILLER_54_191 ();
 FILLCELL_X32 FILLER_54_209 ();
 FILLCELL_X16 FILLER_54_241 ();
 FILLCELL_X8 FILLER_54_257 ();
 FILLCELL_X4 FILLER_54_282 ();
 FILLCELL_X1 FILLER_54_310 ();
 FILLCELL_X8 FILLER_54_328 ();
 FILLCELL_X4 FILLER_54_343 ();
 FILLCELL_X4 FILLER_54_352 ();
 FILLCELL_X2 FILLER_54_363 ();
 FILLCELL_X16 FILLER_54_379 ();
 FILLCELL_X8 FILLER_54_395 ();
 FILLCELL_X2 FILLER_54_403 ();
 FILLCELL_X32 FILLER_54_422 ();
 FILLCELL_X4 FILLER_54_454 ();
 FILLCELL_X2 FILLER_54_458 ();
 FILLCELL_X1 FILLER_54_460 ();
 FILLCELL_X4 FILLER_54_492 ();
 FILLCELL_X2 FILLER_54_496 ();
 FILLCELL_X2 FILLER_54_505 ();
 FILLCELL_X1 FILLER_54_507 ();
 FILLCELL_X2 FILLER_54_518 ();
 FILLCELL_X32 FILLER_54_534 ();
 FILLCELL_X16 FILLER_54_566 ();
 FILLCELL_X8 FILLER_54_582 ();
 FILLCELL_X16 FILLER_54_614 ();
 FILLCELL_X1 FILLER_54_630 ();
 FILLCELL_X2 FILLER_54_632 ();
 FILLCELL_X1 FILLER_54_634 ();
 FILLCELL_X16 FILLER_54_683 ();
 FILLCELL_X2 FILLER_54_699 ();
 FILLCELL_X32 FILLER_54_706 ();
 FILLCELL_X8 FILLER_54_738 ();
 FILLCELL_X2 FILLER_54_746 ();
 FILLCELL_X1 FILLER_54_748 ();
 FILLCELL_X2 FILLER_54_766 ();
 FILLCELL_X4 FILLER_54_774 ();
 FILLCELL_X2 FILLER_54_778 ();
 FILLCELL_X8 FILLER_54_803 ();
 FILLCELL_X1 FILLER_54_811 ();
 FILLCELL_X1 FILLER_54_818 ();
 FILLCELL_X2 FILLER_54_865 ();
 FILLCELL_X2 FILLER_54_880 ();
 FILLCELL_X1 FILLER_54_914 ();
 FILLCELL_X1 FILLER_54_924 ();
 FILLCELL_X1 FILLER_54_928 ();
 FILLCELL_X2 FILLER_54_932 ();
 FILLCELL_X1 FILLER_54_949 ();
 FILLCELL_X4 FILLER_54_954 ();
 FILLCELL_X2 FILLER_54_958 ();
 FILLCELL_X8 FILLER_54_981 ();
 FILLCELL_X2 FILLER_54_989 ();
 FILLCELL_X2 FILLER_54_1037 ();
 FILLCELL_X4 FILLER_54_1063 ();
 FILLCELL_X1 FILLER_54_1091 ();
 FILLCELL_X2 FILLER_54_1109 ();
 FILLCELL_X2 FILLER_54_1128 ();
 FILLCELL_X16 FILLER_54_1139 ();
 FILLCELL_X2 FILLER_54_1155 ();
 FILLCELL_X1 FILLER_54_1157 ();
 FILLCELL_X1 FILLER_54_1165 ();
 FILLCELL_X16 FILLER_54_1179 ();
 FILLCELL_X1 FILLER_54_1195 ();
 FILLCELL_X1 FILLER_54_1239 ();
 FILLCELL_X8 FILLER_55_1 ();
 FILLCELL_X4 FILLER_55_9 ();
 FILLCELL_X2 FILLER_55_13 ();
 FILLCELL_X1 FILLER_55_15 ();
 FILLCELL_X8 FILLER_55_42 ();
 FILLCELL_X4 FILLER_55_50 ();
 FILLCELL_X2 FILLER_55_54 ();
 FILLCELL_X4 FILLER_55_80 ();
 FILLCELL_X2 FILLER_55_84 ();
 FILLCELL_X1 FILLER_55_86 ();
 FILLCELL_X2 FILLER_55_94 ();
 FILLCELL_X1 FILLER_55_96 ();
 FILLCELL_X2 FILLER_55_114 ();
 FILLCELL_X1 FILLER_55_116 ();
 FILLCELL_X2 FILLER_55_124 ();
 FILLCELL_X2 FILLER_55_133 ();
 FILLCELL_X8 FILLER_55_142 ();
 FILLCELL_X1 FILLER_55_150 ();
 FILLCELL_X16 FILLER_55_156 ();
 FILLCELL_X8 FILLER_55_172 ();
 FILLCELL_X2 FILLER_55_180 ();
 FILLCELL_X1 FILLER_55_182 ();
 FILLCELL_X2 FILLER_55_196 ();
 FILLCELL_X1 FILLER_55_198 ();
 FILLCELL_X8 FILLER_55_206 ();
 FILLCELL_X2 FILLER_55_214 ();
 FILLCELL_X4 FILLER_55_223 ();
 FILLCELL_X4 FILLER_55_234 ();
 FILLCELL_X2 FILLER_55_238 ();
 FILLCELL_X1 FILLER_55_240 ();
 FILLCELL_X8 FILLER_55_258 ();
 FILLCELL_X1 FILLER_55_266 ();
 FILLCELL_X1 FILLER_55_308 ();
 FILLCELL_X2 FILLER_55_312 ();
 FILLCELL_X4 FILLER_55_328 ();
 FILLCELL_X1 FILLER_55_332 ();
 FILLCELL_X8 FILLER_55_357 ();
 FILLCELL_X4 FILLER_55_365 ();
 FILLCELL_X2 FILLER_55_369 ();
 FILLCELL_X16 FILLER_55_378 ();
 FILLCELL_X32 FILLER_55_397 ();
 FILLCELL_X16 FILLER_55_429 ();
 FILLCELL_X4 FILLER_55_445 ();
 FILLCELL_X2 FILLER_55_449 ();
 FILLCELL_X8 FILLER_55_478 ();
 FILLCELL_X2 FILLER_55_486 ();
 FILLCELL_X2 FILLER_55_494 ();
 FILLCELL_X4 FILLER_55_519 ();
 FILLCELL_X8 FILLER_55_560 ();
 FILLCELL_X4 FILLER_55_568 ();
 FILLCELL_X1 FILLER_55_572 ();
 FILLCELL_X2 FILLER_55_590 ();
 FILLCELL_X4 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_630 ();
 FILLCELL_X8 FILLER_55_662 ();
 FILLCELL_X4 FILLER_55_670 ();
 FILLCELL_X1 FILLER_55_674 ();
 FILLCELL_X1 FILLER_55_682 ();
 FILLCELL_X16 FILLER_55_696 ();
 FILLCELL_X8 FILLER_55_712 ();
 FILLCELL_X16 FILLER_55_768 ();
 FILLCELL_X1 FILLER_55_784 ();
 FILLCELL_X4 FILLER_55_789 ();
 FILLCELL_X8 FILLER_55_800 ();
 FILLCELL_X2 FILLER_55_808 ();
 FILLCELL_X2 FILLER_55_820 ();
 FILLCELL_X4 FILLER_55_850 ();
 FILLCELL_X2 FILLER_55_854 ();
 FILLCELL_X1 FILLER_55_856 ();
 FILLCELL_X1 FILLER_55_867 ();
 FILLCELL_X2 FILLER_55_871 ();
 FILLCELL_X1 FILLER_55_878 ();
 FILLCELL_X2 FILLER_55_884 ();
 FILLCELL_X4 FILLER_55_895 ();
 FILLCELL_X2 FILLER_55_899 ();
 FILLCELL_X1 FILLER_55_901 ();
 FILLCELL_X4 FILLER_55_916 ();
 FILLCELL_X2 FILLER_55_920 ();
 FILLCELL_X1 FILLER_55_948 ();
 FILLCELL_X8 FILLER_55_954 ();
 FILLCELL_X1 FILLER_55_962 ();
 FILLCELL_X1 FILLER_55_981 ();
 FILLCELL_X8 FILLER_55_986 ();
 FILLCELL_X8 FILLER_55_1015 ();
 FILLCELL_X4 FILLER_55_1023 ();
 FILLCELL_X2 FILLER_55_1027 ();
 FILLCELL_X1 FILLER_55_1046 ();
 FILLCELL_X8 FILLER_55_1068 ();
 FILLCELL_X2 FILLER_55_1076 ();
 FILLCELL_X1 FILLER_55_1078 ();
 FILLCELL_X2 FILLER_55_1086 ();
 FILLCELL_X16 FILLER_55_1134 ();
 FILLCELL_X2 FILLER_55_1150 ();
 FILLCELL_X1 FILLER_55_1176 ();
 FILLCELL_X2 FILLER_55_1194 ();
 FILLCELL_X2 FILLER_55_1217 ();
 FILLCELL_X1 FILLER_55_1219 ();
 FILLCELL_X16 FILLER_56_1 ();
 FILLCELL_X4 FILLER_56_17 ();
 FILLCELL_X1 FILLER_56_39 ();
 FILLCELL_X16 FILLER_56_47 ();
 FILLCELL_X1 FILLER_56_63 ();
 FILLCELL_X4 FILLER_56_92 ();
 FILLCELL_X2 FILLER_56_103 ();
 FILLCELL_X1 FILLER_56_105 ();
 FILLCELL_X8 FILLER_56_113 ();
 FILLCELL_X4 FILLER_56_121 ();
 FILLCELL_X2 FILLER_56_142 ();
 FILLCELL_X2 FILLER_56_161 ();
 FILLCELL_X2 FILLER_56_170 ();
 FILLCELL_X1 FILLER_56_172 ();
 FILLCELL_X4 FILLER_56_190 ();
 FILLCELL_X2 FILLER_56_194 ();
 FILLCELL_X4 FILLER_56_237 ();
 FILLCELL_X2 FILLER_56_241 ();
 FILLCELL_X1 FILLER_56_243 ();
 FILLCELL_X8 FILLER_56_261 ();
 FILLCELL_X2 FILLER_56_269 ();
 FILLCELL_X1 FILLER_56_271 ();
 FILLCELL_X1 FILLER_56_279 ();
 FILLCELL_X4 FILLER_56_294 ();
 FILLCELL_X2 FILLER_56_298 ();
 FILLCELL_X2 FILLER_56_307 ();
 FILLCELL_X4 FILLER_56_340 ();
 FILLCELL_X2 FILLER_56_344 ();
 FILLCELL_X8 FILLER_56_359 ();
 FILLCELL_X4 FILLER_56_367 ();
 FILLCELL_X1 FILLER_56_371 ();
 FILLCELL_X16 FILLER_56_389 ();
 FILLCELL_X2 FILLER_56_405 ();
 FILLCELL_X1 FILLER_56_407 ();
 FILLCELL_X16 FILLER_56_415 ();
 FILLCELL_X4 FILLER_56_431 ();
 FILLCELL_X16 FILLER_56_443 ();
 FILLCELL_X1 FILLER_56_459 ();
 FILLCELL_X2 FILLER_56_472 ();
 FILLCELL_X16 FILLER_56_496 ();
 FILLCELL_X4 FILLER_56_512 ();
 FILLCELL_X1 FILLER_56_516 ();
 FILLCELL_X4 FILLER_56_546 ();
 FILLCELL_X1 FILLER_56_550 ();
 FILLCELL_X4 FILLER_56_558 ();
 FILLCELL_X2 FILLER_56_562 ();
 FILLCELL_X1 FILLER_56_564 ();
 FILLCELL_X8 FILLER_56_579 ();
 FILLCELL_X4 FILLER_56_587 ();
 FILLCELL_X1 FILLER_56_591 ();
 FILLCELL_X8 FILLER_56_620 ();
 FILLCELL_X2 FILLER_56_628 ();
 FILLCELL_X1 FILLER_56_630 ();
 FILLCELL_X8 FILLER_56_632 ();
 FILLCELL_X4 FILLER_56_640 ();
 FILLCELL_X1 FILLER_56_644 ();
 FILLCELL_X2 FILLER_56_669 ();
 FILLCELL_X4 FILLER_56_685 ();
 FILLCELL_X2 FILLER_56_689 ();
 FILLCELL_X1 FILLER_56_691 ();
 FILLCELL_X16 FILLER_56_696 ();
 FILLCELL_X1 FILLER_56_712 ();
 FILLCELL_X4 FILLER_56_730 ();
 FILLCELL_X2 FILLER_56_734 ();
 FILLCELL_X1 FILLER_56_736 ();
 FILLCELL_X1 FILLER_56_744 ();
 FILLCELL_X1 FILLER_56_752 ();
 FILLCELL_X16 FILLER_56_757 ();
 FILLCELL_X8 FILLER_56_773 ();
 FILLCELL_X8 FILLER_56_801 ();
 FILLCELL_X4 FILLER_56_809 ();
 FILLCELL_X2 FILLER_56_813 ();
 FILLCELL_X2 FILLER_56_841 ();
 FILLCELL_X4 FILLER_56_858 ();
 FILLCELL_X4 FILLER_56_872 ();
 FILLCELL_X2 FILLER_56_876 ();
 FILLCELL_X4 FILLER_56_883 ();
 FILLCELL_X2 FILLER_56_887 ();
 FILLCELL_X8 FILLER_56_915 ();
 FILLCELL_X1 FILLER_56_923 ();
 FILLCELL_X32 FILLER_56_933 ();
 FILLCELL_X8 FILLER_56_965 ();
 FILLCELL_X1 FILLER_56_973 ();
 FILLCELL_X16 FILLER_56_984 ();
 FILLCELL_X4 FILLER_56_1000 ();
 FILLCELL_X1 FILLER_56_1004 ();
 FILLCELL_X8 FILLER_56_1008 ();
 FILLCELL_X2 FILLER_56_1016 ();
 FILLCELL_X1 FILLER_56_1018 ();
 FILLCELL_X16 FILLER_56_1043 ();
 FILLCELL_X8 FILLER_56_1059 ();
 FILLCELL_X4 FILLER_56_1067 ();
 FILLCELL_X2 FILLER_56_1071 ();
 FILLCELL_X8 FILLER_56_1086 ();
 FILLCELL_X4 FILLER_56_1094 ();
 FILLCELL_X2 FILLER_56_1098 ();
 FILLCELL_X1 FILLER_56_1100 ();
 FILLCELL_X4 FILLER_56_1106 ();
 FILLCELL_X2 FILLER_56_1110 ();
 FILLCELL_X1 FILLER_56_1112 ();
 FILLCELL_X8 FILLER_56_1137 ();
 FILLCELL_X4 FILLER_56_1145 ();
 FILLCELL_X1 FILLER_56_1149 ();
 FILLCELL_X1 FILLER_56_1167 ();
 FILLCELL_X2 FILLER_56_1206 ();
 FILLCELL_X1 FILLER_56_1221 ();
 FILLCELL_X16 FILLER_57_5 ();
 FILLCELL_X8 FILLER_57_21 ();
 FILLCELL_X8 FILLER_57_46 ();
 FILLCELL_X1 FILLER_57_54 ();
 FILLCELL_X4 FILLER_57_62 ();
 FILLCELL_X2 FILLER_57_66 ();
 FILLCELL_X1 FILLER_57_68 ();
 FILLCELL_X1 FILLER_57_76 ();
 FILLCELL_X8 FILLER_57_89 ();
 FILLCELL_X2 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_103 ();
 FILLCELL_X8 FILLER_57_135 ();
 FILLCELL_X1 FILLER_57_150 ();
 FILLCELL_X8 FILLER_57_154 ();
 FILLCELL_X2 FILLER_57_169 ();
 FILLCELL_X2 FILLER_57_178 ();
 FILLCELL_X1 FILLER_57_187 ();
 FILLCELL_X2 FILLER_57_205 ();
 FILLCELL_X4 FILLER_57_214 ();
 FILLCELL_X2 FILLER_57_225 ();
 FILLCELL_X2 FILLER_57_240 ();
 FILLCELL_X32 FILLER_57_263 ();
 FILLCELL_X4 FILLER_57_295 ();
 FILLCELL_X2 FILLER_57_299 ();
 FILLCELL_X8 FILLER_57_306 ();
 FILLCELL_X2 FILLER_57_314 ();
 FILLCELL_X16 FILLER_57_319 ();
 FILLCELL_X8 FILLER_57_335 ();
 FILLCELL_X1 FILLER_57_343 ();
 FILLCELL_X16 FILLER_57_378 ();
 FILLCELL_X2 FILLER_57_394 ();
 FILLCELL_X1 FILLER_57_396 ();
 FILLCELL_X4 FILLER_57_445 ();
 FILLCELL_X2 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_482 ();
 FILLCELL_X1 FILLER_57_514 ();
 FILLCELL_X2 FILLER_57_532 ();
 FILLCELL_X4 FILLER_57_558 ();
 FILLCELL_X1 FILLER_57_562 ();
 FILLCELL_X16 FILLER_57_575 ();
 FILLCELL_X8 FILLER_57_591 ();
 FILLCELL_X2 FILLER_57_599 ();
 FILLCELL_X1 FILLER_57_601 ();
 FILLCELL_X1 FILLER_57_605 ();
 FILLCELL_X2 FILLER_57_613 ();
 FILLCELL_X1 FILLER_57_615 ();
 FILLCELL_X8 FILLER_57_640 ();
 FILLCELL_X4 FILLER_57_655 ();
 FILLCELL_X1 FILLER_57_676 ();
 FILLCELL_X4 FILLER_57_691 ();
 FILLCELL_X8 FILLER_57_708 ();
 FILLCELL_X8 FILLER_57_733 ();
 FILLCELL_X2 FILLER_57_741 ();
 FILLCELL_X1 FILLER_57_774 ();
 FILLCELL_X2 FILLER_57_787 ();
 FILLCELL_X1 FILLER_57_789 ();
 FILLCELL_X16 FILLER_57_799 ();
 FILLCELL_X8 FILLER_57_815 ();
 FILLCELL_X4 FILLER_57_823 ();
 FILLCELL_X1 FILLER_57_827 ();
 FILLCELL_X16 FILLER_57_833 ();
 FILLCELL_X2 FILLER_57_849 ();
 FILLCELL_X1 FILLER_57_851 ();
 FILLCELL_X2 FILLER_57_857 ();
 FILLCELL_X2 FILLER_57_867 ();
 FILLCELL_X2 FILLER_57_872 ();
 FILLCELL_X4 FILLER_57_887 ();
 FILLCELL_X2 FILLER_57_891 ();
 FILLCELL_X8 FILLER_57_900 ();
 FILLCELL_X4 FILLER_57_908 ();
 FILLCELL_X2 FILLER_57_912 ();
 FILLCELL_X1 FILLER_57_914 ();
 FILLCELL_X8 FILLER_57_920 ();
 FILLCELL_X2 FILLER_57_928 ();
 FILLCELL_X1 FILLER_57_930 ();
 FILLCELL_X8 FILLER_57_941 ();
 FILLCELL_X8 FILLER_57_954 ();
 FILLCELL_X2 FILLER_57_962 ();
 FILLCELL_X2 FILLER_57_969 ();
 FILLCELL_X1 FILLER_57_971 ();
 FILLCELL_X1 FILLER_57_978 ();
 FILLCELL_X4 FILLER_57_986 ();
 FILLCELL_X1 FILLER_57_990 ();
 FILLCELL_X16 FILLER_57_996 ();
 FILLCELL_X4 FILLER_57_1012 ();
 FILLCELL_X1 FILLER_57_1016 ();
 FILLCELL_X1 FILLER_57_1022 ();
 FILLCELL_X4 FILLER_57_1037 ();
 FILLCELL_X16 FILLER_57_1078 ();
 FILLCELL_X8 FILLER_57_1094 ();
 FILLCELL_X2 FILLER_57_1102 ();
 FILLCELL_X2 FILLER_57_1128 ();
 FILLCELL_X16 FILLER_57_1137 ();
 FILLCELL_X2 FILLER_57_1153 ();
 FILLCELL_X4 FILLER_57_1182 ();
 FILLCELL_X2 FILLER_57_1186 ();
 FILLCELL_X1 FILLER_57_1188 ();
 FILLCELL_X8 FILLER_57_1193 ();
 FILLCELL_X2 FILLER_57_1201 ();
 FILLCELL_X2 FILLER_57_1231 ();
 FILLCELL_X1 FILLER_57_1233 ();
 FILLCELL_X2 FILLER_57_1237 ();
 FILLCELL_X1 FILLER_57_1239 ();
 FILLCELL_X4 FILLER_58_1 ();
 FILLCELL_X2 FILLER_58_29 ();
 FILLCELL_X2 FILLER_58_38 ();
 FILLCELL_X1 FILLER_58_40 ();
 FILLCELL_X2 FILLER_58_65 ();
 FILLCELL_X1 FILLER_58_67 ();
 FILLCELL_X8 FILLER_58_75 ();
 FILLCELL_X4 FILLER_58_83 ();
 FILLCELL_X1 FILLER_58_87 ();
 FILLCELL_X32 FILLER_58_112 ();
 FILLCELL_X8 FILLER_58_144 ();
 FILLCELL_X2 FILLER_58_152 ();
 FILLCELL_X1 FILLER_58_154 ();
 FILLCELL_X4 FILLER_58_172 ();
 FILLCELL_X1 FILLER_58_176 ();
 FILLCELL_X2 FILLER_58_191 ();
 FILLCELL_X32 FILLER_58_196 ();
 FILLCELL_X16 FILLER_58_228 ();
 FILLCELL_X1 FILLER_58_244 ();
 FILLCELL_X16 FILLER_58_259 ();
 FILLCELL_X8 FILLER_58_275 ();
 FILLCELL_X4 FILLER_58_283 ();
 FILLCELL_X2 FILLER_58_287 ();
 FILLCELL_X32 FILLER_58_296 ();
 FILLCELL_X8 FILLER_58_328 ();
 FILLCELL_X2 FILLER_58_336 ();
 FILLCELL_X4 FILLER_58_345 ();
 FILLCELL_X1 FILLER_58_349 ();
 FILLCELL_X4 FILLER_58_357 ();
 FILLCELL_X2 FILLER_58_361 ();
 FILLCELL_X1 FILLER_58_363 ();
 FILLCELL_X8 FILLER_58_378 ();
 FILLCELL_X2 FILLER_58_386 ();
 FILLCELL_X1 FILLER_58_412 ();
 FILLCELL_X2 FILLER_58_454 ();
 FILLCELL_X2 FILLER_58_460 ();
 FILLCELL_X1 FILLER_58_462 ();
 FILLCELL_X16 FILLER_58_480 ();
 FILLCELL_X4 FILLER_58_496 ();
 FILLCELL_X4 FILLER_58_531 ();
 FILLCELL_X4 FILLER_58_549 ();
 FILLCELL_X1 FILLER_58_553 ();
 FILLCELL_X8 FILLER_58_586 ();
 FILLCELL_X2 FILLER_58_594 ();
 FILLCELL_X8 FILLER_58_618 ();
 FILLCELL_X4 FILLER_58_626 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X4 FILLER_58_632 ();
 FILLCELL_X16 FILLER_58_661 ();
 FILLCELL_X2 FILLER_58_677 ();
 FILLCELL_X1 FILLER_58_679 ();
 FILLCELL_X1 FILLER_58_704 ();
 FILLCELL_X2 FILLER_58_743 ();
 FILLCELL_X16 FILLER_58_749 ();
 FILLCELL_X4 FILLER_58_765 ();
 FILLCELL_X2 FILLER_58_769 ();
 FILLCELL_X1 FILLER_58_771 ();
 FILLCELL_X8 FILLER_58_779 ();
 FILLCELL_X4 FILLER_58_804 ();
 FILLCELL_X32 FILLER_58_820 ();
 FILLCELL_X4 FILLER_58_852 ();
 FILLCELL_X2 FILLER_58_890 ();
 FILLCELL_X8 FILLER_58_897 ();
 FILLCELL_X1 FILLER_58_922 ();
 FILLCELL_X8 FILLER_58_953 ();
 FILLCELL_X2 FILLER_58_961 ();
 FILLCELL_X1 FILLER_58_963 ();
 FILLCELL_X8 FILLER_58_987 ();
 FILLCELL_X4 FILLER_58_995 ();
 FILLCELL_X2 FILLER_58_1033 ();
 FILLCELL_X16 FILLER_58_1082 ();
 FILLCELL_X8 FILLER_58_1098 ();
 FILLCELL_X2 FILLER_58_1106 ();
 FILLCELL_X2 FILLER_58_1115 ();
 FILLCELL_X1 FILLER_58_1117 ();
 FILLCELL_X32 FILLER_58_1149 ();
 FILLCELL_X4 FILLER_58_1181 ();
 FILLCELL_X2 FILLER_58_1185 ();
 FILLCELL_X4 FILLER_58_1207 ();
 FILLCELL_X2 FILLER_58_1211 ();
 FILLCELL_X1 FILLER_58_1213 ();
 FILLCELL_X1 FILLER_58_1223 ();
 FILLCELL_X16 FILLER_59_1 ();
 FILLCELL_X8 FILLER_59_17 ();
 FILLCELL_X1 FILLER_59_25 ();
 FILLCELL_X8 FILLER_59_43 ();
 FILLCELL_X4 FILLER_59_51 ();
 FILLCELL_X1 FILLER_59_55 ();
 FILLCELL_X1 FILLER_59_73 ();
 FILLCELL_X16 FILLER_59_81 ();
 FILLCELL_X4 FILLER_59_97 ();
 FILLCELL_X1 FILLER_59_101 ();
 FILLCELL_X2 FILLER_59_109 ();
 FILLCELL_X1 FILLER_59_111 ();
 FILLCELL_X4 FILLER_59_126 ();
 FILLCELL_X1 FILLER_59_130 ();
 FILLCELL_X16 FILLER_59_152 ();
 FILLCELL_X8 FILLER_59_168 ();
 FILLCELL_X4 FILLER_59_176 ();
 FILLCELL_X8 FILLER_59_183 ();
 FILLCELL_X4 FILLER_59_191 ();
 FILLCELL_X1 FILLER_59_195 ();
 FILLCELL_X8 FILLER_59_203 ();
 FILLCELL_X4 FILLER_59_211 ();
 FILLCELL_X1 FILLER_59_215 ();
 FILLCELL_X4 FILLER_59_233 ();
 FILLCELL_X2 FILLER_59_237 ();
 FILLCELL_X1 FILLER_59_246 ();
 FILLCELL_X8 FILLER_59_271 ();
 FILLCELL_X2 FILLER_59_279 ();
 FILLCELL_X2 FILLER_59_298 ();
 FILLCELL_X8 FILLER_59_317 ();
 FILLCELL_X2 FILLER_59_356 ();
 FILLCELL_X2 FILLER_59_366 ();
 FILLCELL_X16 FILLER_59_375 ();
 FILLCELL_X2 FILLER_59_391 ();
 FILLCELL_X1 FILLER_59_393 ();
 FILLCELL_X2 FILLER_59_416 ();
 FILLCELL_X1 FILLER_59_418 ();
 FILLCELL_X4 FILLER_59_422 ();
 FILLCELL_X1 FILLER_59_426 ();
 FILLCELL_X16 FILLER_59_447 ();
 FILLCELL_X8 FILLER_59_463 ();
 FILLCELL_X2 FILLER_59_471 ();
 FILLCELL_X4 FILLER_59_480 ();
 FILLCELL_X2 FILLER_59_484 ();
 FILLCELL_X1 FILLER_59_486 ();
 FILLCELL_X8 FILLER_59_497 ();
 FILLCELL_X1 FILLER_59_505 ();
 FILLCELL_X32 FILLER_59_531 ();
 FILLCELL_X16 FILLER_59_577 ();
 FILLCELL_X1 FILLER_59_593 ();
 FILLCELL_X16 FILLER_59_618 ();
 FILLCELL_X1 FILLER_59_634 ();
 FILLCELL_X8 FILLER_59_642 ();
 FILLCELL_X4 FILLER_59_650 ();
 FILLCELL_X16 FILLER_59_661 ();
 FILLCELL_X4 FILLER_59_677 ();
 FILLCELL_X1 FILLER_59_681 ();
 FILLCELL_X32 FILLER_59_704 ();
 FILLCELL_X8 FILLER_59_736 ();
 FILLCELL_X1 FILLER_59_744 ();
 FILLCELL_X32 FILLER_59_776 ();
 FILLCELL_X1 FILLER_59_808 ();
 FILLCELL_X8 FILLER_59_829 ();
 FILLCELL_X8 FILLER_59_842 ();
 FILLCELL_X4 FILLER_59_850 ();
 FILLCELL_X2 FILLER_59_854 ();
 FILLCELL_X1 FILLER_59_873 ();
 FILLCELL_X2 FILLER_59_898 ();
 FILLCELL_X2 FILLER_59_937 ();
 FILLCELL_X1 FILLER_59_952 ();
 FILLCELL_X16 FILLER_59_962 ();
 FILLCELL_X8 FILLER_59_991 ();
 FILLCELL_X1 FILLER_59_999 ();
 FILLCELL_X2 FILLER_59_1033 ();
 FILLCELL_X4 FILLER_59_1039 ();
 FILLCELL_X2 FILLER_59_1043 ();
 FILLCELL_X2 FILLER_59_1062 ();
 FILLCELL_X1 FILLER_59_1064 ();
 FILLCELL_X4 FILLER_59_1072 ();
 FILLCELL_X1 FILLER_59_1076 ();
 FILLCELL_X4 FILLER_59_1094 ();
 FILLCELL_X1 FILLER_59_1098 ();
 FILLCELL_X32 FILLER_59_1136 ();
 FILLCELL_X1 FILLER_59_1168 ();
 FILLCELL_X8 FILLER_59_1184 ();
 FILLCELL_X4 FILLER_59_1192 ();
 FILLCELL_X1 FILLER_59_1196 ();
 FILLCELL_X1 FILLER_59_1204 ();
 FILLCELL_X1 FILLER_59_1236 ();
 FILLCELL_X8 FILLER_60_1 ();
 FILLCELL_X4 FILLER_60_9 ();
 FILLCELL_X32 FILLER_60_17 ();
 FILLCELL_X8 FILLER_60_49 ();
 FILLCELL_X1 FILLER_60_57 ();
 FILLCELL_X4 FILLER_60_63 ();
 FILLCELL_X8 FILLER_60_74 ();
 FILLCELL_X4 FILLER_60_82 ();
 FILLCELL_X1 FILLER_60_86 ();
 FILLCELL_X4 FILLER_60_92 ();
 FILLCELL_X2 FILLER_60_96 ();
 FILLCELL_X8 FILLER_60_149 ();
 FILLCELL_X8 FILLER_60_169 ();
 FILLCELL_X8 FILLER_60_182 ();
 FILLCELL_X2 FILLER_60_190 ();
 FILLCELL_X16 FILLER_60_197 ();
 FILLCELL_X4 FILLER_60_213 ();
 FILLCELL_X2 FILLER_60_217 ();
 FILLCELL_X2 FILLER_60_226 ();
 FILLCELL_X1 FILLER_60_235 ();
 FILLCELL_X1 FILLER_60_256 ();
 FILLCELL_X1 FILLER_60_264 ();
 FILLCELL_X8 FILLER_60_269 ();
 FILLCELL_X2 FILLER_60_277 ();
 FILLCELL_X2 FILLER_60_303 ();
 FILLCELL_X1 FILLER_60_305 ();
 FILLCELL_X1 FILLER_60_323 ();
 FILLCELL_X8 FILLER_60_355 ();
 FILLCELL_X16 FILLER_60_377 ();
 FILLCELL_X8 FILLER_60_393 ();
 FILLCELL_X4 FILLER_60_401 ();
 FILLCELL_X1 FILLER_60_405 ();
 FILLCELL_X32 FILLER_60_409 ();
 FILLCELL_X32 FILLER_60_441 ();
 FILLCELL_X8 FILLER_60_473 ();
 FILLCELL_X2 FILLER_60_481 ();
 FILLCELL_X16 FILLER_60_500 ();
 FILLCELL_X4 FILLER_60_516 ();
 FILLCELL_X8 FILLER_60_557 ();
 FILLCELL_X4 FILLER_60_565 ();
 FILLCELL_X2 FILLER_60_569 ();
 FILLCELL_X1 FILLER_60_571 ();
 FILLCELL_X8 FILLER_60_589 ();
 FILLCELL_X4 FILLER_60_597 ();
 FILLCELL_X2 FILLER_60_601 ();
 FILLCELL_X4 FILLER_60_627 ();
 FILLCELL_X1 FILLER_60_632 ();
 FILLCELL_X4 FILLER_60_657 ();
 FILLCELL_X1 FILLER_60_661 ();
 FILLCELL_X16 FILLER_60_686 ();
 FILLCELL_X2 FILLER_60_702 ();
 FILLCELL_X1 FILLER_60_704 ();
 FILLCELL_X4 FILLER_60_712 ();
 FILLCELL_X2 FILLER_60_716 ();
 FILLCELL_X1 FILLER_60_718 ();
 FILLCELL_X16 FILLER_60_726 ();
 FILLCELL_X8 FILLER_60_742 ();
 FILLCELL_X2 FILLER_60_750 ();
 FILLCELL_X1 FILLER_60_752 ();
 FILLCELL_X16 FILLER_60_777 ();
 FILLCELL_X4 FILLER_60_793 ();
 FILLCELL_X2 FILLER_60_797 ();
 FILLCELL_X1 FILLER_60_799 ();
 FILLCELL_X2 FILLER_60_828 ();
 FILLCELL_X16 FILLER_60_835 ();
 FILLCELL_X8 FILLER_60_851 ();
 FILLCELL_X1 FILLER_60_859 ();
 FILLCELL_X8 FILLER_60_865 ();
 FILLCELL_X4 FILLER_60_873 ();
 FILLCELL_X16 FILLER_60_887 ();
 FILLCELL_X4 FILLER_60_903 ();
 FILLCELL_X2 FILLER_60_907 ();
 FILLCELL_X1 FILLER_60_909 ();
 FILLCELL_X2 FILLER_60_921 ();
 FILLCELL_X16 FILLER_60_926 ();
 FILLCELL_X1 FILLER_60_942 ();
 FILLCELL_X8 FILLER_60_951 ();
 FILLCELL_X4 FILLER_60_959 ();
 FILLCELL_X2 FILLER_60_963 ();
 FILLCELL_X1 FILLER_60_965 ();
 FILLCELL_X8 FILLER_60_990 ();
 FILLCELL_X4 FILLER_60_998 ();
 FILLCELL_X8 FILLER_60_1047 ();
 FILLCELL_X2 FILLER_60_1109 ();
 FILLCELL_X1 FILLER_60_1123 ();
 FILLCELL_X16 FILLER_60_1133 ();
 FILLCELL_X4 FILLER_60_1149 ();
 FILLCELL_X1 FILLER_60_1153 ();
 FILLCELL_X8 FILLER_60_1185 ();
 FILLCELL_X2 FILLER_60_1193 ();
 FILLCELL_X1 FILLER_60_1195 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X16 FILLER_61_33 ();
 FILLCELL_X2 FILLER_61_49 ();
 FILLCELL_X8 FILLER_61_75 ();
 FILLCELL_X2 FILLER_61_83 ();
 FILLCELL_X16 FILLER_61_102 ();
 FILLCELL_X2 FILLER_61_118 ();
 FILLCELL_X1 FILLER_61_120 ();
 FILLCELL_X16 FILLER_61_126 ();
 FILLCELL_X8 FILLER_61_142 ();
 FILLCELL_X2 FILLER_61_150 ();
 FILLCELL_X1 FILLER_61_152 ();
 FILLCELL_X1 FILLER_61_170 ();
 FILLCELL_X1 FILLER_61_219 ();
 FILLCELL_X1 FILLER_61_227 ();
 FILLCELL_X1 FILLER_61_235 ();
 FILLCELL_X1 FILLER_61_243 ();
 FILLCELL_X2 FILLER_61_251 ();
 FILLCELL_X8 FILLER_61_270 ();
 FILLCELL_X4 FILLER_61_278 ();
 FILLCELL_X2 FILLER_61_293 ();
 FILLCELL_X2 FILLER_61_330 ();
 FILLCELL_X1 FILLER_61_332 ();
 FILLCELL_X8 FILLER_61_385 ();
 FILLCELL_X4 FILLER_61_393 ();
 FILLCELL_X2 FILLER_61_421 ();
 FILLCELL_X8 FILLER_61_430 ();
 FILLCELL_X1 FILLER_61_438 ();
 FILLCELL_X8 FILLER_61_470 ();
 FILLCELL_X4 FILLER_61_478 ();
 FILLCELL_X2 FILLER_61_482 ();
 FILLCELL_X4 FILLER_61_508 ();
 FILLCELL_X1 FILLER_61_512 ();
 FILLCELL_X2 FILLER_61_516 ();
 FILLCELL_X1 FILLER_61_525 ();
 FILLCELL_X4 FILLER_61_550 ();
 FILLCELL_X2 FILLER_61_557 ();
 FILLCELL_X1 FILLER_61_559 ();
 FILLCELL_X4 FILLER_61_577 ();
 FILLCELL_X2 FILLER_61_581 ();
 FILLCELL_X2 FILLER_61_607 ();
 FILLCELL_X8 FILLER_61_633 ();
 FILLCELL_X4 FILLER_61_641 ();
 FILLCELL_X2 FILLER_61_645 ();
 FILLCELL_X1 FILLER_61_647 ();
 FILLCELL_X2 FILLER_61_672 ();
 FILLCELL_X16 FILLER_61_678 ();
 FILLCELL_X8 FILLER_61_694 ();
 FILLCELL_X32 FILLER_61_736 ();
 FILLCELL_X16 FILLER_61_768 ();
 FILLCELL_X8 FILLER_61_784 ();
 FILLCELL_X8 FILLER_61_797 ();
 FILLCELL_X8 FILLER_61_841 ();
 FILLCELL_X4 FILLER_61_849 ();
 FILLCELL_X8 FILLER_61_862 ();
 FILLCELL_X4 FILLER_61_870 ();
 FILLCELL_X1 FILLER_61_874 ();
 FILLCELL_X4 FILLER_61_880 ();
 FILLCELL_X1 FILLER_61_884 ();
 FILLCELL_X8 FILLER_61_890 ();
 FILLCELL_X4 FILLER_61_898 ();
 FILLCELL_X1 FILLER_61_912 ();
 FILLCELL_X4 FILLER_61_917 ();
 FILLCELL_X2 FILLER_61_921 ();
 FILLCELL_X2 FILLER_61_926 ();
 FILLCELL_X1 FILLER_61_928 ();
 FILLCELL_X32 FILLER_61_932 ();
 FILLCELL_X4 FILLER_61_964 ();
 FILLCELL_X1 FILLER_61_968 ();
 FILLCELL_X16 FILLER_61_979 ();
 FILLCELL_X8 FILLER_61_995 ();
 FILLCELL_X4 FILLER_61_1003 ();
 FILLCELL_X2 FILLER_61_1007 ();
 FILLCELL_X8 FILLER_61_1014 ();
 FILLCELL_X4 FILLER_61_1022 ();
 FILLCELL_X2 FILLER_61_1026 ();
 FILLCELL_X1 FILLER_61_1028 ();
 FILLCELL_X1 FILLER_61_1060 ();
 FILLCELL_X8 FILLER_61_1078 ();
 FILLCELL_X2 FILLER_61_1086 ();
 FILLCELL_X2 FILLER_61_1112 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X4 FILLER_61_1153 ();
 FILLCELL_X2 FILLER_61_1157 ();
 FILLCELL_X1 FILLER_61_1189 ();
 FILLCELL_X8 FILLER_61_1210 ();
 FILLCELL_X4 FILLER_61_1218 ();
 FILLCELL_X2 FILLER_61_1229 ();
 FILLCELL_X1 FILLER_61_1231 ();
 FILLCELL_X4 FILLER_61_1235 ();
 FILLCELL_X1 FILLER_61_1239 ();
 FILLCELL_X16 FILLER_62_1 ();
 FILLCELL_X4 FILLER_62_17 ();
 FILLCELL_X2 FILLER_62_24 ();
 FILLCELL_X1 FILLER_62_26 ();
 FILLCELL_X2 FILLER_62_80 ();
 FILLCELL_X1 FILLER_62_82 ();
 FILLCELL_X1 FILLER_62_111 ();
 FILLCELL_X1 FILLER_62_138 ();
 FILLCELL_X1 FILLER_62_203 ();
 FILLCELL_X4 FILLER_62_221 ();
 FILLCELL_X1 FILLER_62_225 ();
 FILLCELL_X2 FILLER_62_233 ();
 FILLCELL_X16 FILLER_62_248 ();
 FILLCELL_X8 FILLER_62_264 ();
 FILLCELL_X4 FILLER_62_272 ();
 FILLCELL_X2 FILLER_62_276 ();
 FILLCELL_X1 FILLER_62_278 ();
 FILLCELL_X2 FILLER_62_286 ();
 FILLCELL_X1 FILLER_62_288 ();
 FILLCELL_X8 FILLER_62_296 ();
 FILLCELL_X4 FILLER_62_304 ();
 FILLCELL_X2 FILLER_62_311 ();
 FILLCELL_X1 FILLER_62_313 ();
 FILLCELL_X1 FILLER_62_328 ();
 FILLCELL_X2 FILLER_62_336 ();
 FILLCELL_X4 FILLER_62_352 ();
 FILLCELL_X2 FILLER_62_356 ();
 FILLCELL_X4 FILLER_62_365 ();
 FILLCELL_X1 FILLER_62_376 ();
 FILLCELL_X2 FILLER_62_384 ();
 FILLCELL_X4 FILLER_62_403 ();
 FILLCELL_X2 FILLER_62_414 ();
 FILLCELL_X4 FILLER_62_433 ();
 FILLCELL_X8 FILLER_62_475 ();
 FILLCELL_X4 FILLER_62_483 ();
 FILLCELL_X1 FILLER_62_487 ();
 FILLCELL_X8 FILLER_62_506 ();
 FILLCELL_X8 FILLER_62_538 ();
 FILLCELL_X2 FILLER_62_546 ();
 FILLCELL_X1 FILLER_62_548 ();
 FILLCELL_X1 FILLER_62_565 ();
 FILLCELL_X8 FILLER_62_573 ();
 FILLCELL_X1 FILLER_62_581 ();
 FILLCELL_X4 FILLER_62_589 ();
 FILLCELL_X2 FILLER_62_593 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X8 FILLER_62_664 ();
 FILLCELL_X4 FILLER_62_672 ();
 FILLCELL_X8 FILLER_62_689 ();
 FILLCELL_X4 FILLER_62_697 ();
 FILLCELL_X2 FILLER_62_701 ();
 FILLCELL_X4 FILLER_62_727 ();
 FILLCELL_X2 FILLER_62_736 ();
 FILLCELL_X4 FILLER_62_755 ();
 FILLCELL_X8 FILLER_62_776 ();
 FILLCELL_X4 FILLER_62_784 ();
 FILLCELL_X2 FILLER_62_788 ();
 FILLCELL_X1 FILLER_62_790 ();
 FILLCELL_X1 FILLER_62_820 ();
 FILLCELL_X1 FILLER_62_826 ();
 FILLCELL_X2 FILLER_62_832 ();
 FILLCELL_X1 FILLER_62_839 ();
 FILLCELL_X1 FILLER_62_845 ();
 FILLCELL_X1 FILLER_62_855 ();
 FILLCELL_X2 FILLER_62_870 ();
 FILLCELL_X8 FILLER_62_886 ();
 FILLCELL_X2 FILLER_62_898 ();
 FILLCELL_X2 FILLER_62_905 ();
 FILLCELL_X1 FILLER_62_917 ();
 FILLCELL_X8 FILLER_62_934 ();
 FILLCELL_X4 FILLER_62_942 ();
 FILLCELL_X2 FILLER_62_946 ();
 FILLCELL_X1 FILLER_62_948 ();
 FILLCELL_X8 FILLER_62_952 ();
 FILLCELL_X4 FILLER_62_960 ();
 FILLCELL_X1 FILLER_62_964 ();
 FILLCELL_X1 FILLER_62_968 ();
 FILLCELL_X16 FILLER_62_989 ();
 FILLCELL_X2 FILLER_62_1005 ();
 FILLCELL_X1 FILLER_62_1007 ();
 FILLCELL_X32 FILLER_62_1013 ();
 FILLCELL_X32 FILLER_62_1045 ();
 FILLCELL_X16 FILLER_62_1077 ();
 FILLCELL_X4 FILLER_62_1093 ();
 FILLCELL_X1 FILLER_62_1097 ();
 FILLCELL_X2 FILLER_62_1105 ();
 FILLCELL_X32 FILLER_62_1131 ();
 FILLCELL_X8 FILLER_62_1163 ();
 FILLCELL_X1 FILLER_62_1171 ();
 FILLCELL_X4 FILLER_62_1189 ();
 FILLCELL_X16 FILLER_62_1196 ();
 FILLCELL_X4 FILLER_62_1212 ();
 FILLCELL_X2 FILLER_62_1229 ();
 FILLCELL_X2 FILLER_62_1237 ();
 FILLCELL_X1 FILLER_62_1239 ();
 FILLCELL_X16 FILLER_63_1 ();
 FILLCELL_X8 FILLER_63_17 ();
 FILLCELL_X4 FILLER_63_32 ();
 FILLCELL_X1 FILLER_63_36 ();
 FILLCELL_X4 FILLER_63_44 ();
 FILLCELL_X1 FILLER_63_48 ();
 FILLCELL_X16 FILLER_63_56 ();
 FILLCELL_X4 FILLER_63_72 ();
 FILLCELL_X2 FILLER_63_76 ();
 FILLCELL_X8 FILLER_63_85 ();
 FILLCELL_X1 FILLER_63_100 ();
 FILLCELL_X2 FILLER_63_108 ();
 FILLCELL_X4 FILLER_63_127 ();
 FILLCELL_X2 FILLER_63_138 ();
 FILLCELL_X4 FILLER_63_145 ();
 FILLCELL_X16 FILLER_63_154 ();
 FILLCELL_X8 FILLER_63_170 ();
 FILLCELL_X1 FILLER_63_178 ();
 FILLCELL_X4 FILLER_63_182 ();
 FILLCELL_X2 FILLER_63_186 ();
 FILLCELL_X1 FILLER_63_188 ();
 FILLCELL_X1 FILLER_63_199 ();
 FILLCELL_X8 FILLER_63_236 ();
 FILLCELL_X4 FILLER_63_251 ();
 FILLCELL_X2 FILLER_63_255 ();
 FILLCELL_X1 FILLER_63_257 ();
 FILLCELL_X2 FILLER_63_265 ();
 FILLCELL_X2 FILLER_63_284 ();
 FILLCELL_X1 FILLER_63_286 ();
 FILLCELL_X1 FILLER_63_294 ();
 FILLCELL_X2 FILLER_63_305 ();
 FILLCELL_X1 FILLER_63_345 ();
 FILLCELL_X1 FILLER_63_353 ();
 FILLCELL_X1 FILLER_63_361 ();
 FILLCELL_X1 FILLER_63_375 ();
 FILLCELL_X4 FILLER_63_393 ();
 FILLCELL_X2 FILLER_63_397 ();
 FILLCELL_X1 FILLER_63_399 ();
 FILLCELL_X4 FILLER_63_407 ();
 FILLCELL_X1 FILLER_63_411 ();
 FILLCELL_X2 FILLER_63_419 ();
 FILLCELL_X1 FILLER_63_421 ();
 FILLCELL_X2 FILLER_63_432 ();
 FILLCELL_X1 FILLER_63_434 ();
 FILLCELL_X2 FILLER_63_459 ();
 FILLCELL_X1 FILLER_63_461 ();
 FILLCELL_X32 FILLER_63_466 ();
 FILLCELL_X2 FILLER_63_498 ();
 FILLCELL_X1 FILLER_63_500 ();
 FILLCELL_X16 FILLER_63_532 ();
 FILLCELL_X2 FILLER_63_548 ();
 FILLCELL_X1 FILLER_63_550 ();
 FILLCELL_X4 FILLER_63_556 ();
 FILLCELL_X1 FILLER_63_560 ();
 FILLCELL_X8 FILLER_63_585 ();
 FILLCELL_X4 FILLER_63_600 ();
 FILLCELL_X2 FILLER_63_604 ();
 FILLCELL_X1 FILLER_63_606 ();
 FILLCELL_X32 FILLER_63_611 ();
 FILLCELL_X4 FILLER_63_643 ();
 FILLCELL_X2 FILLER_63_647 ();
 FILLCELL_X1 FILLER_63_649 ();
 FILLCELL_X4 FILLER_63_655 ();
 FILLCELL_X1 FILLER_63_659 ();
 FILLCELL_X2 FILLER_63_667 ();
 FILLCELL_X16 FILLER_63_686 ();
 FILLCELL_X4 FILLER_63_702 ();
 FILLCELL_X2 FILLER_63_720 ();
 FILLCELL_X1 FILLER_63_722 ();
 FILLCELL_X2 FILLER_63_750 ();
 FILLCELL_X1 FILLER_63_752 ();
 FILLCELL_X4 FILLER_63_784 ();
 FILLCELL_X2 FILLER_63_788 ();
 FILLCELL_X2 FILLER_63_812 ();
 FILLCELL_X1 FILLER_63_825 ();
 FILLCELL_X8 FILLER_63_831 ();
 FILLCELL_X4 FILLER_63_839 ();
 FILLCELL_X2 FILLER_63_843 ();
 FILLCELL_X8 FILLER_63_864 ();
 FILLCELL_X2 FILLER_63_872 ();
 FILLCELL_X4 FILLER_63_904 ();
 FILLCELL_X2 FILLER_63_908 ();
 FILLCELL_X16 FILLER_63_942 ();
 FILLCELL_X2 FILLER_63_958 ();
 FILLCELL_X1 FILLER_63_974 ();
 FILLCELL_X4 FILLER_63_978 ();
 FILLCELL_X4 FILLER_63_989 ();
 FILLCELL_X4 FILLER_63_996 ();
 FILLCELL_X2 FILLER_63_1000 ();
 FILLCELL_X4 FILLER_63_1033 ();
 FILLCELL_X1 FILLER_63_1037 ();
 FILLCELL_X4 FILLER_63_1047 ();
 FILLCELL_X2 FILLER_63_1051 ();
 FILLCELL_X1 FILLER_63_1053 ();
 FILLCELL_X16 FILLER_63_1075 ();
 FILLCELL_X4 FILLER_63_1091 ();
 FILLCELL_X2 FILLER_63_1095 ();
 FILLCELL_X8 FILLER_63_1104 ();
 FILLCELL_X4 FILLER_63_1112 ();
 FILLCELL_X2 FILLER_63_1116 ();
 FILLCELL_X1 FILLER_63_1118 ();
 FILLCELL_X2 FILLER_63_1143 ();
 FILLCELL_X1 FILLER_63_1145 ();
 FILLCELL_X4 FILLER_63_1163 ();
 FILLCELL_X1 FILLER_63_1167 ();
 FILLCELL_X8 FILLER_63_1192 ();
 FILLCELL_X2 FILLER_63_1200 ();
 FILLCELL_X1 FILLER_63_1202 ();
 FILLCELL_X1 FILLER_63_1213 ();
 FILLCELL_X2 FILLER_63_1238 ();
 FILLCELL_X16 FILLER_64_1 ();
 FILLCELL_X8 FILLER_64_17 ();
 FILLCELL_X1 FILLER_64_25 ();
 FILLCELL_X4 FILLER_64_43 ();
 FILLCELL_X1 FILLER_64_47 ();
 FILLCELL_X32 FILLER_64_53 ();
 FILLCELL_X8 FILLER_64_85 ();
 FILLCELL_X4 FILLER_64_93 ();
 FILLCELL_X1 FILLER_64_97 ();
 FILLCELL_X8 FILLER_64_103 ();
 FILLCELL_X4 FILLER_64_111 ();
 FILLCELL_X2 FILLER_64_115 ();
 FILLCELL_X1 FILLER_64_117 ();
 FILLCELL_X4 FILLER_64_123 ();
 FILLCELL_X1 FILLER_64_127 ();
 FILLCELL_X32 FILLER_64_145 ();
 FILLCELL_X32 FILLER_64_177 ();
 FILLCELL_X8 FILLER_64_209 ();
 FILLCELL_X4 FILLER_64_217 ();
 FILLCELL_X2 FILLER_64_221 ();
 FILLCELL_X8 FILLER_64_230 ();
 FILLCELL_X4 FILLER_64_238 ();
 FILLCELL_X2 FILLER_64_242 ();
 FILLCELL_X1 FILLER_64_244 ();
 FILLCELL_X4 FILLER_64_262 ();
 FILLCELL_X4 FILLER_64_307 ();
 FILLCELL_X2 FILLER_64_342 ();
 FILLCELL_X1 FILLER_64_365 ();
 FILLCELL_X16 FILLER_64_373 ();
 FILLCELL_X8 FILLER_64_389 ();
 FILLCELL_X4 FILLER_64_397 ();
 FILLCELL_X8 FILLER_64_418 ();
 FILLCELL_X2 FILLER_64_439 ();
 FILLCELL_X1 FILLER_64_471 ();
 FILLCELL_X16 FILLER_64_483 ();
 FILLCELL_X2 FILLER_64_499 ();
 FILLCELL_X32 FILLER_64_527 ();
 FILLCELL_X16 FILLER_64_559 ();
 FILLCELL_X4 FILLER_64_575 ();
 FILLCELL_X2 FILLER_64_579 ();
 FILLCELL_X1 FILLER_64_581 ();
 FILLCELL_X1 FILLER_64_630 ();
 FILLCELL_X16 FILLER_64_632 ();
 FILLCELL_X4 FILLER_64_648 ();
 FILLCELL_X2 FILLER_64_652 ();
 FILLCELL_X2 FILLER_64_699 ();
 FILLCELL_X1 FILLER_64_701 ();
 FILLCELL_X1 FILLER_64_726 ();
 FILLCELL_X1 FILLER_64_731 ();
 FILLCELL_X1 FILLER_64_739 ();
 FILLCELL_X2 FILLER_64_754 ();
 FILLCELL_X2 FILLER_64_763 ();
 FILLCELL_X1 FILLER_64_765 ();
 FILLCELL_X1 FILLER_64_770 ();
 FILLCELL_X2 FILLER_64_784 ();
 FILLCELL_X1 FILLER_64_786 ();
 FILLCELL_X1 FILLER_64_800 ();
 FILLCELL_X1 FILLER_64_805 ();
 FILLCELL_X32 FILLER_64_819 ();
 FILLCELL_X2 FILLER_64_851 ();
 FILLCELL_X1 FILLER_64_860 ();
 FILLCELL_X8 FILLER_64_866 ();
 FILLCELL_X2 FILLER_64_874 ();
 FILLCELL_X8 FILLER_64_886 ();
 FILLCELL_X2 FILLER_64_894 ();
 FILLCELL_X4 FILLER_64_901 ();
 FILLCELL_X1 FILLER_64_905 ();
 FILLCELL_X2 FILLER_64_930 ();
 FILLCELL_X16 FILLER_64_942 ();
 FILLCELL_X8 FILLER_64_958 ();
 FILLCELL_X8 FILLER_64_980 ();
 FILLCELL_X4 FILLER_64_988 ();
 FILLCELL_X2 FILLER_64_992 ();
 FILLCELL_X1 FILLER_64_994 ();
 FILLCELL_X2 FILLER_64_1005 ();
 FILLCELL_X1 FILLER_64_1007 ();
 FILLCELL_X1 FILLER_64_1022 ();
 FILLCELL_X1 FILLER_64_1040 ();
 FILLCELL_X1 FILLER_64_1058 ();
 FILLCELL_X8 FILLER_64_1072 ();
 FILLCELL_X4 FILLER_64_1080 ();
 FILLCELL_X2 FILLER_64_1084 ();
 FILLCELL_X8 FILLER_64_1103 ();
 FILLCELL_X4 FILLER_64_1111 ();
 FILLCELL_X2 FILLER_64_1115 ();
 FILLCELL_X1 FILLER_64_1117 ();
 FILLCELL_X1 FILLER_64_1135 ();
 FILLCELL_X1 FILLER_64_1160 ();
 FILLCELL_X2 FILLER_64_1174 ();
 FILLCELL_X1 FILLER_64_1183 ();
 FILLCELL_X1 FILLER_64_1191 ();
 FILLCELL_X1 FILLER_64_1209 ();
 FILLCELL_X2 FILLER_64_1217 ();
 FILLCELL_X1 FILLER_64_1236 ();
 FILLCELL_X16 FILLER_65_1 ();
 FILLCELL_X8 FILLER_65_17 ();
 FILLCELL_X16 FILLER_65_29 ();
 FILLCELL_X4 FILLER_65_45 ();
 FILLCELL_X2 FILLER_65_49 ();
 FILLCELL_X16 FILLER_65_56 ();
 FILLCELL_X8 FILLER_65_72 ();
 FILLCELL_X4 FILLER_65_104 ();
 FILLCELL_X8 FILLER_65_115 ();
 FILLCELL_X2 FILLER_65_123 ();
 FILLCELL_X2 FILLER_65_149 ();
 FILLCELL_X8 FILLER_65_163 ();
 FILLCELL_X1 FILLER_65_171 ();
 FILLCELL_X8 FILLER_65_179 ();
 FILLCELL_X2 FILLER_65_204 ();
 FILLCELL_X16 FILLER_65_223 ();
 FILLCELL_X4 FILLER_65_239 ();
 FILLCELL_X2 FILLER_65_243 ();
 FILLCELL_X2 FILLER_65_259 ();
 FILLCELL_X1 FILLER_65_261 ();
 FILLCELL_X4 FILLER_65_269 ();
 FILLCELL_X1 FILLER_65_280 ();
 FILLCELL_X16 FILLER_65_312 ();
 FILLCELL_X1 FILLER_65_335 ();
 FILLCELL_X32 FILLER_65_343 ();
 FILLCELL_X32 FILLER_65_375 ();
 FILLCELL_X16 FILLER_65_407 ();
 FILLCELL_X8 FILLER_65_423 ();
 FILLCELL_X4 FILLER_65_431 ();
 FILLCELL_X1 FILLER_65_435 ();
 FILLCELL_X16 FILLER_65_440 ();
 FILLCELL_X8 FILLER_65_456 ();
 FILLCELL_X4 FILLER_65_464 ();
 FILLCELL_X1 FILLER_65_468 ();
 FILLCELL_X2 FILLER_65_500 ();
 FILLCELL_X1 FILLER_65_509 ();
 FILLCELL_X1 FILLER_65_525 ();
 FILLCELL_X8 FILLER_65_538 ();
 FILLCELL_X2 FILLER_65_546 ();
 FILLCELL_X1 FILLER_65_548 ();
 FILLCELL_X1 FILLER_65_566 ();
 FILLCELL_X1 FILLER_65_591 ();
 FILLCELL_X1 FILLER_65_630 ();
 FILLCELL_X8 FILLER_65_648 ();
 FILLCELL_X2 FILLER_65_694 ();
 FILLCELL_X1 FILLER_65_696 ();
 FILLCELL_X32 FILLER_65_710 ();
 FILLCELL_X32 FILLER_65_742 ();
 FILLCELL_X16 FILLER_65_774 ();
 FILLCELL_X2 FILLER_65_790 ();
 FILLCELL_X2 FILLER_65_795 ();
 FILLCELL_X1 FILLER_65_797 ();
 FILLCELL_X2 FILLER_65_802 ();
 FILLCELL_X2 FILLER_65_819 ();
 FILLCELL_X1 FILLER_65_821 ();
 FILLCELL_X1 FILLER_65_827 ();
 FILLCELL_X2 FILLER_65_836 ();
 FILLCELL_X32 FILLER_65_843 ();
 FILLCELL_X1 FILLER_65_875 ();
 FILLCELL_X2 FILLER_65_904 ();
 FILLCELL_X1 FILLER_65_906 ();
 FILLCELL_X4 FILLER_65_926 ();
 FILLCELL_X1 FILLER_65_930 ();
 FILLCELL_X16 FILLER_65_938 ();
 FILLCELL_X2 FILLER_65_954 ();
 FILLCELL_X8 FILLER_65_961 ();
 FILLCELL_X2 FILLER_65_969 ();
 FILLCELL_X1 FILLER_65_971 ();
 FILLCELL_X8 FILLER_65_982 ();
 FILLCELL_X1 FILLER_65_990 ();
 FILLCELL_X1 FILLER_65_1015 ();
 FILLCELL_X1 FILLER_65_1050 ();
 FILLCELL_X1 FILLER_65_1058 ();
 FILLCELL_X2 FILLER_65_1064 ();
 FILLCELL_X1 FILLER_65_1066 ();
 FILLCELL_X8 FILLER_65_1074 ();
 FILLCELL_X1 FILLER_65_1082 ();
 FILLCELL_X8 FILLER_65_1114 ();
 FILLCELL_X4 FILLER_65_1129 ();
 FILLCELL_X2 FILLER_65_1133 ();
 FILLCELL_X1 FILLER_65_1135 ();
 FILLCELL_X4 FILLER_65_1143 ();
 FILLCELL_X1 FILLER_65_1147 ();
 FILLCELL_X1 FILLER_65_1169 ();
 FILLCELL_X4 FILLER_65_1174 ();
 FILLCELL_X2 FILLER_65_1178 ();
 FILLCELL_X1 FILLER_65_1180 ();
 FILLCELL_X2 FILLER_65_1235 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X8 FILLER_66_33 ();
 FILLCELL_X4 FILLER_66_41 ();
 FILLCELL_X32 FILLER_66_62 ();
 FILLCELL_X8 FILLER_66_122 ();
 FILLCELL_X2 FILLER_66_130 ();
 FILLCELL_X2 FILLER_66_149 ();
 FILLCELL_X1 FILLER_66_151 ();
 FILLCELL_X2 FILLER_66_193 ();
 FILLCELL_X1 FILLER_66_195 ();
 FILLCELL_X2 FILLER_66_210 ();
 FILLCELL_X1 FILLER_66_212 ();
 FILLCELL_X16 FILLER_66_220 ();
 FILLCELL_X4 FILLER_66_236 ();
 FILLCELL_X2 FILLER_66_240 ();
 FILLCELL_X1 FILLER_66_250 ();
 FILLCELL_X32 FILLER_66_268 ();
 FILLCELL_X16 FILLER_66_300 ();
 FILLCELL_X1 FILLER_66_316 ();
 FILLCELL_X2 FILLER_66_324 ();
 FILLCELL_X1 FILLER_66_326 ();
 FILLCELL_X2 FILLER_66_341 ();
 FILLCELL_X2 FILLER_66_350 ();
 FILLCELL_X1 FILLER_66_352 ();
 FILLCELL_X4 FILLER_66_377 ();
 FILLCELL_X1 FILLER_66_381 ();
 FILLCELL_X32 FILLER_66_387 ();
 FILLCELL_X2 FILLER_66_419 ();
 FILLCELL_X1 FILLER_66_421 ();
 FILLCELL_X4 FILLER_66_439 ();
 FILLCELL_X2 FILLER_66_443 ();
 FILLCELL_X1 FILLER_66_445 ();
 FILLCELL_X8 FILLER_66_463 ();
 FILLCELL_X4 FILLER_66_471 ();
 FILLCELL_X2 FILLER_66_475 ();
 FILLCELL_X8 FILLER_66_484 ();
 FILLCELL_X4 FILLER_66_492 ();
 FILLCELL_X1 FILLER_66_496 ();
 FILLCELL_X2 FILLER_66_514 ();
 FILLCELL_X1 FILLER_66_516 ();
 FILLCELL_X2 FILLER_66_530 ();
 FILLCELL_X8 FILLER_66_570 ();
 FILLCELL_X4 FILLER_66_578 ();
 FILLCELL_X4 FILLER_66_589 ();
 FILLCELL_X2 FILLER_66_593 ();
 FILLCELL_X4 FILLER_66_609 ();
 FILLCELL_X2 FILLER_66_613 ();
 FILLCELL_X1 FILLER_66_615 ();
 FILLCELL_X1 FILLER_66_623 ();
 FILLCELL_X2 FILLER_66_632 ();
 FILLCELL_X16 FILLER_66_651 ();
 FILLCELL_X2 FILLER_66_667 ();
 FILLCELL_X1 FILLER_66_669 ();
 FILLCELL_X1 FILLER_66_694 ();
 FILLCELL_X8 FILLER_66_699 ();
 FILLCELL_X2 FILLER_66_707 ();
 FILLCELL_X1 FILLER_66_709 ();
 FILLCELL_X2 FILLER_66_727 ();
 FILLCELL_X1 FILLER_66_729 ();
 FILLCELL_X32 FILLER_66_743 ();
 FILLCELL_X16 FILLER_66_775 ();
 FILLCELL_X2 FILLER_66_791 ();
 FILLCELL_X2 FILLER_66_800 ();
 FILLCELL_X2 FILLER_66_807 ();
 FILLCELL_X1 FILLER_66_816 ();
 FILLCELL_X1 FILLER_66_826 ();
 FILLCELL_X16 FILLER_66_841 ();
 FILLCELL_X16 FILLER_66_867 ();
 FILLCELL_X1 FILLER_66_883 ();
 FILLCELL_X32 FILLER_66_893 ();
 FILLCELL_X32 FILLER_66_925 ();
 FILLCELL_X4 FILLER_66_957 ();
 FILLCELL_X2 FILLER_66_961 ();
 FILLCELL_X1 FILLER_66_963 ();
 FILLCELL_X2 FILLER_66_991 ();
 FILLCELL_X8 FILLER_66_996 ();
 FILLCELL_X8 FILLER_66_1024 ();
 FILLCELL_X2 FILLER_66_1040 ();
 FILLCELL_X4 FILLER_66_1083 ();
 FILLCELL_X8 FILLER_66_1108 ();
 FILLCELL_X4 FILLER_66_1116 ();
 FILLCELL_X1 FILLER_66_1120 ();
 FILLCELL_X16 FILLER_66_1135 ();
 FILLCELL_X8 FILLER_66_1151 ();
 FILLCELL_X1 FILLER_66_1159 ();
 FILLCELL_X16 FILLER_66_1177 ();
 FILLCELL_X8 FILLER_66_1193 ();
 FILLCELL_X2 FILLER_66_1201 ();
 FILLCELL_X1 FILLER_66_1203 ();
 FILLCELL_X1 FILLER_66_1207 ();
 FILLCELL_X1 FILLER_66_1219 ();
 FILLCELL_X2 FILLER_66_1237 ();
 FILLCELL_X1 FILLER_66_1239 ();
 FILLCELL_X8 FILLER_67_1 ();
 FILLCELL_X16 FILLER_67_12 ();
 FILLCELL_X8 FILLER_67_28 ();
 FILLCELL_X4 FILLER_67_36 ();
 FILLCELL_X1 FILLER_67_40 ();
 FILLCELL_X8 FILLER_67_75 ();
 FILLCELL_X4 FILLER_67_83 ();
 FILLCELL_X4 FILLER_67_94 ();
 FILLCELL_X1 FILLER_67_98 ();
 FILLCELL_X4 FILLER_67_106 ();
 FILLCELL_X1 FILLER_67_110 ();
 FILLCELL_X8 FILLER_67_125 ();
 FILLCELL_X4 FILLER_67_133 ();
 FILLCELL_X2 FILLER_67_144 ();
 FILLCELL_X1 FILLER_67_146 ();
 FILLCELL_X8 FILLER_67_154 ();
 FILLCELL_X4 FILLER_67_162 ();
 FILLCELL_X2 FILLER_67_166 ();
 FILLCELL_X16 FILLER_67_173 ();
 FILLCELL_X8 FILLER_67_189 ();
 FILLCELL_X2 FILLER_67_197 ();
 FILLCELL_X1 FILLER_67_199 ();
 FILLCELL_X16 FILLER_67_207 ();
 FILLCELL_X2 FILLER_67_223 ();
 FILLCELL_X1 FILLER_67_225 ();
 FILLCELL_X16 FILLER_67_257 ();
 FILLCELL_X8 FILLER_67_273 ();
 FILLCELL_X2 FILLER_67_281 ();
 FILLCELL_X1 FILLER_67_283 ();
 FILLCELL_X16 FILLER_67_289 ();
 FILLCELL_X4 FILLER_67_305 ();
 FILLCELL_X1 FILLER_67_309 ();
 FILLCELL_X2 FILLER_67_334 ();
 FILLCELL_X4 FILLER_67_344 ();
 FILLCELL_X1 FILLER_67_348 ();
 FILLCELL_X4 FILLER_67_373 ();
 FILLCELL_X1 FILLER_67_377 ();
 FILLCELL_X4 FILLER_67_419 ();
 FILLCELL_X2 FILLER_67_423 ();
 FILLCELL_X2 FILLER_67_473 ();
 FILLCELL_X1 FILLER_67_475 ();
 FILLCELL_X16 FILLER_67_493 ();
 FILLCELL_X2 FILLER_67_509 ();
 FILLCELL_X2 FILLER_67_518 ();
 FILLCELL_X4 FILLER_67_523 ();
 FILLCELL_X16 FILLER_67_534 ();
 FILLCELL_X4 FILLER_67_550 ();
 FILLCELL_X1 FILLER_67_554 ();
 FILLCELL_X8 FILLER_67_572 ();
 FILLCELL_X2 FILLER_67_580 ();
 FILLCELL_X1 FILLER_67_582 ();
 FILLCELL_X4 FILLER_67_600 ();
 FILLCELL_X2 FILLER_67_604 ();
 FILLCELL_X32 FILLER_67_644 ();
 FILLCELL_X8 FILLER_67_676 ();
 FILLCELL_X4 FILLER_67_684 ();
 FILLCELL_X2 FILLER_67_688 ();
 FILLCELL_X8 FILLER_67_702 ();
 FILLCELL_X4 FILLER_67_710 ();
 FILLCELL_X8 FILLER_67_745 ();
 FILLCELL_X2 FILLER_67_753 ();
 FILLCELL_X4 FILLER_67_796 ();
 FILLCELL_X2 FILLER_67_800 ();
 FILLCELL_X1 FILLER_67_802 ();
 FILLCELL_X8 FILLER_67_808 ();
 FILLCELL_X2 FILLER_67_816 ();
 FILLCELL_X1 FILLER_67_821 ();
 FILLCELL_X1 FILLER_67_841 ();
 FILLCELL_X4 FILLER_67_847 ();
 FILLCELL_X2 FILLER_67_851 ();
 FILLCELL_X2 FILLER_67_877 ();
 FILLCELL_X4 FILLER_67_893 ();
 FILLCELL_X4 FILLER_67_902 ();
 FILLCELL_X1 FILLER_67_906 ();
 FILLCELL_X2 FILLER_67_916 ();
 FILLCELL_X1 FILLER_67_918 ();
 FILLCELL_X2 FILLER_67_922 ();
 FILLCELL_X1 FILLER_67_929 ();
 FILLCELL_X1 FILLER_67_933 ();
 FILLCELL_X1 FILLER_67_956 ();
 FILLCELL_X4 FILLER_67_962 ();
 FILLCELL_X2 FILLER_67_966 ();
 FILLCELL_X1 FILLER_67_968 ();
 FILLCELL_X1 FILLER_67_978 ();
 FILLCELL_X16 FILLER_67_987 ();
 FILLCELL_X8 FILLER_67_1003 ();
 FILLCELL_X2 FILLER_67_1011 ();
 FILLCELL_X1 FILLER_67_1013 ();
 FILLCELL_X32 FILLER_67_1021 ();
 FILLCELL_X16 FILLER_67_1053 ();
 FILLCELL_X8 FILLER_67_1069 ();
 FILLCELL_X4 FILLER_67_1077 ();
 FILLCELL_X2 FILLER_67_1081 ();
 FILLCELL_X1 FILLER_67_1083 ();
 FILLCELL_X8 FILLER_67_1110 ();
 FILLCELL_X4 FILLER_67_1118 ();
 FILLCELL_X8 FILLER_67_1139 ();
 FILLCELL_X2 FILLER_67_1147 ();
 FILLCELL_X1 FILLER_67_1166 ();
 FILLCELL_X8 FILLER_67_1184 ();
 FILLCELL_X2 FILLER_67_1192 ();
 FILLCELL_X1 FILLER_67_1234 ();
 FILLCELL_X2 FILLER_67_1238 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X2 FILLER_68_33 ();
 FILLCELL_X4 FILLER_68_39 ();
 FILLCELL_X8 FILLER_68_67 ();
 FILLCELL_X1 FILLER_68_75 ();
 FILLCELL_X8 FILLER_68_100 ();
 FILLCELL_X4 FILLER_68_108 ();
 FILLCELL_X16 FILLER_68_129 ();
 FILLCELL_X4 FILLER_68_145 ();
 FILLCELL_X2 FILLER_68_149 ();
 FILLCELL_X8 FILLER_68_196 ();
 FILLCELL_X2 FILLER_68_204 ();
 FILLCELL_X2 FILLER_68_229 ();
 FILLCELL_X1 FILLER_68_231 ();
 FILLCELL_X8 FILLER_68_263 ();
 FILLCELL_X1 FILLER_68_271 ();
 FILLCELL_X2 FILLER_68_279 ();
 FILLCELL_X1 FILLER_68_281 ();
 FILLCELL_X1 FILLER_68_289 ();
 FILLCELL_X4 FILLER_68_338 ();
 FILLCELL_X1 FILLER_68_342 ();
 FILLCELL_X4 FILLER_68_346 ();
 FILLCELL_X2 FILLER_68_350 ();
 FILLCELL_X2 FILLER_68_359 ();
 FILLCELL_X1 FILLER_68_361 ();
 FILLCELL_X2 FILLER_68_379 ();
 FILLCELL_X1 FILLER_68_381 ();
 FILLCELL_X2 FILLER_68_389 ();
 FILLCELL_X1 FILLER_68_391 ();
 FILLCELL_X2 FILLER_68_409 ();
 FILLCELL_X1 FILLER_68_418 ();
 FILLCELL_X2 FILLER_68_433 ();
 FILLCELL_X1 FILLER_68_435 ();
 FILLCELL_X4 FILLER_68_443 ();
 FILLCELL_X1 FILLER_68_447 ();
 FILLCELL_X2 FILLER_68_455 ();
 FILLCELL_X1 FILLER_68_461 ();
 FILLCELL_X1 FILLER_68_478 ();
 FILLCELL_X16 FILLER_68_486 ();
 FILLCELL_X8 FILLER_68_502 ();
 FILLCELL_X4 FILLER_68_534 ();
 FILLCELL_X2 FILLER_68_538 ();
 FILLCELL_X32 FILLER_68_547 ();
 FILLCELL_X16 FILLER_68_579 ();
 FILLCELL_X8 FILLER_68_595 ();
 FILLCELL_X8 FILLER_68_620 ();
 FILLCELL_X2 FILLER_68_628 ();
 FILLCELL_X1 FILLER_68_630 ();
 FILLCELL_X16 FILLER_68_632 ();
 FILLCELL_X2 FILLER_68_648 ();
 FILLCELL_X16 FILLER_68_658 ();
 FILLCELL_X4 FILLER_68_674 ();
 FILLCELL_X1 FILLER_68_685 ();
 FILLCELL_X2 FILLER_68_703 ();
 FILLCELL_X2 FILLER_68_722 ();
 FILLCELL_X2 FILLER_68_741 ();
 FILLCELL_X1 FILLER_68_743 ();
 FILLCELL_X1 FILLER_68_748 ();
 FILLCELL_X8 FILLER_68_756 ();
 FILLCELL_X1 FILLER_68_764 ();
 FILLCELL_X16 FILLER_68_803 ();
 FILLCELL_X4 FILLER_68_819 ();
 FILLCELL_X4 FILLER_68_830 ();
 FILLCELL_X1 FILLER_68_834 ();
 FILLCELL_X8 FILLER_68_838 ();
 FILLCELL_X4 FILLER_68_846 ();
 FILLCELL_X2 FILLER_68_850 ();
 FILLCELL_X2 FILLER_68_859 ();
 FILLCELL_X2 FILLER_68_877 ();
 FILLCELL_X2 FILLER_68_891 ();
 FILLCELL_X2 FILLER_68_915 ();
 FILLCELL_X1 FILLER_68_933 ();
 FILLCELL_X2 FILLER_68_944 ();
 FILLCELL_X2 FILLER_68_951 ();
 FILLCELL_X32 FILLER_68_962 ();
 FILLCELL_X4 FILLER_68_994 ();
 FILLCELL_X2 FILLER_68_998 ();
 FILLCELL_X1 FILLER_68_1000 ();
 FILLCELL_X16 FILLER_68_1025 ();
 FILLCELL_X4 FILLER_68_1041 ();
 FILLCELL_X1 FILLER_68_1045 ();
 FILLCELL_X8 FILLER_68_1060 ();
 FILLCELL_X4 FILLER_68_1068 ();
 FILLCELL_X1 FILLER_68_1072 ();
 FILLCELL_X8 FILLER_68_1078 ();
 FILLCELL_X2 FILLER_68_1086 ();
 FILLCELL_X1 FILLER_68_1088 ();
 FILLCELL_X4 FILLER_68_1111 ();
 FILLCELL_X2 FILLER_68_1115 ();
 FILLCELL_X8 FILLER_68_1141 ();
 FILLCELL_X2 FILLER_68_1149 ();
 FILLCELL_X1 FILLER_68_1151 ();
 FILLCELL_X2 FILLER_68_1159 ();
 FILLCELL_X8 FILLER_68_1185 ();
 FILLCELL_X2 FILLER_68_1193 ();
 FILLCELL_X1 FILLER_68_1195 ();
 FILLCELL_X2 FILLER_68_1217 ();
 FILLCELL_X1 FILLER_68_1219 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_33 ();
 FILLCELL_X2 FILLER_69_37 ();
 FILLCELL_X4 FILLER_69_46 ();
 FILLCELL_X1 FILLER_69_50 ();
 FILLCELL_X4 FILLER_69_58 ();
 FILLCELL_X1 FILLER_69_62 ();
 FILLCELL_X8 FILLER_69_70 ();
 FILLCELL_X4 FILLER_69_78 ();
 FILLCELL_X2 FILLER_69_82 ();
 FILLCELL_X32 FILLER_69_91 ();
 FILLCELL_X8 FILLER_69_123 ();
 FILLCELL_X4 FILLER_69_131 ();
 FILLCELL_X4 FILLER_69_142 ();
 FILLCELL_X8 FILLER_69_153 ();
 FILLCELL_X4 FILLER_69_161 ();
 FILLCELL_X2 FILLER_69_165 ();
 FILLCELL_X1 FILLER_69_167 ();
 FILLCELL_X8 FILLER_69_170 ();
 FILLCELL_X2 FILLER_69_178 ();
 FILLCELL_X1 FILLER_69_197 ();
 FILLCELL_X2 FILLER_69_201 ();
 FILLCELL_X1 FILLER_69_203 ();
 FILLCELL_X32 FILLER_69_211 ();
 FILLCELL_X4 FILLER_69_243 ();
 FILLCELL_X1 FILLER_69_247 ();
 FILLCELL_X4 FILLER_69_269 ();
 FILLCELL_X1 FILLER_69_273 ();
 FILLCELL_X16 FILLER_69_291 ();
 FILLCELL_X8 FILLER_69_307 ();
 FILLCELL_X1 FILLER_69_315 ();
 FILLCELL_X2 FILLER_69_340 ();
 FILLCELL_X4 FILLER_69_349 ();
 FILLCELL_X1 FILLER_69_353 ();
 FILLCELL_X2 FILLER_69_406 ();
 FILLCELL_X1 FILLER_69_408 ();
 FILLCELL_X32 FILLER_69_416 ();
 FILLCELL_X8 FILLER_69_448 ();
 FILLCELL_X4 FILLER_69_456 ();
 FILLCELL_X1 FILLER_69_460 ();
 FILLCELL_X8 FILLER_69_472 ();
 FILLCELL_X32 FILLER_69_485 ();
 FILLCELL_X16 FILLER_69_517 ();
 FILLCELL_X8 FILLER_69_533 ();
 FILLCELL_X2 FILLER_69_541 ();
 FILLCELL_X1 FILLER_69_543 ();
 FILLCELL_X16 FILLER_69_547 ();
 FILLCELL_X1 FILLER_69_563 ();
 FILLCELL_X2 FILLER_69_611 ();
 FILLCELL_X1 FILLER_69_613 ();
 FILLCELL_X16 FILLER_69_631 ();
 FILLCELL_X8 FILLER_69_647 ();
 FILLCELL_X2 FILLER_69_655 ();
 FILLCELL_X8 FILLER_69_674 ();
 FILLCELL_X1 FILLER_69_682 ();
 FILLCELL_X4 FILLER_69_707 ();
 FILLCELL_X2 FILLER_69_711 ();
 FILLCELL_X1 FILLER_69_713 ();
 FILLCELL_X4 FILLER_69_735 ();
 FILLCELL_X2 FILLER_69_739 ();
 FILLCELL_X1 FILLER_69_741 ();
 FILLCELL_X4 FILLER_69_749 ();
 FILLCELL_X2 FILLER_69_753 ();
 FILLCELL_X8 FILLER_69_799 ();
 FILLCELL_X4 FILLER_69_807 ();
 FILLCELL_X16 FILLER_69_816 ();
 FILLCELL_X8 FILLER_69_832 ();
 FILLCELL_X2 FILLER_69_840 ();
 FILLCELL_X1 FILLER_69_842 ();
 FILLCELL_X2 FILLER_69_853 ();
 FILLCELL_X1 FILLER_69_855 ();
 FILLCELL_X1 FILLER_69_861 ();
 FILLCELL_X1 FILLER_69_865 ();
 FILLCELL_X2 FILLER_69_869 ();
 FILLCELL_X1 FILLER_69_875 ();
 FILLCELL_X4 FILLER_69_881 ();
 FILLCELL_X2 FILLER_69_889 ();
 FILLCELL_X16 FILLER_69_896 ();
 FILLCELL_X4 FILLER_69_912 ();
 FILLCELL_X4 FILLER_69_928 ();
 FILLCELL_X2 FILLER_69_946 ();
 FILLCELL_X1 FILLER_69_948 ();
 FILLCELL_X8 FILLER_69_952 ();
 FILLCELL_X2 FILLER_69_960 ();
 FILLCELL_X4 FILLER_69_965 ();
 FILLCELL_X1 FILLER_69_972 ();
 FILLCELL_X2 FILLER_69_982 ();
 FILLCELL_X1 FILLER_69_984 ();
 FILLCELL_X4 FILLER_69_988 ();
 FILLCELL_X2 FILLER_69_992 ();
 FILLCELL_X1 FILLER_69_994 ();
 FILLCELL_X1 FILLER_69_1036 ();
 FILLCELL_X1 FILLER_69_1054 ();
 FILLCELL_X1 FILLER_69_1062 ();
 FILLCELL_X2 FILLER_69_1070 ();
 FILLCELL_X2 FILLER_69_1096 ();
 FILLCELL_X1 FILLER_69_1098 ();
 FILLCELL_X32 FILLER_69_1102 ();
 FILLCELL_X2 FILLER_69_1134 ();
 FILLCELL_X16 FILLER_69_1181 ();
 FILLCELL_X1 FILLER_69_1197 ();
 FILLCELL_X1 FILLER_69_1222 ();
 FILLCELL_X4 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_9 ();
 FILLCELL_X8 FILLER_70_41 ();
 FILLCELL_X1 FILLER_70_49 ();
 FILLCELL_X8 FILLER_70_67 ();
 FILLCELL_X2 FILLER_70_75 ();
 FILLCELL_X1 FILLER_70_77 ();
 FILLCELL_X4 FILLER_70_95 ();
 FILLCELL_X2 FILLER_70_99 ();
 FILLCELL_X2 FILLER_70_125 ();
 FILLCELL_X2 FILLER_70_151 ();
 FILLCELL_X2 FILLER_70_167 ();
 FILLCELL_X2 FILLER_70_223 ();
 FILLCELL_X1 FILLER_70_225 ();
 FILLCELL_X4 FILLER_70_233 ();
 FILLCELL_X2 FILLER_70_237 ();
 FILLCELL_X4 FILLER_70_256 ();
 FILLCELL_X2 FILLER_70_260 ();
 FILLCELL_X4 FILLER_70_279 ();
 FILLCELL_X16 FILLER_70_290 ();
 FILLCELL_X4 FILLER_70_306 ();
 FILLCELL_X2 FILLER_70_310 ();
 FILLCELL_X1 FILLER_70_312 ();
 FILLCELL_X4 FILLER_70_320 ();
 FILLCELL_X8 FILLER_70_334 ();
 FILLCELL_X1 FILLER_70_342 ();
 FILLCELL_X4 FILLER_70_356 ();
 FILLCELL_X2 FILLER_70_360 ();
 FILLCELL_X1 FILLER_70_362 ();
 FILLCELL_X1 FILLER_70_380 ();
 FILLCELL_X16 FILLER_70_386 ();
 FILLCELL_X8 FILLER_70_402 ();
 FILLCELL_X4 FILLER_70_410 ();
 FILLCELL_X2 FILLER_70_414 ();
 FILLCELL_X1 FILLER_70_416 ();
 FILLCELL_X32 FILLER_70_421 ();
 FILLCELL_X4 FILLER_70_453 ();
 FILLCELL_X8 FILLER_70_508 ();
 FILLCELL_X4 FILLER_70_516 ();
 FILLCELL_X1 FILLER_70_520 ();
 FILLCELL_X1 FILLER_70_528 ();
 FILLCELL_X8 FILLER_70_536 ();
 FILLCELL_X4 FILLER_70_544 ();
 FILLCELL_X2 FILLER_70_548 ();
 FILLCELL_X8 FILLER_70_557 ();
 FILLCELL_X4 FILLER_70_565 ();
 FILLCELL_X8 FILLER_70_620 ();
 FILLCELL_X2 FILLER_70_628 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X16 FILLER_70_632 ();
 FILLCELL_X8 FILLER_70_648 ();
 FILLCELL_X1 FILLER_70_680 ();
 FILLCELL_X4 FILLER_70_688 ();
 FILLCELL_X2 FILLER_70_692 ();
 FILLCELL_X4 FILLER_70_701 ();
 FILLCELL_X2 FILLER_70_705 ();
 FILLCELL_X1 FILLER_70_707 ();
 FILLCELL_X32 FILLER_70_715 ();
 FILLCELL_X2 FILLER_70_747 ();
 FILLCELL_X1 FILLER_70_749 ();
 FILLCELL_X8 FILLER_70_757 ();
 FILLCELL_X4 FILLER_70_765 ();
 FILLCELL_X2 FILLER_70_769 ();
 FILLCELL_X1 FILLER_70_771 ();
 FILLCELL_X2 FILLER_70_776 ();
 FILLCELL_X8 FILLER_70_785 ();
 FILLCELL_X2 FILLER_70_793 ();
 FILLCELL_X1 FILLER_70_795 ();
 FILLCELL_X1 FILLER_70_801 ();
 FILLCELL_X2 FILLER_70_807 ();
 FILLCELL_X1 FILLER_70_809 ();
 FILLCELL_X1 FILLER_70_818 ();
 FILLCELL_X2 FILLER_70_828 ();
 FILLCELL_X1 FILLER_70_830 ();
 FILLCELL_X2 FILLER_70_839 ();
 FILLCELL_X16 FILLER_70_845 ();
 FILLCELL_X8 FILLER_70_861 ();
 FILLCELL_X4 FILLER_70_869 ();
 FILLCELL_X2 FILLER_70_873 ();
 FILLCELL_X1 FILLER_70_875 ();
 FILLCELL_X8 FILLER_70_881 ();
 FILLCELL_X2 FILLER_70_889 ();
 FILLCELL_X1 FILLER_70_891 ();
 FILLCELL_X2 FILLER_70_895 ();
 FILLCELL_X4 FILLER_70_902 ();
 FILLCELL_X2 FILLER_70_906 ();
 FILLCELL_X32 FILLER_70_911 ();
 FILLCELL_X16 FILLER_70_943 ();
 FILLCELL_X8 FILLER_70_991 ();
 FILLCELL_X4 FILLER_70_999 ();
 FILLCELL_X4 FILLER_70_1036 ();
 FILLCELL_X32 FILLER_70_1084 ();
 FILLCELL_X16 FILLER_70_1116 ();
 FILLCELL_X4 FILLER_70_1132 ();
 FILLCELL_X1 FILLER_70_1136 ();
 FILLCELL_X8 FILLER_70_1154 ();
 FILLCELL_X1 FILLER_70_1162 ();
 FILLCELL_X8 FILLER_70_1168 ();
 FILLCELL_X1 FILLER_70_1176 ();
 FILLCELL_X4 FILLER_70_1184 ();
 FILLCELL_X2 FILLER_70_1188 ();
 FILLCELL_X1 FILLER_70_1190 ();
 FILLCELL_X2 FILLER_70_1198 ();
 FILLCELL_X1 FILLER_70_1200 ();
 FILLCELL_X4 FILLER_70_1204 ();
 FILLCELL_X1 FILLER_70_1208 ();
 FILLCELL_X4 FILLER_70_1212 ();
 FILLCELL_X4 FILLER_70_1219 ();
 FILLCELL_X1 FILLER_70_1223 ();
 FILLCELL_X4 FILLER_70_1230 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X16 FILLER_71_33 ();
 FILLCELL_X4 FILLER_71_49 ();
 FILLCELL_X2 FILLER_71_53 ();
 FILLCELL_X1 FILLER_71_55 ();
 FILLCELL_X8 FILLER_71_73 ();
 FILLCELL_X2 FILLER_71_81 ();
 FILLCELL_X2 FILLER_71_107 ();
 FILLCELL_X1 FILLER_71_109 ();
 FILLCELL_X2 FILLER_71_117 ();
 FILLCELL_X4 FILLER_71_141 ();
 FILLCELL_X1 FILLER_71_145 ();
 FILLCELL_X16 FILLER_71_153 ();
 FILLCELL_X2 FILLER_71_169 ();
 FILLCELL_X2 FILLER_71_178 ();
 FILLCELL_X1 FILLER_71_180 ();
 FILLCELL_X2 FILLER_71_188 ();
 FILLCELL_X1 FILLER_71_190 ();
 FILLCELL_X4 FILLER_71_194 ();
 FILLCELL_X2 FILLER_71_211 ();
 FILLCELL_X16 FILLER_71_237 ();
 FILLCELL_X4 FILLER_71_281 ();
 FILLCELL_X2 FILLER_71_285 ();
 FILLCELL_X16 FILLER_71_294 ();
 FILLCELL_X8 FILLER_71_313 ();
 FILLCELL_X2 FILLER_71_321 ();
 FILLCELL_X1 FILLER_71_323 ();
 FILLCELL_X8 FILLER_71_331 ();
 FILLCELL_X4 FILLER_71_339 ();
 FILLCELL_X2 FILLER_71_343 ();
 FILLCELL_X1 FILLER_71_345 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X4 FILLER_71_385 ();
 FILLCELL_X8 FILLER_71_396 ();
 FILLCELL_X4 FILLER_71_404 ();
 FILLCELL_X2 FILLER_71_408 ();
 FILLCELL_X4 FILLER_71_465 ();
 FILLCELL_X1 FILLER_71_469 ();
 FILLCELL_X8 FILLER_71_474 ();
 FILLCELL_X1 FILLER_71_482 ();
 FILLCELL_X1 FILLER_71_490 ();
 FILLCELL_X2 FILLER_71_508 ();
 FILLCELL_X1 FILLER_71_527 ();
 FILLCELL_X2 FILLER_71_545 ();
 FILLCELL_X16 FILLER_71_564 ();
 FILLCELL_X4 FILLER_71_580 ();
 FILLCELL_X2 FILLER_71_584 ();
 FILLCELL_X1 FILLER_71_612 ();
 FILLCELL_X16 FILLER_71_630 ();
 FILLCELL_X8 FILLER_71_646 ();
 FILLCELL_X4 FILLER_71_654 ();
 FILLCELL_X2 FILLER_71_658 ();
 FILLCELL_X4 FILLER_71_667 ();
 FILLCELL_X4 FILLER_71_708 ();
 FILLCELL_X1 FILLER_71_712 ();
 FILLCELL_X8 FILLER_71_724 ();
 FILLCELL_X1 FILLER_71_732 ();
 FILLCELL_X8 FILLER_71_740 ();
 FILLCELL_X4 FILLER_71_748 ();
 FILLCELL_X1 FILLER_71_752 ();
 FILLCELL_X2 FILLER_71_763 ();
 FILLCELL_X1 FILLER_71_775 ();
 FILLCELL_X8 FILLER_71_783 ();
 FILLCELL_X4 FILLER_71_791 ();
 FILLCELL_X2 FILLER_71_795 ();
 FILLCELL_X1 FILLER_71_797 ();
 FILLCELL_X2 FILLER_71_826 ();
 FILLCELL_X4 FILLER_71_833 ();
 FILLCELL_X16 FILLER_71_851 ();
 FILLCELL_X2 FILLER_71_867 ();
 FILLCELL_X1 FILLER_71_869 ();
 FILLCELL_X1 FILLER_71_875 ();
 FILLCELL_X2 FILLER_71_879 ();
 FILLCELL_X1 FILLER_71_890 ();
 FILLCELL_X4 FILLER_71_898 ();
 FILLCELL_X1 FILLER_71_902 ();
 FILLCELL_X2 FILLER_71_915 ();
 FILLCELL_X32 FILLER_71_920 ();
 FILLCELL_X2 FILLER_71_952 ();
 FILLCELL_X2 FILLER_71_959 ();
 FILLCELL_X1 FILLER_71_961 ();
 FILLCELL_X4 FILLER_71_965 ();
 FILLCELL_X2 FILLER_71_969 ();
 FILLCELL_X1 FILLER_71_976 ();
 FILLCELL_X2 FILLER_71_982 ();
 FILLCELL_X2 FILLER_71_987 ();
 FILLCELL_X4 FILLER_71_996 ();
 FILLCELL_X2 FILLER_71_1000 ();
 FILLCELL_X1 FILLER_71_1002 ();
 FILLCELL_X8 FILLER_71_1006 ();
 FILLCELL_X1 FILLER_71_1014 ();
 FILLCELL_X16 FILLER_71_1032 ();
 FILLCELL_X8 FILLER_71_1053 ();
 FILLCELL_X2 FILLER_71_1061 ();
 FILLCELL_X1 FILLER_71_1063 ();
 FILLCELL_X8 FILLER_71_1073 ();
 FILLCELL_X2 FILLER_71_1081 ();
 FILLCELL_X16 FILLER_71_1100 ();
 FILLCELL_X2 FILLER_71_1116 ();
 FILLCELL_X1 FILLER_71_1118 ();
 FILLCELL_X2 FILLER_71_1143 ();
 FILLCELL_X1 FILLER_71_1145 ();
 FILLCELL_X4 FILLER_71_1163 ();
 FILLCELL_X1 FILLER_71_1167 ();
 FILLCELL_X16 FILLER_71_1175 ();
 FILLCELL_X2 FILLER_71_1191 ();
 FILLCELL_X2 FILLER_71_1217 ();
 FILLCELL_X1 FILLER_71_1219 ();
 FILLCELL_X4 FILLER_71_1223 ();
 FILLCELL_X2 FILLER_72_1 ();
 FILLCELL_X1 FILLER_72_3 ();
 FILLCELL_X32 FILLER_72_7 ();
 FILLCELL_X4 FILLER_72_39 ();
 FILLCELL_X2 FILLER_72_43 ();
 FILLCELL_X1 FILLER_72_45 ();
 FILLCELL_X1 FILLER_72_53 ();
 FILLCELL_X8 FILLER_72_61 ();
 FILLCELL_X2 FILLER_72_69 ();
 FILLCELL_X16 FILLER_72_78 ();
 FILLCELL_X2 FILLER_72_94 ();
 FILLCELL_X1 FILLER_72_96 ();
 FILLCELL_X1 FILLER_72_111 ();
 FILLCELL_X16 FILLER_72_123 ();
 FILLCELL_X16 FILLER_72_156 ();
 FILLCELL_X2 FILLER_72_189 ();
 FILLCELL_X4 FILLER_72_194 ();
 FILLCELL_X2 FILLER_72_198 ();
 FILLCELL_X2 FILLER_72_207 ();
 FILLCELL_X2 FILLER_72_226 ();
 FILLCELL_X8 FILLER_72_242 ();
 FILLCELL_X4 FILLER_72_257 ();
 FILLCELL_X1 FILLER_72_261 ();
 FILLCELL_X4 FILLER_72_282 ();
 FILLCELL_X1 FILLER_72_286 ();
 FILLCELL_X4 FILLER_72_294 ();
 FILLCELL_X4 FILLER_72_305 ();
 FILLCELL_X2 FILLER_72_309 ();
 FILLCELL_X1 FILLER_72_311 ();
 FILLCELL_X4 FILLER_72_336 ();
 FILLCELL_X2 FILLER_72_340 ();
 FILLCELL_X1 FILLER_72_342 ();
 FILLCELL_X32 FILLER_72_355 ();
 FILLCELL_X1 FILLER_72_387 ();
 FILLCELL_X4 FILLER_72_405 ();
 FILLCELL_X2 FILLER_72_409 ();
 FILLCELL_X2 FILLER_72_445 ();
 FILLCELL_X1 FILLER_72_447 ();
 FILLCELL_X4 FILLER_72_455 ();
 FILLCELL_X1 FILLER_72_470 ();
 FILLCELL_X4 FILLER_72_484 ();
 FILLCELL_X4 FILLER_72_495 ();
 FILLCELL_X2 FILLER_72_499 ();
 FILLCELL_X8 FILLER_72_508 ();
 FILLCELL_X2 FILLER_72_516 ();
 FILLCELL_X4 FILLER_72_547 ();
 FILLCELL_X2 FILLER_72_551 ();
 FILLCELL_X1 FILLER_72_553 ();
 FILLCELL_X16 FILLER_72_561 ();
 FILLCELL_X4 FILLER_72_594 ();
 FILLCELL_X2 FILLER_72_598 ();
 FILLCELL_X1 FILLER_72_600 ();
 FILLCELL_X2 FILLER_72_628 ();
 FILLCELL_X1 FILLER_72_630 ();
 FILLCELL_X16 FILLER_72_656 ();
 FILLCELL_X8 FILLER_72_672 ();
 FILLCELL_X4 FILLER_72_680 ();
 FILLCELL_X4 FILLER_72_691 ();
 FILLCELL_X4 FILLER_72_702 ();
 FILLCELL_X2 FILLER_72_706 ();
 FILLCELL_X1 FILLER_72_708 ();
 FILLCELL_X1 FILLER_72_739 ();
 FILLCELL_X4 FILLER_72_747 ();
 FILLCELL_X1 FILLER_72_751 ();
 FILLCELL_X8 FILLER_72_770 ();
 FILLCELL_X1 FILLER_72_778 ();
 FILLCELL_X4 FILLER_72_796 ();
 FILLCELL_X2 FILLER_72_807 ();
 FILLCELL_X1 FILLER_72_809 ();
 FILLCELL_X1 FILLER_72_818 ();
 FILLCELL_X1 FILLER_72_827 ();
 FILLCELL_X2 FILLER_72_838 ();
 FILLCELL_X8 FILLER_72_863 ();
 FILLCELL_X4 FILLER_72_871 ();
 FILLCELL_X2 FILLER_72_875 ();
 FILLCELL_X1 FILLER_72_877 ();
 FILLCELL_X1 FILLER_72_904 ();
 FILLCELL_X16 FILLER_72_914 ();
 FILLCELL_X4 FILLER_72_930 ();
 FILLCELL_X2 FILLER_72_939 ();
 FILLCELL_X16 FILLER_72_946 ();
 FILLCELL_X4 FILLER_72_962 ();
 FILLCELL_X1 FILLER_72_966 ();
 FILLCELL_X4 FILLER_72_981 ();
 FILLCELL_X8 FILLER_72_989 ();
 FILLCELL_X4 FILLER_72_997 ();
 FILLCELL_X2 FILLER_72_1001 ();
 FILLCELL_X4 FILLER_72_1006 ();
 FILLCELL_X1 FILLER_72_1010 ();
 FILLCELL_X16 FILLER_72_1016 ();
 FILLCELL_X8 FILLER_72_1032 ();
 FILLCELL_X1 FILLER_72_1040 ();
 FILLCELL_X16 FILLER_72_1058 ();
 FILLCELL_X8 FILLER_72_1074 ();
 FILLCELL_X4 FILLER_72_1082 ();
 FILLCELL_X2 FILLER_72_1086 ();
 FILLCELL_X8 FILLER_72_1095 ();
 FILLCELL_X2 FILLER_72_1103 ();
 FILLCELL_X16 FILLER_72_1112 ();
 FILLCELL_X8 FILLER_72_1142 ();
 FILLCELL_X1 FILLER_72_1150 ();
 FILLCELL_X1 FILLER_72_1158 ();
 FILLCELL_X4 FILLER_72_1187 ();
 FILLCELL_X2 FILLER_72_1238 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X2 FILLER_73_33 ();
 FILLCELL_X1 FILLER_73_59 ();
 FILLCELL_X1 FILLER_73_67 ();
 FILLCELL_X4 FILLER_73_75 ();
 FILLCELL_X2 FILLER_73_86 ();
 FILLCELL_X16 FILLER_73_95 ();
 FILLCELL_X8 FILLER_73_111 ();
 FILLCELL_X2 FILLER_73_126 ();
 FILLCELL_X2 FILLER_73_135 ();
 FILLCELL_X1 FILLER_73_137 ();
 FILLCELL_X8 FILLER_73_162 ();
 FILLCELL_X4 FILLER_73_170 ();
 FILLCELL_X2 FILLER_73_174 ();
 FILLCELL_X1 FILLER_73_176 ();
 FILLCELL_X8 FILLER_73_201 ();
 FILLCELL_X2 FILLER_73_209 ();
 FILLCELL_X1 FILLER_73_211 ();
 FILLCELL_X8 FILLER_73_217 ();
 FILLCELL_X2 FILLER_73_225 ();
 FILLCELL_X1 FILLER_73_227 ();
 FILLCELL_X16 FILLER_73_242 ();
 FILLCELL_X8 FILLER_73_258 ();
 FILLCELL_X2 FILLER_73_266 ();
 FILLCELL_X1 FILLER_73_268 ();
 FILLCELL_X1 FILLER_73_279 ();
 FILLCELL_X2 FILLER_73_297 ();
 FILLCELL_X2 FILLER_73_306 ();
 FILLCELL_X1 FILLER_73_308 ();
 FILLCELL_X4 FILLER_73_347 ();
 FILLCELL_X4 FILLER_73_358 ();
 FILLCELL_X4 FILLER_73_369 ();
 FILLCELL_X2 FILLER_73_380 ();
 FILLCELL_X1 FILLER_73_382 ();
 FILLCELL_X4 FILLER_73_400 ();
 FILLCELL_X1 FILLER_73_404 ();
 FILLCELL_X4 FILLER_73_419 ();
 FILLCELL_X1 FILLER_73_452 ();
 FILLCELL_X2 FILLER_73_463 ();
 FILLCELL_X1 FILLER_73_465 ();
 FILLCELL_X8 FILLER_73_471 ();
 FILLCELL_X1 FILLER_73_479 ();
 FILLCELL_X1 FILLER_73_504 ();
 FILLCELL_X16 FILLER_73_520 ();
 FILLCELL_X2 FILLER_73_536 ();
 FILLCELL_X1 FILLER_73_538 ();
 FILLCELL_X2 FILLER_73_546 ();
 FILLCELL_X8 FILLER_73_572 ();
 FILLCELL_X2 FILLER_73_580 ();
 FILLCELL_X4 FILLER_73_610 ();
 FILLCELL_X16 FILLER_73_635 ();
 FILLCELL_X8 FILLER_73_651 ();
 FILLCELL_X2 FILLER_73_659 ();
 FILLCELL_X8 FILLER_73_678 ();
 FILLCELL_X2 FILLER_73_686 ();
 FILLCELL_X16 FILLER_73_695 ();
 FILLCELL_X4 FILLER_73_773 ();
 FILLCELL_X2 FILLER_73_777 ();
 FILLCELL_X1 FILLER_73_779 ();
 FILLCELL_X4 FILLER_73_787 ();
 FILLCELL_X2 FILLER_73_791 ();
 FILLCELL_X16 FILLER_73_797 ();
 FILLCELL_X4 FILLER_73_813 ();
 FILLCELL_X1 FILLER_73_838 ();
 FILLCELL_X1 FILLER_73_854 ();
 FILLCELL_X16 FILLER_73_865 ();
 FILLCELL_X4 FILLER_73_881 ();
 FILLCELL_X2 FILLER_73_885 ();
 FILLCELL_X1 FILLER_73_896 ();
 FILLCELL_X16 FILLER_73_912 ();
 FILLCELL_X2 FILLER_73_928 ();
 FILLCELL_X1 FILLER_73_930 ();
 FILLCELL_X32 FILLER_73_955 ();
 FILLCELL_X16 FILLER_73_987 ();
 FILLCELL_X2 FILLER_73_1022 ();
 FILLCELL_X1 FILLER_73_1024 ();
 FILLCELL_X4 FILLER_73_1032 ();
 FILLCELL_X2 FILLER_73_1036 ();
 FILLCELL_X1 FILLER_73_1038 ();
 FILLCELL_X16 FILLER_73_1053 ();
 FILLCELL_X2 FILLER_73_1069 ();
 FILLCELL_X1 FILLER_73_1071 ();
 FILLCELL_X4 FILLER_73_1096 ();
 FILLCELL_X1 FILLER_73_1100 ();
 FILLCELL_X16 FILLER_73_1121 ();
 FILLCELL_X2 FILLER_73_1161 ();
 FILLCELL_X1 FILLER_73_1163 ();
 FILLCELL_X1 FILLER_73_1188 ();
 FILLCELL_X2 FILLER_73_1203 ();
 FILLCELL_X1 FILLER_73_1218 ();
 FILLCELL_X4 FILLER_73_1236 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X4 FILLER_74_33 ();
 FILLCELL_X2 FILLER_74_37 ();
 FILLCELL_X8 FILLER_74_56 ();
 FILLCELL_X2 FILLER_74_64 ();
 FILLCELL_X1 FILLER_74_66 ();
 FILLCELL_X2 FILLER_74_84 ();
 FILLCELL_X4 FILLER_74_110 ();
 FILLCELL_X1 FILLER_74_114 ();
 FILLCELL_X16 FILLER_74_139 ();
 FILLCELL_X4 FILLER_74_155 ();
 FILLCELL_X2 FILLER_74_159 ();
 FILLCELL_X2 FILLER_74_189 ();
 FILLCELL_X16 FILLER_74_202 ();
 FILLCELL_X2 FILLER_74_218 ();
 FILLCELL_X2 FILLER_74_261 ();
 FILLCELL_X2 FILLER_74_290 ();
 FILLCELL_X1 FILLER_74_292 ();
 FILLCELL_X4 FILLER_74_324 ();
 FILLCELL_X1 FILLER_74_393 ();
 FILLCELL_X32 FILLER_74_425 ();
 FILLCELL_X2 FILLER_74_457 ();
 FILLCELL_X1 FILLER_74_459 ();
 FILLCELL_X4 FILLER_74_464 ();
 FILLCELL_X16 FILLER_74_472 ();
 FILLCELL_X4 FILLER_74_488 ();
 FILLCELL_X2 FILLER_74_492 ();
 FILLCELL_X1 FILLER_74_494 ();
 FILLCELL_X1 FILLER_74_519 ();
 FILLCELL_X8 FILLER_74_527 ();
 FILLCELL_X4 FILLER_74_535 ();
 FILLCELL_X1 FILLER_74_539 ();
 FILLCELL_X8 FILLER_74_547 ();
 FILLCELL_X2 FILLER_74_555 ();
 FILLCELL_X1 FILLER_74_557 ();
 FILLCELL_X16 FILLER_74_565 ();
 FILLCELL_X1 FILLER_74_581 ();
 FILLCELL_X32 FILLER_74_589 ();
 FILLCELL_X8 FILLER_74_621 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X16 FILLER_74_632 ();
 FILLCELL_X2 FILLER_74_648 ();
 FILLCELL_X4 FILLER_74_655 ();
 FILLCELL_X2 FILLER_74_683 ();
 FILLCELL_X2 FILLER_74_764 ();
 FILLCELL_X2 FILLER_74_773 ();
 FILLCELL_X1 FILLER_74_775 ();
 FILLCELL_X4 FILLER_74_783 ();
 FILLCELL_X2 FILLER_74_787 ();
 FILLCELL_X1 FILLER_74_789 ();
 FILLCELL_X16 FILLER_74_814 ();
 FILLCELL_X2 FILLER_74_830 ();
 FILLCELL_X2 FILLER_74_837 ();
 FILLCELL_X32 FILLER_74_858 ();
 FILLCELL_X8 FILLER_74_890 ();
 FILLCELL_X2 FILLER_74_898 ();
 FILLCELL_X8 FILLER_74_907 ();
 FILLCELL_X4 FILLER_74_915 ();
 FILLCELL_X2 FILLER_74_919 ();
 FILLCELL_X2 FILLER_74_941 ();
 FILLCELL_X32 FILLER_74_948 ();
 FILLCELL_X4 FILLER_74_980 ();
 FILLCELL_X8 FILLER_74_990 ();
 FILLCELL_X4 FILLER_74_998 ();
 FILLCELL_X2 FILLER_74_1002 ();
 FILLCELL_X1 FILLER_74_1021 ();
 FILLCELL_X4 FILLER_74_1029 ();
 FILLCELL_X1 FILLER_74_1033 ();
 FILLCELL_X2 FILLER_74_1038 ();
 FILLCELL_X2 FILLER_74_1108 ();
 FILLCELL_X2 FILLER_74_1127 ();
 FILLCELL_X1 FILLER_74_1129 ();
 FILLCELL_X2 FILLER_74_1143 ();
 FILLCELL_X1 FILLER_74_1145 ();
 FILLCELL_X2 FILLER_74_1164 ();
 FILLCELL_X16 FILLER_74_1173 ();
 FILLCELL_X4 FILLER_74_1189 ();
 FILLCELL_X2 FILLER_74_1193 ();
 FILLCELL_X2 FILLER_74_1206 ();
 FILLCELL_X2 FILLER_74_1225 ();
 FILLCELL_X8 FILLER_75_1 ();
 FILLCELL_X4 FILLER_75_9 ();
 FILLCELL_X2 FILLER_75_13 ();
 FILLCELL_X1 FILLER_75_15 ();
 FILLCELL_X2 FILLER_75_20 ();
 FILLCELL_X32 FILLER_75_25 ();
 FILLCELL_X16 FILLER_75_57 ();
 FILLCELL_X8 FILLER_75_73 ();
 FILLCELL_X4 FILLER_75_81 ();
 FILLCELL_X8 FILLER_75_109 ();
 FILLCELL_X4 FILLER_75_117 ();
 FILLCELL_X2 FILLER_75_121 ();
 FILLCELL_X1 FILLER_75_123 ();
 FILLCELL_X16 FILLER_75_141 ();
 FILLCELL_X2 FILLER_75_157 ();
 FILLCELL_X2 FILLER_75_176 ();
 FILLCELL_X1 FILLER_75_178 ();
 FILLCELL_X4 FILLER_75_186 ();
 FILLCELL_X4 FILLER_75_214 ();
 FILLCELL_X2 FILLER_75_218 ();
 FILLCELL_X4 FILLER_75_244 ();
 FILLCELL_X4 FILLER_75_262 ();
 FILLCELL_X2 FILLER_75_266 ();
 FILLCELL_X2 FILLER_75_296 ();
 FILLCELL_X1 FILLER_75_298 ();
 FILLCELL_X2 FILLER_75_330 ();
 FILLCELL_X1 FILLER_75_332 ();
 FILLCELL_X32 FILLER_75_357 ();
 FILLCELL_X32 FILLER_75_389 ();
 FILLCELL_X16 FILLER_75_421 ();
 FILLCELL_X8 FILLER_75_437 ();
 FILLCELL_X2 FILLER_75_445 ();
 FILLCELL_X1 FILLER_75_447 ();
 FILLCELL_X8 FILLER_75_455 ();
 FILLCELL_X4 FILLER_75_463 ();
 FILLCELL_X2 FILLER_75_467 ();
 FILLCELL_X1 FILLER_75_469 ();
 FILLCELL_X4 FILLER_75_524 ();
 FILLCELL_X1 FILLER_75_528 ();
 FILLCELL_X16 FILLER_75_536 ();
 FILLCELL_X2 FILLER_75_552 ();
 FILLCELL_X2 FILLER_75_595 ();
 FILLCELL_X2 FILLER_75_604 ();
 FILLCELL_X4 FILLER_75_637 ();
 FILLCELL_X2 FILLER_75_641 ();
 FILLCELL_X2 FILLER_75_669 ();
 FILLCELL_X1 FILLER_75_671 ();
 FILLCELL_X32 FILLER_75_683 ();
 FILLCELL_X32 FILLER_75_715 ();
 FILLCELL_X4 FILLER_75_747 ();
 FILLCELL_X1 FILLER_75_751 ();
 FILLCELL_X1 FILLER_75_763 ();
 FILLCELL_X8 FILLER_75_794 ();
 FILLCELL_X4 FILLER_75_802 ();
 FILLCELL_X4 FILLER_75_811 ();
 FILLCELL_X1 FILLER_75_818 ();
 FILLCELL_X8 FILLER_75_824 ();
 FILLCELL_X32 FILLER_75_842 ();
 FILLCELL_X8 FILLER_75_874 ();
 FILLCELL_X4 FILLER_75_882 ();
 FILLCELL_X2 FILLER_75_886 ();
 FILLCELL_X1 FILLER_75_888 ();
 FILLCELL_X16 FILLER_75_896 ();
 FILLCELL_X8 FILLER_75_912 ();
 FILLCELL_X2 FILLER_75_920 ();
 FILLCELL_X4 FILLER_75_940 ();
 FILLCELL_X1 FILLER_75_949 ();
 FILLCELL_X8 FILLER_75_953 ();
 FILLCELL_X4 FILLER_75_961 ();
 FILLCELL_X2 FILLER_75_978 ();
 FILLCELL_X2 FILLER_75_992 ();
 FILLCELL_X1 FILLER_75_994 ();
 FILLCELL_X16 FILLER_75_1001 ();
 FILLCELL_X1 FILLER_75_1017 ();
 FILLCELL_X4 FILLER_75_1025 ();
 FILLCELL_X2 FILLER_75_1029 ();
 FILLCELL_X1 FILLER_75_1038 ();
 FILLCELL_X2 FILLER_75_1052 ();
 FILLCELL_X2 FILLER_75_1071 ();
 FILLCELL_X2 FILLER_75_1080 ();
 FILLCELL_X4 FILLER_75_1096 ();
 FILLCELL_X2 FILLER_75_1100 ();
 FILLCELL_X1 FILLER_75_1109 ();
 FILLCELL_X16 FILLER_75_1139 ();
 FILLCELL_X2 FILLER_75_1155 ();
 FILLCELL_X1 FILLER_75_1157 ();
 FILLCELL_X16 FILLER_75_1165 ();
 FILLCELL_X8 FILLER_75_1181 ();
 FILLCELL_X2 FILLER_75_1189 ();
 FILLCELL_X1 FILLER_75_1222 ();
 FILLCELL_X8 FILLER_76_1 ();
 FILLCELL_X4 FILLER_76_9 ();
 FILLCELL_X1 FILLER_76_13 ();
 FILLCELL_X32 FILLER_76_21 ();
 FILLCELL_X4 FILLER_76_53 ();
 FILLCELL_X2 FILLER_76_57 ();
 FILLCELL_X16 FILLER_76_76 ();
 FILLCELL_X1 FILLER_76_92 ();
 FILLCELL_X8 FILLER_76_98 ();
 FILLCELL_X1 FILLER_76_106 ();
 FILLCELL_X32 FILLER_76_138 ();
 FILLCELL_X16 FILLER_76_170 ();
 FILLCELL_X8 FILLER_76_186 ();
 FILLCELL_X2 FILLER_76_194 ();
 FILLCELL_X1 FILLER_76_196 ();
 FILLCELL_X2 FILLER_76_204 ();
 FILLCELL_X1 FILLER_76_206 ();
 FILLCELL_X8 FILLER_76_255 ();
 FILLCELL_X4 FILLER_76_263 ();
 FILLCELL_X2 FILLER_76_267 ();
 FILLCELL_X1 FILLER_76_269 ();
 FILLCELL_X16 FILLER_76_302 ();
 FILLCELL_X8 FILLER_76_318 ();
 FILLCELL_X1 FILLER_76_326 ();
 FILLCELL_X2 FILLER_76_334 ();
 FILLCELL_X32 FILLER_76_357 ();
 FILLCELL_X16 FILLER_76_389 ();
 FILLCELL_X4 FILLER_76_405 ();
 FILLCELL_X2 FILLER_76_409 ();
 FILLCELL_X2 FILLER_76_444 ();
 FILLCELL_X1 FILLER_76_446 ();
 FILLCELL_X2 FILLER_76_464 ();
 FILLCELL_X4 FILLER_76_490 ();
 FILLCELL_X2 FILLER_76_494 ();
 FILLCELL_X2 FILLER_76_502 ();
 FILLCELL_X8 FILLER_76_508 ();
 FILLCELL_X1 FILLER_76_516 ();
 FILLCELL_X8 FILLER_76_520 ();
 FILLCELL_X1 FILLER_76_528 ();
 FILLCELL_X1 FILLER_76_540 ();
 FILLCELL_X1 FILLER_76_558 ();
 FILLCELL_X1 FILLER_76_566 ();
 FILLCELL_X1 FILLER_76_591 ();
 FILLCELL_X1 FILLER_76_599 ();
 FILLCELL_X16 FILLER_76_639 ();
 FILLCELL_X8 FILLER_76_655 ();
 FILLCELL_X2 FILLER_76_663 ();
 FILLCELL_X1 FILLER_76_665 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X16 FILLER_76_728 ();
 FILLCELL_X2 FILLER_76_744 ();
 FILLCELL_X32 FILLER_76_753 ();
 FILLCELL_X2 FILLER_76_785 ();
 FILLCELL_X1 FILLER_76_787 ();
 FILLCELL_X8 FILLER_76_795 ();
 FILLCELL_X1 FILLER_76_812 ();
 FILLCELL_X1 FILLER_76_816 ();
 FILLCELL_X2 FILLER_76_826 ();
 FILLCELL_X4 FILLER_76_833 ();
 FILLCELL_X2 FILLER_76_837 ();
 FILLCELL_X8 FILLER_76_843 ();
 FILLCELL_X1 FILLER_76_851 ();
 FILLCELL_X4 FILLER_76_857 ();
 FILLCELL_X2 FILLER_76_861 ();
 FILLCELL_X1 FILLER_76_863 ();
 FILLCELL_X4 FILLER_76_871 ();
 FILLCELL_X1 FILLER_76_875 ();
 FILLCELL_X8 FILLER_76_904 ();
 FILLCELL_X1 FILLER_76_912 ();
 FILLCELL_X2 FILLER_76_920 ();
 FILLCELL_X1 FILLER_76_922 ();
 FILLCELL_X2 FILLER_76_929 ();
 FILLCELL_X8 FILLER_76_949 ();
 FILLCELL_X4 FILLER_76_957 ();
 FILLCELL_X1 FILLER_76_961 ();
 FILLCELL_X2 FILLER_76_993 ();
 FILLCELL_X8 FILLER_76_999 ();
 FILLCELL_X4 FILLER_76_1007 ();
 FILLCELL_X1 FILLER_76_1011 ();
 FILLCELL_X32 FILLER_76_1025 ();
 FILLCELL_X8 FILLER_76_1057 ();
 FILLCELL_X4 FILLER_76_1065 ();
 FILLCELL_X1 FILLER_76_1069 ();
 FILLCELL_X8 FILLER_76_1081 ();
 FILLCELL_X4 FILLER_76_1089 ();
 FILLCELL_X4 FILLER_76_1106 ();
 FILLCELL_X1 FILLER_76_1110 ();
 FILLCELL_X4 FILLER_76_1118 ();
 FILLCELL_X1 FILLER_76_1122 ();
 FILLCELL_X2 FILLER_76_1130 ();
 FILLCELL_X8 FILLER_76_1145 ();
 FILLCELL_X4 FILLER_76_1153 ();
 FILLCELL_X16 FILLER_76_1170 ();
 FILLCELL_X2 FILLER_76_1186 ();
 FILLCELL_X1 FILLER_76_1239 ();
 FILLCELL_X4 FILLER_77_1 ();
 FILLCELL_X1 FILLER_77_5 ();
 FILLCELL_X32 FILLER_77_9 ();
 FILLCELL_X4 FILLER_77_41 ();
 FILLCELL_X1 FILLER_77_45 ();
 FILLCELL_X4 FILLER_77_53 ();
 FILLCELL_X2 FILLER_77_57 ();
 FILLCELL_X1 FILLER_77_59 ();
 FILLCELL_X8 FILLER_77_67 ();
 FILLCELL_X2 FILLER_77_75 ();
 FILLCELL_X1 FILLER_77_77 ();
 FILLCELL_X8 FILLER_77_82 ();
 FILLCELL_X1 FILLER_77_90 ();
 FILLCELL_X2 FILLER_77_123 ();
 FILLCELL_X1 FILLER_77_125 ();
 FILLCELL_X2 FILLER_77_133 ();
 FILLCELL_X4 FILLER_77_142 ();
 FILLCELL_X2 FILLER_77_146 ();
 FILLCELL_X1 FILLER_77_148 ();
 FILLCELL_X16 FILLER_77_152 ();
 FILLCELL_X4 FILLER_77_168 ();
 FILLCELL_X2 FILLER_77_172 ();
 FILLCELL_X1 FILLER_77_174 ();
 FILLCELL_X2 FILLER_77_192 ();
 FILLCELL_X1 FILLER_77_194 ();
 FILLCELL_X8 FILLER_77_214 ();
 FILLCELL_X2 FILLER_77_222 ();
 FILLCELL_X1 FILLER_77_224 ();
 FILLCELL_X2 FILLER_77_232 ();
 FILLCELL_X4 FILLER_77_263 ();
 FILLCELL_X2 FILLER_77_267 ();
 FILLCELL_X16 FILLER_77_286 ();
 FILLCELL_X8 FILLER_77_302 ();
 FILLCELL_X4 FILLER_77_310 ();
 FILLCELL_X2 FILLER_77_314 ();
 FILLCELL_X1 FILLER_77_316 ();
 FILLCELL_X2 FILLER_77_331 ();
 FILLCELL_X4 FILLER_77_360 ();
 FILLCELL_X1 FILLER_77_364 ();
 FILLCELL_X4 FILLER_77_382 ();
 FILLCELL_X8 FILLER_77_408 ();
 FILLCELL_X4 FILLER_77_440 ();
 FILLCELL_X2 FILLER_77_444 ();
 FILLCELL_X2 FILLER_77_470 ();
 FILLCELL_X1 FILLER_77_472 ();
 FILLCELL_X16 FILLER_77_490 ();
 FILLCELL_X2 FILLER_77_506 ();
 FILLCELL_X1 FILLER_77_508 ();
 FILLCELL_X4 FILLER_77_515 ();
 FILLCELL_X2 FILLER_77_524 ();
 FILLCELL_X1 FILLER_77_526 ();
 FILLCELL_X2 FILLER_77_539 ();
 FILLCELL_X1 FILLER_77_541 ();
 FILLCELL_X2 FILLER_77_551 ();
 FILLCELL_X1 FILLER_77_553 ();
 FILLCELL_X4 FILLER_77_571 ();
 FILLCELL_X2 FILLER_77_575 ();
 FILLCELL_X2 FILLER_77_591 ();
 FILLCELL_X4 FILLER_77_600 ();
 FILLCELL_X2 FILLER_77_613 ();
 FILLCELL_X1 FILLER_77_615 ();
 FILLCELL_X8 FILLER_77_623 ();
 FILLCELL_X2 FILLER_77_631 ();
 FILLCELL_X8 FILLER_77_650 ();
 FILLCELL_X1 FILLER_77_658 ();
 FILLCELL_X4 FILLER_77_666 ();
 FILLCELL_X2 FILLER_77_677 ();
 FILLCELL_X4 FILLER_77_690 ();
 FILLCELL_X1 FILLER_77_725 ();
 FILLCELL_X8 FILLER_77_730 ();
 FILLCELL_X4 FILLER_77_738 ();
 FILLCELL_X4 FILLER_77_759 ();
 FILLCELL_X2 FILLER_77_763 ();
 FILLCELL_X4 FILLER_77_782 ();
 FILLCELL_X2 FILLER_77_786 ();
 FILLCELL_X1 FILLER_77_816 ();
 FILLCELL_X2 FILLER_77_835 ();
 FILLCELL_X4 FILLER_77_846 ();
 FILLCELL_X2 FILLER_77_850 ();
 FILLCELL_X4 FILLER_77_857 ();
 FILLCELL_X1 FILLER_77_884 ();
 FILLCELL_X32 FILLER_77_902 ();
 FILLCELL_X16 FILLER_77_934 ();
 FILLCELL_X8 FILLER_77_950 ();
 FILLCELL_X4 FILLER_77_958 ();
 FILLCELL_X1 FILLER_77_975 ();
 FILLCELL_X2 FILLER_77_979 ();
 FILLCELL_X1 FILLER_77_981 ();
 FILLCELL_X4 FILLER_77_991 ();
 FILLCELL_X1 FILLER_77_995 ();
 FILLCELL_X1 FILLER_77_999 ();
 FILLCELL_X1 FILLER_77_1013 ();
 FILLCELL_X8 FILLER_77_1024 ();
 FILLCELL_X2 FILLER_77_1032 ();
 FILLCELL_X4 FILLER_77_1038 ();
 FILLCELL_X1 FILLER_77_1042 ();
 FILLCELL_X16 FILLER_77_1065 ();
 FILLCELL_X8 FILLER_77_1081 ();
 FILLCELL_X4 FILLER_77_1089 ();
 FILLCELL_X2 FILLER_77_1104 ();
 FILLCELL_X4 FILLER_77_1130 ();
 FILLCELL_X1 FILLER_77_1193 ();
 FILLCELL_X1 FILLER_77_1201 ();
 FILLCELL_X2 FILLER_77_1215 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X2 FILLER_78_33 ();
 FILLCELL_X1 FILLER_78_83 ();
 FILLCELL_X8 FILLER_78_91 ();
 FILLCELL_X8 FILLER_78_113 ();
 FILLCELL_X4 FILLER_78_121 ();
 FILLCELL_X1 FILLER_78_125 ();
 FILLCELL_X2 FILLER_78_133 ();
 FILLCELL_X1 FILLER_78_135 ();
 FILLCELL_X1 FILLER_78_158 ();
 FILLCELL_X1 FILLER_78_173 ();
 FILLCELL_X2 FILLER_78_188 ();
 FILLCELL_X1 FILLER_78_190 ();
 FILLCELL_X2 FILLER_78_198 ();
 FILLCELL_X1 FILLER_78_200 ();
 FILLCELL_X8 FILLER_78_208 ();
 FILLCELL_X4 FILLER_78_216 ();
 FILLCELL_X1 FILLER_78_220 ();
 FILLCELL_X2 FILLER_78_228 ();
 FILLCELL_X1 FILLER_78_230 ();
 FILLCELL_X8 FILLER_78_252 ();
 FILLCELL_X4 FILLER_78_260 ();
 FILLCELL_X1 FILLER_78_264 ();
 FILLCELL_X16 FILLER_78_282 ();
 FILLCELL_X2 FILLER_78_298 ();
 FILLCELL_X1 FILLER_78_300 ();
 FILLCELL_X4 FILLER_78_323 ();
 FILLCELL_X2 FILLER_78_327 ();
 FILLCELL_X8 FILLER_78_336 ();
 FILLCELL_X4 FILLER_78_344 ();
 FILLCELL_X2 FILLER_78_348 ();
 FILLCELL_X1 FILLER_78_350 ();
 FILLCELL_X1 FILLER_78_382 ();
 FILLCELL_X4 FILLER_78_407 ();
 FILLCELL_X2 FILLER_78_411 ();
 FILLCELL_X2 FILLER_78_422 ();
 FILLCELL_X2 FILLER_78_433 ();
 FILLCELL_X1 FILLER_78_435 ();
 FILLCELL_X2 FILLER_78_443 ();
 FILLCELL_X1 FILLER_78_453 ();
 FILLCELL_X2 FILLER_78_468 ();
 FILLCELL_X4 FILLER_78_502 ();
 FILLCELL_X2 FILLER_78_506 ();
 FILLCELL_X1 FILLER_78_534 ();
 FILLCELL_X4 FILLER_78_539 ();
 FILLCELL_X16 FILLER_78_546 ();
 FILLCELL_X2 FILLER_78_562 ();
 FILLCELL_X16 FILLER_78_581 ();
 FILLCELL_X1 FILLER_78_597 ();
 FILLCELL_X8 FILLER_78_618 ();
 FILLCELL_X4 FILLER_78_626 ();
 FILLCELL_X1 FILLER_78_630 ();
 FILLCELL_X16 FILLER_78_632 ();
 FILLCELL_X8 FILLER_78_648 ();
 FILLCELL_X2 FILLER_78_656 ();
 FILLCELL_X8 FILLER_78_675 ();
 FILLCELL_X2 FILLER_78_683 ();
 FILLCELL_X1 FILLER_78_709 ();
 FILLCELL_X2 FILLER_78_727 ();
 FILLCELL_X2 FILLER_78_742 ();
 FILLCELL_X1 FILLER_78_778 ();
 FILLCELL_X1 FILLER_78_786 ();
 FILLCELL_X2 FILLER_78_804 ();
 FILLCELL_X1 FILLER_78_806 ();
 FILLCELL_X4 FILLER_78_844 ();
 FILLCELL_X1 FILLER_78_848 ();
 FILLCELL_X1 FILLER_78_861 ();
 FILLCELL_X2 FILLER_78_871 ();
 FILLCELL_X2 FILLER_78_897 ();
 FILLCELL_X2 FILLER_78_919 ();
 FILLCELL_X2 FILLER_78_933 ();
 FILLCELL_X1 FILLER_78_935 ();
 FILLCELL_X2 FILLER_78_943 ();
 FILLCELL_X4 FILLER_78_952 ();
 FILLCELL_X1 FILLER_78_956 ();
 FILLCELL_X8 FILLER_78_960 ();
 FILLCELL_X8 FILLER_78_973 ();
 FILLCELL_X4 FILLER_78_981 ();
 FILLCELL_X8 FILLER_78_992 ();
 FILLCELL_X2 FILLER_78_1000 ();
 FILLCELL_X1 FILLER_78_1034 ();
 FILLCELL_X4 FILLER_78_1048 ();
 FILLCELL_X1 FILLER_78_1066 ();
 FILLCELL_X32 FILLER_78_1084 ();
 FILLCELL_X4 FILLER_78_1116 ();
 FILLCELL_X1 FILLER_78_1120 ();
 FILLCELL_X4 FILLER_78_1135 ();
 FILLCELL_X2 FILLER_78_1139 ();
 FILLCELL_X8 FILLER_78_1148 ();
 FILLCELL_X4 FILLER_78_1156 ();
 FILLCELL_X2 FILLER_78_1160 ();
 FILLCELL_X4 FILLER_78_1176 ();
 FILLCELL_X2 FILLER_78_1180 ();
 FILLCELL_X1 FILLER_78_1189 ();
 FILLCELL_X8 FILLER_78_1210 ();
 FILLCELL_X16 FILLER_78_1221 ();
 FILLCELL_X2 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_7 ();
 FILLCELL_X2 FILLER_79_39 ();
 FILLCELL_X1 FILLER_79_41 ();
 FILLCELL_X1 FILLER_79_59 ();
 FILLCELL_X8 FILLER_79_79 ();
 FILLCELL_X1 FILLER_79_87 ();
 FILLCELL_X16 FILLER_79_105 ();
 FILLCELL_X2 FILLER_79_121 ();
 FILLCELL_X16 FILLER_79_140 ();
 FILLCELL_X1 FILLER_79_156 ();
 FILLCELL_X4 FILLER_79_174 ();
 FILLCELL_X32 FILLER_79_202 ();
 FILLCELL_X32 FILLER_79_234 ();
 FILLCELL_X8 FILLER_79_294 ();
 FILLCELL_X4 FILLER_79_302 ();
 FILLCELL_X1 FILLER_79_306 ();
 FILLCELL_X4 FILLER_79_324 ();
 FILLCELL_X1 FILLER_79_328 ();
 FILLCELL_X8 FILLER_79_360 ();
 FILLCELL_X2 FILLER_79_368 ();
 FILLCELL_X1 FILLER_79_370 ();
 FILLCELL_X2 FILLER_79_385 ();
 FILLCELL_X1 FILLER_79_387 ();
 FILLCELL_X8 FILLER_79_402 ();
 FILLCELL_X2 FILLER_79_410 ();
 FILLCELL_X8 FILLER_79_429 ();
 FILLCELL_X1 FILLER_79_437 ();
 FILLCELL_X16 FILLER_79_449 ();
 FILLCELL_X8 FILLER_79_465 ();
 FILLCELL_X4 FILLER_79_473 ();
 FILLCELL_X32 FILLER_79_480 ();
 FILLCELL_X4 FILLER_79_512 ();
 FILLCELL_X1 FILLER_79_516 ();
 FILLCELL_X2 FILLER_79_543 ();
 FILLCELL_X16 FILLER_79_554 ();
 FILLCELL_X4 FILLER_79_570 ();
 FILLCELL_X2 FILLER_79_574 ();
 FILLCELL_X1 FILLER_79_576 ();
 FILLCELL_X16 FILLER_79_582 ();
 FILLCELL_X4 FILLER_79_598 ();
 FILLCELL_X2 FILLER_79_602 ();
 FILLCELL_X1 FILLER_79_608 ();
 FILLCELL_X32 FILLER_79_618 ();
 FILLCELL_X4 FILLER_79_650 ();
 FILLCELL_X2 FILLER_79_654 ();
 FILLCELL_X16 FILLER_79_680 ();
 FILLCELL_X1 FILLER_79_696 ();
 FILLCELL_X2 FILLER_79_712 ();
 FILLCELL_X1 FILLER_79_714 ();
 FILLCELL_X2 FILLER_79_722 ();
 FILLCELL_X1 FILLER_79_724 ();
 FILLCELL_X2 FILLER_79_732 ();
 FILLCELL_X4 FILLER_79_741 ();
 FILLCELL_X1 FILLER_79_759 ();
 FILLCELL_X2 FILLER_79_767 ();
 FILLCELL_X2 FILLER_79_776 ();
 FILLCELL_X2 FILLER_79_785 ();
 FILLCELL_X4 FILLER_79_805 ();
 FILLCELL_X2 FILLER_79_809 ();
 FILLCELL_X4 FILLER_79_818 ();
 FILLCELL_X2 FILLER_79_825 ();
 FILLCELL_X1 FILLER_79_834 ();
 FILLCELL_X4 FILLER_79_838 ();
 FILLCELL_X1 FILLER_79_842 ();
 FILLCELL_X1 FILLER_79_860 ();
 FILLCELL_X4 FILLER_79_876 ();
 FILLCELL_X2 FILLER_79_880 ();
 FILLCELL_X1 FILLER_79_882 ();
 FILLCELL_X4 FILLER_79_926 ();
 FILLCELL_X2 FILLER_79_930 ();
 FILLCELL_X1 FILLER_79_951 ();
 FILLCELL_X2 FILLER_79_967 ();
 FILLCELL_X1 FILLER_79_969 ();
 FILLCELL_X16 FILLER_79_982 ();
 FILLCELL_X1 FILLER_79_998 ();
 FILLCELL_X1 FILLER_79_1033 ();
 FILLCELL_X2 FILLER_79_1076 ();
 FILLCELL_X1 FILLER_79_1078 ();
 FILLCELL_X4 FILLER_79_1103 ();
 FILLCELL_X2 FILLER_79_1107 ();
 FILLCELL_X2 FILLER_79_1140 ();
 FILLCELL_X1 FILLER_79_1142 ();
 FILLCELL_X2 FILLER_79_1160 ();
 FILLCELL_X8 FILLER_79_1191 ();
 FILLCELL_X2 FILLER_79_1199 ();
 FILLCELL_X1 FILLER_79_1208 ();
 FILLCELL_X1 FILLER_79_1219 ();
 FILLCELL_X2 FILLER_79_1238 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X16 FILLER_80_33 ();
 FILLCELL_X8 FILLER_80_49 ();
 FILLCELL_X1 FILLER_80_57 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X16 FILLER_80_129 ();
 FILLCELL_X2 FILLER_80_145 ();
 FILLCELL_X1 FILLER_80_147 ();
 FILLCELL_X16 FILLER_80_172 ();
 FILLCELL_X4 FILLER_80_188 ();
 FILLCELL_X1 FILLER_80_192 ();
 FILLCELL_X4 FILLER_80_200 ();
 FILLCELL_X2 FILLER_80_204 ();
 FILLCELL_X8 FILLER_80_213 ();
 FILLCELL_X4 FILLER_80_221 ();
 FILLCELL_X2 FILLER_80_225 ();
 FILLCELL_X1 FILLER_80_227 ();
 FILLCELL_X32 FILLER_80_235 ();
 FILLCELL_X1 FILLER_80_267 ();
 FILLCELL_X8 FILLER_80_292 ();
 FILLCELL_X4 FILLER_80_300 ();
 FILLCELL_X2 FILLER_80_304 ();
 FILLCELL_X1 FILLER_80_306 ();
 FILLCELL_X2 FILLER_80_321 ();
 FILLCELL_X1 FILLER_80_323 ();
 FILLCELL_X1 FILLER_80_338 ();
 FILLCELL_X32 FILLER_80_363 ();
 FILLCELL_X4 FILLER_80_395 ();
 FILLCELL_X4 FILLER_80_413 ();
 FILLCELL_X2 FILLER_80_417 ();
 FILLCELL_X1 FILLER_80_419 ();
 FILLCELL_X16 FILLER_80_470 ();
 FILLCELL_X8 FILLER_80_486 ();
 FILLCELL_X2 FILLER_80_494 ();
 FILLCELL_X1 FILLER_80_509 ();
 FILLCELL_X1 FILLER_80_516 ();
 FILLCELL_X1 FILLER_80_521 ();
 FILLCELL_X2 FILLER_80_528 ();
 FILLCELL_X1 FILLER_80_534 ();
 FILLCELL_X2 FILLER_80_552 ();
 FILLCELL_X2 FILLER_80_571 ();
 FILLCELL_X2 FILLER_80_580 ();
 FILLCELL_X4 FILLER_80_592 ();
 FILLCELL_X8 FILLER_80_603 ();
 FILLCELL_X8 FILLER_80_618 ();
 FILLCELL_X4 FILLER_80_626 ();
 FILLCELL_X1 FILLER_80_630 ();
 FILLCELL_X8 FILLER_80_639 ();
 FILLCELL_X32 FILLER_80_678 ();
 FILLCELL_X1 FILLER_80_710 ();
 FILLCELL_X8 FILLER_80_728 ();
 FILLCELL_X4 FILLER_80_736 ();
 FILLCELL_X2 FILLER_80_740 ();
 FILLCELL_X8 FILLER_80_748 ();
 FILLCELL_X4 FILLER_80_756 ();
 FILLCELL_X2 FILLER_80_760 ();
 FILLCELL_X16 FILLER_80_770 ();
 FILLCELL_X4 FILLER_80_786 ();
 FILLCELL_X2 FILLER_80_790 ();
 FILLCELL_X1 FILLER_80_792 ();
 FILLCELL_X16 FILLER_80_811 ();
 FILLCELL_X8 FILLER_80_827 ();
 FILLCELL_X1 FILLER_80_835 ();
 FILLCELL_X4 FILLER_80_843 ();
 FILLCELL_X2 FILLER_80_847 ();
 FILLCELL_X1 FILLER_80_849 ();
 FILLCELL_X2 FILLER_80_855 ();
 FILLCELL_X1 FILLER_80_857 ();
 FILLCELL_X2 FILLER_80_885 ();
 FILLCELL_X1 FILLER_80_887 ();
 FILLCELL_X1 FILLER_80_896 ();
 FILLCELL_X1 FILLER_80_900 ();
 FILLCELL_X2 FILLER_80_906 ();
 FILLCELL_X2 FILLER_80_913 ();
 FILLCELL_X2 FILLER_80_928 ();
 FILLCELL_X1 FILLER_80_930 ();
 FILLCELL_X1 FILLER_80_948 ();
 FILLCELL_X1 FILLER_80_961 ();
 FILLCELL_X1 FILLER_80_967 ();
 FILLCELL_X8 FILLER_80_987 ();
 FILLCELL_X1 FILLER_80_1001 ();
 FILLCELL_X2 FILLER_80_1011 ();
 FILLCELL_X2 FILLER_80_1030 ();
 FILLCELL_X4 FILLER_80_1039 ();
 FILLCELL_X8 FILLER_80_1050 ();
 FILLCELL_X4 FILLER_80_1058 ();
 FILLCELL_X1 FILLER_80_1062 ();
 FILLCELL_X1 FILLER_80_1087 ();
 FILLCELL_X8 FILLER_80_1095 ();
 FILLCELL_X2 FILLER_80_1103 ();
 FILLCELL_X1 FILLER_80_1105 ();
 FILLCELL_X16 FILLER_80_1147 ();
 FILLCELL_X4 FILLER_80_1163 ();
 FILLCELL_X2 FILLER_80_1167 ();
 FILLCELL_X8 FILLER_80_1172 ();
 FILLCELL_X1 FILLER_80_1180 ();
 FILLCELL_X2 FILLER_80_1194 ();
 FILLCELL_X1 FILLER_80_1203 ();
 FILLCELL_X2 FILLER_80_1207 ();
 FILLCELL_X1 FILLER_80_1209 ();
 FILLCELL_X2 FILLER_80_1213 ();
 FILLCELL_X1 FILLER_80_1215 ();
 FILLCELL_X2 FILLER_80_1219 ();
 FILLCELL_X1 FILLER_80_1221 ();
 FILLCELL_X1 FILLER_80_1239 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X16 FILLER_81_33 ();
 FILLCELL_X8 FILLER_81_49 ();
 FILLCELL_X2 FILLER_81_57 ();
 FILLCELL_X8 FILLER_81_66 ();
 FILLCELL_X2 FILLER_81_74 ();
 FILLCELL_X8 FILLER_81_100 ();
 FILLCELL_X2 FILLER_81_108 ();
 FILLCELL_X1 FILLER_81_110 ();
 FILLCELL_X16 FILLER_81_125 ();
 FILLCELL_X4 FILLER_81_141 ();
 FILLCELL_X2 FILLER_81_145 ();
 FILLCELL_X1 FILLER_81_154 ();
 FILLCELL_X1 FILLER_81_172 ();
 FILLCELL_X2 FILLER_81_190 ();
 FILLCELL_X1 FILLER_81_199 ();
 FILLCELL_X2 FILLER_81_207 ();
 FILLCELL_X16 FILLER_81_226 ();
 FILLCELL_X8 FILLER_81_266 ();
 FILLCELL_X2 FILLER_81_274 ();
 FILLCELL_X1 FILLER_81_276 ();
 FILLCELL_X32 FILLER_81_284 ();
 FILLCELL_X8 FILLER_81_316 ();
 FILLCELL_X2 FILLER_81_324 ();
 FILLCELL_X4 FILLER_81_343 ();
 FILLCELL_X2 FILLER_81_347 ();
 FILLCELL_X1 FILLER_81_349 ();
 FILLCELL_X2 FILLER_81_362 ();
 FILLCELL_X8 FILLER_81_371 ();
 FILLCELL_X2 FILLER_81_379 ();
 FILLCELL_X1 FILLER_81_381 ();
 FILLCELL_X16 FILLER_81_406 ();
 FILLCELL_X2 FILLER_81_453 ();
 FILLCELL_X1 FILLER_81_455 ();
 FILLCELL_X4 FILLER_81_480 ();
 FILLCELL_X2 FILLER_81_484 ();
 FILLCELL_X1 FILLER_81_530 ();
 FILLCELL_X2 FILLER_81_572 ();
 FILLCELL_X4 FILLER_81_591 ();
 FILLCELL_X1 FILLER_81_595 ();
 FILLCELL_X8 FILLER_81_647 ();
 FILLCELL_X4 FILLER_81_655 ();
 FILLCELL_X1 FILLER_81_659 ();
 FILLCELL_X16 FILLER_81_668 ();
 FILLCELL_X4 FILLER_81_698 ();
 FILLCELL_X32 FILLER_81_709 ();
 FILLCELL_X1 FILLER_81_741 ();
 FILLCELL_X2 FILLER_81_749 ();
 FILLCELL_X16 FILLER_81_775 ();
 FILLCELL_X4 FILLER_81_805 ();
 FILLCELL_X2 FILLER_81_809 ();
 FILLCELL_X1 FILLER_81_828 ();
 FILLCELL_X2 FILLER_81_837 ();
 FILLCELL_X1 FILLER_81_839 ();
 FILLCELL_X1 FILLER_81_849 ();
 FILLCELL_X2 FILLER_81_853 ();
 FILLCELL_X2 FILLER_81_874 ();
 FILLCELL_X8 FILLER_81_883 ();
 FILLCELL_X1 FILLER_81_891 ();
 FILLCELL_X8 FILLER_81_897 ();
 FILLCELL_X1 FILLER_81_905 ();
 FILLCELL_X2 FILLER_81_911 ();
 FILLCELL_X1 FILLER_81_913 ();
 FILLCELL_X2 FILLER_81_920 ();
 FILLCELL_X1 FILLER_81_922 ();
 FILLCELL_X2 FILLER_81_947 ();
 FILLCELL_X1 FILLER_81_968 ();
 FILLCELL_X1 FILLER_81_992 ();
 FILLCELL_X4 FILLER_81_1011 ();
 FILLCELL_X1 FILLER_81_1015 ();
 FILLCELL_X32 FILLER_81_1019 ();
 FILLCELL_X16 FILLER_81_1051 ();
 FILLCELL_X2 FILLER_81_1067 ();
 FILLCELL_X8 FILLER_81_1100 ();
 FILLCELL_X4 FILLER_81_1108 ();
 FILLCELL_X2 FILLER_81_1112 ();
 FILLCELL_X1 FILLER_81_1126 ();
 FILLCELL_X2 FILLER_81_1134 ();
 FILLCELL_X16 FILLER_81_1170 ();
 FILLCELL_X8 FILLER_81_1186 ();
 FILLCELL_X4 FILLER_81_1194 ();
 FILLCELL_X2 FILLER_81_1238 ();
 FILLCELL_X8 FILLER_82_1 ();
 FILLCELL_X4 FILLER_82_9 ();
 FILLCELL_X1 FILLER_82_13 ();
 FILLCELL_X32 FILLER_82_17 ();
 FILLCELL_X8 FILLER_82_87 ();
 FILLCELL_X1 FILLER_82_95 ();
 FILLCELL_X8 FILLER_82_113 ();
 FILLCELL_X4 FILLER_82_121 ();
 FILLCELL_X2 FILLER_82_125 ();
 FILLCELL_X4 FILLER_82_151 ();
 FILLCELL_X2 FILLER_82_155 ();
 FILLCELL_X4 FILLER_82_164 ();
 FILLCELL_X2 FILLER_82_168 ();
 FILLCELL_X1 FILLER_82_170 ();
 FILLCELL_X1 FILLER_82_195 ();
 FILLCELL_X2 FILLER_82_203 ();
 FILLCELL_X1 FILLER_82_218 ();
 FILLCELL_X2 FILLER_82_226 ();
 FILLCELL_X8 FILLER_82_231 ();
 FILLCELL_X4 FILLER_82_239 ();
 FILLCELL_X1 FILLER_82_243 ();
 FILLCELL_X16 FILLER_82_251 ();
 FILLCELL_X8 FILLER_82_267 ();
 FILLCELL_X1 FILLER_82_275 ();
 FILLCELL_X4 FILLER_82_280 ();
 FILLCELL_X8 FILLER_82_308 ();
 FILLCELL_X4 FILLER_82_316 ();
 FILLCELL_X2 FILLER_82_320 ();
 FILLCELL_X1 FILLER_82_322 ();
 FILLCELL_X8 FILLER_82_340 ();
 FILLCELL_X4 FILLER_82_348 ();
 FILLCELL_X8 FILLER_82_376 ();
 FILLCELL_X1 FILLER_82_384 ();
 FILLCELL_X1 FILLER_82_402 ();
 FILLCELL_X2 FILLER_82_410 ();
 FILLCELL_X1 FILLER_82_412 ();
 FILLCELL_X4 FILLER_82_430 ();
 FILLCELL_X4 FILLER_82_441 ();
 FILLCELL_X1 FILLER_82_445 ();
 FILLCELL_X4 FILLER_82_509 ();
 FILLCELL_X4 FILLER_82_521 ();
 FILLCELL_X2 FILLER_82_525 ();
 FILLCELL_X1 FILLER_82_539 ();
 FILLCELL_X2 FILLER_82_544 ();
 FILLCELL_X4 FILLER_82_567 ();
 FILLCELL_X2 FILLER_82_571 ();
 FILLCELL_X1 FILLER_82_573 ();
 FILLCELL_X2 FILLER_82_598 ();
 FILLCELL_X1 FILLER_82_607 ();
 FILLCELL_X4 FILLER_82_615 ();
 FILLCELL_X16 FILLER_82_649 ();
 FILLCELL_X8 FILLER_82_665 ();
 FILLCELL_X4 FILLER_82_673 ();
 FILLCELL_X2 FILLER_82_677 ();
 FILLCELL_X2 FILLER_82_713 ();
 FILLCELL_X4 FILLER_82_732 ();
 FILLCELL_X1 FILLER_82_736 ();
 FILLCELL_X16 FILLER_82_761 ();
 FILLCELL_X1 FILLER_82_777 ();
 FILLCELL_X4 FILLER_82_809 ();
 FILLCELL_X2 FILLER_82_813 ();
 FILLCELL_X1 FILLER_82_824 ();
 FILLCELL_X1 FILLER_82_839 ();
 FILLCELL_X1 FILLER_82_850 ();
 FILLCELL_X2 FILLER_82_869 ();
 FILLCELL_X1 FILLER_82_885 ();
 FILLCELL_X8 FILLER_82_923 ();
 FILLCELL_X1 FILLER_82_931 ();
 FILLCELL_X2 FILLER_82_940 ();
 FILLCELL_X2 FILLER_82_956 ();
 FILLCELL_X1 FILLER_82_992 ();
 FILLCELL_X32 FILLER_82_996 ();
 FILLCELL_X2 FILLER_82_1028 ();
 FILLCELL_X16 FILLER_82_1037 ();
 FILLCELL_X4 FILLER_82_1053 ();
 FILLCELL_X1 FILLER_82_1057 ();
 FILLCELL_X32 FILLER_82_1071 ();
 FILLCELL_X8 FILLER_82_1103 ();
 FILLCELL_X4 FILLER_82_1111 ();
 FILLCELL_X2 FILLER_82_1115 ();
 FILLCELL_X1 FILLER_82_1117 ();
 FILLCELL_X4 FILLER_82_1131 ();
 FILLCELL_X8 FILLER_82_1139 ();
 FILLCELL_X4 FILLER_82_1147 ();
 FILLCELL_X1 FILLER_82_1188 ();
 FILLCELL_X2 FILLER_82_1192 ();
 FILLCELL_X1 FILLER_82_1211 ();
 FILLCELL_X1 FILLER_82_1215 ();
 FILLCELL_X1 FILLER_82_1223 ();
 FILLCELL_X4 FILLER_82_1234 ();
 FILLCELL_X2 FILLER_82_1238 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X4 FILLER_83_33 ();
 FILLCELL_X1 FILLER_83_37 ();
 FILLCELL_X1 FILLER_83_62 ();
 FILLCELL_X8 FILLER_83_80 ();
 FILLCELL_X4 FILLER_83_88 ();
 FILLCELL_X2 FILLER_83_92 ();
 FILLCELL_X8 FILLER_83_108 ();
 FILLCELL_X2 FILLER_83_120 ();
 FILLCELL_X4 FILLER_83_136 ();
 FILLCELL_X1 FILLER_83_140 ();
 FILLCELL_X2 FILLER_83_148 ();
 FILLCELL_X1 FILLER_83_150 ();
 FILLCELL_X4 FILLER_83_158 ();
 FILLCELL_X8 FILLER_83_169 ();
 FILLCELL_X1 FILLER_83_190 ();
 FILLCELL_X1 FILLER_83_198 ();
 FILLCELL_X1 FILLER_83_223 ();
 FILLCELL_X1 FILLER_83_241 ();
 FILLCELL_X2 FILLER_83_249 ();
 FILLCELL_X2 FILLER_83_272 ();
 FILLCELL_X16 FILLER_83_283 ();
 FILLCELL_X8 FILLER_83_299 ();
 FILLCELL_X4 FILLER_83_307 ();
 FILLCELL_X1 FILLER_83_311 ();
 FILLCELL_X2 FILLER_83_319 ();
 FILLCELL_X1 FILLER_83_328 ();
 FILLCELL_X2 FILLER_83_336 ();
 FILLCELL_X1 FILLER_83_338 ();
 FILLCELL_X2 FILLER_83_360 ();
 FILLCELL_X1 FILLER_83_362 ();
 FILLCELL_X8 FILLER_83_370 ();
 FILLCELL_X4 FILLER_83_378 ();
 FILLCELL_X1 FILLER_83_382 ();
 FILLCELL_X2 FILLER_83_400 ();
 FILLCELL_X1 FILLER_83_402 ();
 FILLCELL_X4 FILLER_83_410 ();
 FILLCELL_X16 FILLER_83_452 ();
 FILLCELL_X8 FILLER_83_468 ();
 FILLCELL_X4 FILLER_83_476 ();
 FILLCELL_X2 FILLER_83_480 ();
 FILLCELL_X1 FILLER_83_482 ();
 FILLCELL_X16 FILLER_83_490 ();
 FILLCELL_X2 FILLER_83_506 ();
 FILLCELL_X1 FILLER_83_522 ();
 FILLCELL_X4 FILLER_83_528 ();
 FILLCELL_X8 FILLER_83_549 ();
 FILLCELL_X1 FILLER_83_557 ();
 FILLCELL_X32 FILLER_83_565 ();
 FILLCELL_X4 FILLER_83_597 ();
 FILLCELL_X32 FILLER_83_618 ();
 FILLCELL_X16 FILLER_83_650 ();
 FILLCELL_X4 FILLER_83_666 ();
 FILLCELL_X4 FILLER_83_687 ();
 FILLCELL_X16 FILLER_83_729 ();
 FILLCELL_X8 FILLER_83_755 ();
 FILLCELL_X4 FILLER_83_763 ();
 FILLCELL_X2 FILLER_83_767 ();
 FILLCELL_X1 FILLER_83_769 ();
 FILLCELL_X1 FILLER_83_787 ();
 FILLCELL_X4 FILLER_83_812 ();
 FILLCELL_X2 FILLER_83_816 ();
 FILLCELL_X1 FILLER_83_818 ();
 FILLCELL_X2 FILLER_83_828 ();
 FILLCELL_X4 FILLER_83_853 ();
 FILLCELL_X2 FILLER_83_871 ();
 FILLCELL_X1 FILLER_83_873 ();
 FILLCELL_X2 FILLER_83_890 ();
 FILLCELL_X1 FILLER_83_901 ();
 FILLCELL_X2 FILLER_83_927 ();
 FILLCELL_X8 FILLER_83_943 ();
 FILLCELL_X2 FILLER_83_951 ();
 FILLCELL_X8 FILLER_83_992 ();
 FILLCELL_X4 FILLER_83_1000 ();
 FILLCELL_X1 FILLER_83_1021 ();
 FILLCELL_X2 FILLER_83_1029 ();
 FILLCELL_X8 FILLER_83_1048 ();
 FILLCELL_X1 FILLER_83_1056 ();
 FILLCELL_X8 FILLER_83_1068 ();
 FILLCELL_X1 FILLER_83_1076 ();
 FILLCELL_X4 FILLER_83_1084 ();
 FILLCELL_X2 FILLER_83_1088 ();
 FILLCELL_X1 FILLER_83_1090 ();
 FILLCELL_X8 FILLER_83_1098 ();
 FILLCELL_X4 FILLER_83_1106 ();
 FILLCELL_X2 FILLER_83_1110 ();
 FILLCELL_X1 FILLER_83_1112 ();
 FILLCELL_X32 FILLER_83_1120 ();
 FILLCELL_X2 FILLER_83_1172 ();
 FILLCELL_X16 FILLER_83_1178 ();
 FILLCELL_X2 FILLER_83_1194 ();
 FILLCELL_X1 FILLER_83_1206 ();
 FILLCELL_X4 FILLER_83_1214 ();
 FILLCELL_X1 FILLER_83_1224 ();
 FILLCELL_X4 FILLER_83_1235 ();
 FILLCELL_X1 FILLER_83_1239 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X8 FILLER_84_33 ();
 FILLCELL_X2 FILLER_84_41 ();
 FILLCELL_X2 FILLER_84_60 ();
 FILLCELL_X1 FILLER_84_62 ();
 FILLCELL_X4 FILLER_84_70 ();
 FILLCELL_X1 FILLER_84_74 ();
 FILLCELL_X8 FILLER_84_82 ();
 FILLCELL_X1 FILLER_84_90 ();
 FILLCELL_X8 FILLER_84_108 ();
 FILLCELL_X1 FILLER_84_116 ();
 FILLCELL_X4 FILLER_84_134 ();
 FILLCELL_X2 FILLER_84_138 ();
 FILLCELL_X32 FILLER_84_157 ();
 FILLCELL_X32 FILLER_84_189 ();
 FILLCELL_X8 FILLER_84_221 ();
 FILLCELL_X4 FILLER_84_229 ();
 FILLCELL_X1 FILLER_84_233 ();
 FILLCELL_X4 FILLER_84_275 ();
 FILLCELL_X1 FILLER_84_279 ();
 FILLCELL_X16 FILLER_84_294 ();
 FILLCELL_X2 FILLER_84_310 ();
 FILLCELL_X8 FILLER_84_343 ();
 FILLCELL_X4 FILLER_84_351 ();
 FILLCELL_X8 FILLER_84_372 ();
 FILLCELL_X4 FILLER_84_380 ();
 FILLCELL_X2 FILLER_84_384 ();
 FILLCELL_X8 FILLER_84_410 ();
 FILLCELL_X4 FILLER_84_423 ();
 FILLCELL_X1 FILLER_84_427 ();
 FILLCELL_X4 FILLER_84_433 ();
 FILLCELL_X32 FILLER_84_444 ();
 FILLCELL_X4 FILLER_84_476 ();
 FILLCELL_X4 FILLER_84_492 ();
 FILLCELL_X2 FILLER_84_496 ();
 FILLCELL_X2 FILLER_84_504 ();
 FILLCELL_X1 FILLER_84_506 ();
 FILLCELL_X8 FILLER_84_528 ();
 FILLCELL_X4 FILLER_84_550 ();
 FILLCELL_X2 FILLER_84_554 ();
 FILLCELL_X8 FILLER_84_573 ();
 FILLCELL_X2 FILLER_84_619 ();
 FILLCELL_X1 FILLER_84_621 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_639 ();
 FILLCELL_X4 FILLER_84_671 ();
 FILLCELL_X8 FILLER_84_682 ();
 FILLCELL_X4 FILLER_84_690 ();
 FILLCELL_X1 FILLER_84_694 ();
 FILLCELL_X16 FILLER_84_719 ();
 FILLCELL_X4 FILLER_84_742 ();
 FILLCELL_X1 FILLER_84_746 ();
 FILLCELL_X1 FILLER_84_754 ();
 FILLCELL_X4 FILLER_84_786 ();
 FILLCELL_X8 FILLER_84_800 ();
 FILLCELL_X4 FILLER_84_808 ();
 FILLCELL_X2 FILLER_84_812 ();
 FILLCELL_X8 FILLER_84_849 ();
 FILLCELL_X1 FILLER_84_866 ();
 FILLCELL_X4 FILLER_84_890 ();
 FILLCELL_X1 FILLER_84_901 ();
 FILLCELL_X2 FILLER_84_929 ();
 FILLCELL_X2 FILLER_84_941 ();
 FILLCELL_X4 FILLER_84_948 ();
 FILLCELL_X2 FILLER_84_952 ();
 FILLCELL_X1 FILLER_84_981 ();
 FILLCELL_X8 FILLER_84_987 ();
 FILLCELL_X4 FILLER_84_995 ();
 FILLCELL_X2 FILLER_84_999 ();
 FILLCELL_X1 FILLER_84_1001 ();
 FILLCELL_X4 FILLER_84_1081 ();
 FILLCELL_X4 FILLER_84_1102 ();
 FILLCELL_X4 FILLER_84_1126 ();
 FILLCELL_X2 FILLER_84_1130 ();
 FILLCELL_X1 FILLER_84_1132 ();
 FILLCELL_X8 FILLER_84_1150 ();
 FILLCELL_X4 FILLER_84_1158 ();
 FILLCELL_X2 FILLER_84_1183 ();
 FILLCELL_X1 FILLER_84_1185 ();
 FILLCELL_X2 FILLER_84_1223 ();
 FILLCELL_X1 FILLER_84_1239 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X16 FILLER_85_97 ();
 FILLCELL_X1 FILLER_85_113 ();
 FILLCELL_X32 FILLER_85_117 ();
 FILLCELL_X16 FILLER_85_149 ();
 FILLCELL_X2 FILLER_85_165 ();
 FILLCELL_X8 FILLER_85_174 ();
 FILLCELL_X1 FILLER_85_182 ();
 FILLCELL_X1 FILLER_85_189 ();
 FILLCELL_X4 FILLER_85_197 ();
 FILLCELL_X1 FILLER_85_201 ();
 FILLCELL_X8 FILLER_85_217 ();
 FILLCELL_X2 FILLER_85_238 ();
 FILLCELL_X1 FILLER_85_240 ();
 FILLCELL_X8 FILLER_85_265 ();
 FILLCELL_X4 FILLER_85_273 ();
 FILLCELL_X2 FILLER_85_277 ();
 FILLCELL_X1 FILLER_85_279 ();
 FILLCELL_X2 FILLER_85_297 ();
 FILLCELL_X1 FILLER_85_316 ();
 FILLCELL_X2 FILLER_85_334 ();
 FILLCELL_X32 FILLER_85_343 ();
 FILLCELL_X8 FILLER_85_375 ();
 FILLCELL_X4 FILLER_85_383 ();
 FILLCELL_X2 FILLER_85_387 ();
 FILLCELL_X4 FILLER_85_413 ();
 FILLCELL_X2 FILLER_85_417 ();
 FILLCELL_X1 FILLER_85_419 ();
 FILLCELL_X4 FILLER_85_427 ();
 FILLCELL_X2 FILLER_85_431 ();
 FILLCELL_X2 FILLER_85_450 ();
 FILLCELL_X4 FILLER_85_459 ();
 FILLCELL_X2 FILLER_85_480 ();
 FILLCELL_X1 FILLER_85_506 ();
 FILLCELL_X4 FILLER_85_533 ();
 FILLCELL_X16 FILLER_85_594 ();
 FILLCELL_X8 FILLER_85_610 ();
 FILLCELL_X1 FILLER_85_625 ();
 FILLCELL_X2 FILLER_85_633 ();
 FILLCELL_X1 FILLER_85_652 ();
 FILLCELL_X1 FILLER_85_670 ();
 FILLCELL_X4 FILLER_85_685 ();
 FILLCELL_X1 FILLER_85_689 ();
 FILLCELL_X2 FILLER_85_694 ();
 FILLCELL_X1 FILLER_85_696 ();
 FILLCELL_X8 FILLER_85_710 ();
 FILLCELL_X4 FILLER_85_718 ();
 FILLCELL_X1 FILLER_85_722 ();
 FILLCELL_X4 FILLER_85_730 ();
 FILLCELL_X1 FILLER_85_734 ();
 FILLCELL_X1 FILLER_85_752 ();
 FILLCELL_X1 FILLER_85_760 ();
 FILLCELL_X2 FILLER_85_787 ();
 FILLCELL_X16 FILLER_85_799 ();
 FILLCELL_X1 FILLER_85_815 ();
 FILLCELL_X8 FILLER_85_847 ();
 FILLCELL_X2 FILLER_85_872 ();
 FILLCELL_X1 FILLER_85_874 ();
 FILLCELL_X2 FILLER_85_883 ();
 FILLCELL_X2 FILLER_85_890 ();
 FILLCELL_X1 FILLER_85_892 ();
 FILLCELL_X1 FILLER_85_903 ();
 FILLCELL_X2 FILLER_85_907 ();
 FILLCELL_X1 FILLER_85_909 ();
 FILLCELL_X2 FILLER_85_953 ();
 FILLCELL_X1 FILLER_85_955 ();
 FILLCELL_X1 FILLER_85_963 ();
 FILLCELL_X4 FILLER_85_971 ();
 FILLCELL_X2 FILLER_85_975 ();
 FILLCELL_X1 FILLER_85_977 ();
 FILLCELL_X16 FILLER_85_992 ();
 FILLCELL_X8 FILLER_85_1063 ();
 FILLCELL_X2 FILLER_85_1071 ();
 FILLCELL_X1 FILLER_85_1073 ();
 FILLCELL_X4 FILLER_85_1094 ();
 FILLCELL_X1 FILLER_85_1098 ();
 FILLCELL_X1 FILLER_85_1169 ();
 FILLCELL_X4 FILLER_85_1187 ();
 FILLCELL_X2 FILLER_85_1191 ();
 FILLCELL_X1 FILLER_85_1193 ();
 FILLCELL_X4 FILLER_85_1201 ();
 FILLCELL_X1 FILLER_85_1205 ();
 FILLCELL_X1 FILLER_85_1222 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X8 FILLER_86_33 ();
 FILLCELL_X2 FILLER_86_41 ();
 FILLCELL_X16 FILLER_86_69 ();
 FILLCELL_X2 FILLER_86_85 ();
 FILLCELL_X1 FILLER_86_87 ();
 FILLCELL_X2 FILLER_86_105 ();
 FILLCELL_X1 FILLER_86_119 ();
 FILLCELL_X1 FILLER_86_134 ();
 FILLCELL_X2 FILLER_86_169 ();
 FILLCELL_X1 FILLER_86_171 ();
 FILLCELL_X1 FILLER_86_189 ();
 FILLCELL_X1 FILLER_86_204 ();
 FILLCELL_X16 FILLER_86_227 ();
 FILLCELL_X8 FILLER_86_243 ();
 FILLCELL_X4 FILLER_86_251 ();
 FILLCELL_X2 FILLER_86_255 ();
 FILLCELL_X1 FILLER_86_257 ();
 FILLCELL_X1 FILLER_86_265 ();
 FILLCELL_X32 FILLER_86_301 ();
 FILLCELL_X8 FILLER_86_333 ();
 FILLCELL_X4 FILLER_86_341 ();
 FILLCELL_X1 FILLER_86_345 ();
 FILLCELL_X2 FILLER_86_353 ();
 FILLCELL_X1 FILLER_86_379 ();
 FILLCELL_X16 FILLER_86_391 ();
 FILLCELL_X8 FILLER_86_407 ();
 FILLCELL_X4 FILLER_86_415 ();
 FILLCELL_X2 FILLER_86_419 ();
 FILLCELL_X2 FILLER_86_427 ();
 FILLCELL_X1 FILLER_86_429 ();
 FILLCELL_X1 FILLER_86_459 ();
 FILLCELL_X1 FILLER_86_517 ();
 FILLCELL_X4 FILLER_86_527 ();
 FILLCELL_X16 FILLER_86_561 ();
 FILLCELL_X4 FILLER_86_577 ();
 FILLCELL_X4 FILLER_86_584 ();
 FILLCELL_X1 FILLER_86_588 ();
 FILLCELL_X8 FILLER_86_613 ();
 FILLCELL_X2 FILLER_86_621 ();
 FILLCELL_X1 FILLER_86_623 ();
 FILLCELL_X8 FILLER_86_649 ();
 FILLCELL_X4 FILLER_86_657 ();
 FILLCELL_X32 FILLER_86_697 ();
 FILLCELL_X8 FILLER_86_729 ();
 FILLCELL_X1 FILLER_86_737 ();
 FILLCELL_X8 FILLER_86_749 ();
 FILLCELL_X16 FILLER_86_770 ();
 FILLCELL_X2 FILLER_86_786 ();
 FILLCELL_X8 FILLER_86_806 ();
 FILLCELL_X2 FILLER_86_814 ();
 FILLCELL_X1 FILLER_86_816 ();
 FILLCELL_X4 FILLER_86_820 ();
 FILLCELL_X1 FILLER_86_824 ();
 FILLCELL_X2 FILLER_86_835 ();
 FILLCELL_X2 FILLER_86_841 ();
 FILLCELL_X1 FILLER_86_843 ();
 FILLCELL_X2 FILLER_86_849 ();
 FILLCELL_X2 FILLER_86_856 ();
 FILLCELL_X1 FILLER_86_858 ();
 FILLCELL_X1 FILLER_86_864 ();
 FILLCELL_X2 FILLER_86_870 ();
 FILLCELL_X1 FILLER_86_872 ();
 FILLCELL_X1 FILLER_86_892 ();
 FILLCELL_X1 FILLER_86_896 ();
 FILLCELL_X2 FILLER_86_911 ();
 FILLCELL_X2 FILLER_86_916 ();
 FILLCELL_X2 FILLER_86_921 ();
 FILLCELL_X1 FILLER_86_923 ();
 FILLCELL_X1 FILLER_86_941 ();
 FILLCELL_X4 FILLER_86_949 ();
 FILLCELL_X1 FILLER_86_953 ();
 FILLCELL_X1 FILLER_86_957 ();
 FILLCELL_X8 FILLER_86_971 ();
 FILLCELL_X2 FILLER_86_979 ();
 FILLCELL_X1 FILLER_86_981 ();
 FILLCELL_X8 FILLER_86_985 ();
 FILLCELL_X1 FILLER_86_993 ();
 FILLCELL_X32 FILLER_86_1001 ();
 FILLCELL_X8 FILLER_86_1033 ();
 FILLCELL_X2 FILLER_86_1041 ();
 FILLCELL_X8 FILLER_86_1065 ();
 FILLCELL_X4 FILLER_86_1073 ();
 FILLCELL_X1 FILLER_86_1077 ();
 FILLCELL_X4 FILLER_86_1103 ();
 FILLCELL_X2 FILLER_86_1107 ();
 FILLCELL_X2 FILLER_86_1123 ();
 FILLCELL_X1 FILLER_86_1125 ();
 FILLCELL_X16 FILLER_86_1140 ();
 FILLCELL_X8 FILLER_86_1156 ();
 FILLCELL_X2 FILLER_86_1164 ();
 FILLCELL_X1 FILLER_86_1166 ();
 FILLCELL_X8 FILLER_86_1171 ();
 FILLCELL_X4 FILLER_86_1179 ();
 FILLCELL_X2 FILLER_86_1183 ();
 FILLCELL_X1 FILLER_86_1185 ();
 FILLCELL_X8 FILLER_86_1193 ();
 FILLCELL_X4 FILLER_86_1201 ();
 FILLCELL_X2 FILLER_86_1205 ();
 FILLCELL_X2 FILLER_86_1238 ();
 FILLCELL_X8 FILLER_87_1 ();
 FILLCELL_X4 FILLER_87_9 ();
 FILLCELL_X1 FILLER_87_13 ();
 FILLCELL_X16 FILLER_87_17 ();
 FILLCELL_X8 FILLER_87_33 ();
 FILLCELL_X2 FILLER_87_41 ();
 FILLCELL_X1 FILLER_87_70 ();
 FILLCELL_X2 FILLER_87_78 ();
 FILLCELL_X2 FILLER_87_98 ();
 FILLCELL_X4 FILLER_87_107 ();
 FILLCELL_X2 FILLER_87_169 ();
 FILLCELL_X4 FILLER_87_226 ();
 FILLCELL_X16 FILLER_87_237 ();
 FILLCELL_X1 FILLER_87_253 ();
 FILLCELL_X8 FILLER_87_261 ();
 FILLCELL_X4 FILLER_87_269 ();
 FILLCELL_X2 FILLER_87_273 ();
 FILLCELL_X1 FILLER_87_275 ();
 FILLCELL_X4 FILLER_87_283 ();
 FILLCELL_X1 FILLER_87_287 ();
 FILLCELL_X32 FILLER_87_295 ();
 FILLCELL_X4 FILLER_87_327 ();
 FILLCELL_X2 FILLER_87_331 ();
 FILLCELL_X1 FILLER_87_333 ();
 FILLCELL_X4 FILLER_87_341 ();
 FILLCELL_X1 FILLER_87_393 ();
 FILLCELL_X8 FILLER_87_401 ();
 FILLCELL_X4 FILLER_87_409 ();
 FILLCELL_X16 FILLER_87_437 ();
 FILLCELL_X8 FILLER_87_453 ();
 FILLCELL_X2 FILLER_87_461 ();
 FILLCELL_X1 FILLER_87_463 ();
 FILLCELL_X8 FILLER_87_481 ();
 FILLCELL_X2 FILLER_87_489 ();
 FILLCELL_X1 FILLER_87_491 ();
 FILLCELL_X1 FILLER_87_499 ();
 FILLCELL_X2 FILLER_87_504 ();
 FILLCELL_X1 FILLER_87_512 ();
 FILLCELL_X1 FILLER_87_530 ();
 FILLCELL_X2 FILLER_87_542 ();
 FILLCELL_X4 FILLER_87_547 ();
 FILLCELL_X16 FILLER_87_574 ();
 FILLCELL_X4 FILLER_87_590 ();
 FILLCELL_X2 FILLER_87_594 ();
 FILLCELL_X1 FILLER_87_596 ();
 FILLCELL_X32 FILLER_87_614 ();
 FILLCELL_X16 FILLER_87_646 ();
 FILLCELL_X4 FILLER_87_662 ();
 FILLCELL_X4 FILLER_87_690 ();
 FILLCELL_X1 FILLER_87_694 ();
 FILLCELL_X4 FILLER_87_719 ();
 FILLCELL_X4 FILLER_87_747 ();
 FILLCELL_X1 FILLER_87_751 ();
 FILLCELL_X16 FILLER_87_774 ();
 FILLCELL_X16 FILLER_87_800 ();
 FILLCELL_X1 FILLER_87_816 ();
 FILLCELL_X1 FILLER_87_878 ();
 FILLCELL_X4 FILLER_87_900 ();
 FILLCELL_X2 FILLER_87_904 ();
 FILLCELL_X1 FILLER_87_906 ();
 FILLCELL_X4 FILLER_87_921 ();
 FILLCELL_X1 FILLER_87_932 ();
 FILLCELL_X4 FILLER_87_940 ();
 FILLCELL_X2 FILLER_87_944 ();
 FILLCELL_X1 FILLER_87_946 ();
 FILLCELL_X4 FILLER_87_969 ();
 FILLCELL_X4 FILLER_87_985 ();
 FILLCELL_X1 FILLER_87_989 ();
 FILLCELL_X8 FILLER_87_1014 ();
 FILLCELL_X2 FILLER_87_1022 ();
 FILLCELL_X16 FILLER_87_1044 ();
 FILLCELL_X8 FILLER_87_1060 ();
 FILLCELL_X4 FILLER_87_1068 ();
 FILLCELL_X2 FILLER_87_1072 ();
 FILLCELL_X8 FILLER_87_1077 ();
 FILLCELL_X2 FILLER_87_1085 ();
 FILLCELL_X16 FILLER_87_1098 ();
 FILLCELL_X4 FILLER_87_1114 ();
 FILLCELL_X1 FILLER_87_1118 ();
 FILLCELL_X16 FILLER_87_1128 ();
 FILLCELL_X4 FILLER_87_1144 ();
 FILLCELL_X2 FILLER_87_1148 ();
 FILLCELL_X8 FILLER_87_1179 ();
 FILLCELL_X1 FILLER_87_1204 ();
 FILLCELL_X2 FILLER_87_1234 ();
 FILLCELL_X1 FILLER_87_1236 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X8 FILLER_88_33 ();
 FILLCELL_X1 FILLER_88_41 ();
 FILLCELL_X8 FILLER_88_83 ();
 FILLCELL_X2 FILLER_88_91 ();
 FILLCELL_X2 FILLER_88_100 ();
 FILLCELL_X1 FILLER_88_119 ();
 FILLCELL_X1 FILLER_88_127 ();
 FILLCELL_X2 FILLER_88_135 ();
 FILLCELL_X2 FILLER_88_144 ();
 FILLCELL_X2 FILLER_88_153 ();
 FILLCELL_X1 FILLER_88_155 ();
 FILLCELL_X16 FILLER_88_170 ();
 FILLCELL_X2 FILLER_88_186 ();
 FILLCELL_X4 FILLER_88_195 ();
 FILLCELL_X8 FILLER_88_213 ();
 FILLCELL_X1 FILLER_88_221 ();
 FILLCELL_X8 FILLER_88_250 ();
 FILLCELL_X4 FILLER_88_258 ();
 FILLCELL_X1 FILLER_88_262 ();
 FILLCELL_X2 FILLER_88_270 ();
 FILLCELL_X1 FILLER_88_272 ();
 FILLCELL_X4 FILLER_88_290 ();
 FILLCELL_X4 FILLER_88_327 ();
 FILLCELL_X1 FILLER_88_331 ();
 FILLCELL_X4 FILLER_88_340 ();
 FILLCELL_X1 FILLER_88_344 ();
 FILLCELL_X8 FILLER_88_352 ();
 FILLCELL_X16 FILLER_88_391 ();
 FILLCELL_X4 FILLER_88_407 ();
 FILLCELL_X2 FILLER_88_411 ();
 FILLCELL_X1 FILLER_88_413 ();
 FILLCELL_X4 FILLER_88_431 ();
 FILLCELL_X1 FILLER_88_435 ();
 FILLCELL_X2 FILLER_88_460 ();
 FILLCELL_X1 FILLER_88_462 ();
 FILLCELL_X4 FILLER_88_470 ();
 FILLCELL_X2 FILLER_88_474 ();
 FILLCELL_X1 FILLER_88_476 ();
 FILLCELL_X2 FILLER_88_484 ();
 FILLCELL_X16 FILLER_88_493 ();
 FILLCELL_X8 FILLER_88_548 ();
 FILLCELL_X16 FILLER_88_570 ();
 FILLCELL_X8 FILLER_88_586 ();
 FILLCELL_X4 FILLER_88_594 ();
 FILLCELL_X1 FILLER_88_598 ();
 FILLCELL_X16 FILLER_88_613 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X16 FILLER_88_664 ();
 FILLCELL_X8 FILLER_88_680 ();
 FILLCELL_X4 FILLER_88_688 ();
 FILLCELL_X2 FILLER_88_692 ();
 FILLCELL_X2 FILLER_88_718 ();
 FILLCELL_X1 FILLER_88_720 ();
 FILLCELL_X4 FILLER_88_731 ();
 FILLCELL_X2 FILLER_88_735 ();
 FILLCELL_X2 FILLER_88_755 ();
 FILLCELL_X1 FILLER_88_757 ();
 FILLCELL_X2 FILLER_88_771 ();
 FILLCELL_X1 FILLER_88_773 ();
 FILLCELL_X8 FILLER_88_808 ();
 FILLCELL_X4 FILLER_88_816 ();
 FILLCELL_X2 FILLER_88_823 ();
 FILLCELL_X1 FILLER_88_834 ();
 FILLCELL_X8 FILLER_88_845 ();
 FILLCELL_X4 FILLER_88_853 ();
 FILLCELL_X1 FILLER_88_857 ();
 FILLCELL_X2 FILLER_88_865 ();
 FILLCELL_X4 FILLER_88_871 ();
 FILLCELL_X2 FILLER_88_875 ();
 FILLCELL_X2 FILLER_88_892 ();
 FILLCELL_X2 FILLER_88_911 ();
 FILLCELL_X8 FILLER_88_936 ();
 FILLCELL_X2 FILLER_88_944 ();
 FILLCELL_X4 FILLER_88_974 ();
 FILLCELL_X2 FILLER_88_978 ();
 FILLCELL_X1 FILLER_88_980 ();
 FILLCELL_X1 FILLER_88_986 ();
 FILLCELL_X2 FILLER_88_1014 ();
 FILLCELL_X1 FILLER_88_1016 ();
 FILLCELL_X2 FILLER_88_1034 ();
 FILLCELL_X8 FILLER_88_1043 ();
 FILLCELL_X4 FILLER_88_1051 ();
 FILLCELL_X2 FILLER_88_1055 ();
 FILLCELL_X2 FILLER_88_1084 ();
 FILLCELL_X1 FILLER_88_1086 ();
 FILLCELL_X16 FILLER_88_1100 ();
 FILLCELL_X1 FILLER_88_1116 ();
 FILLCELL_X8 FILLER_88_1137 ();
 FILLCELL_X2 FILLER_88_1145 ();
 FILLCELL_X1 FILLER_88_1154 ();
 FILLCELL_X16 FILLER_88_1182 ();
 FILLCELL_X2 FILLER_88_1198 ();
 FILLCELL_X1 FILLER_88_1200 ();
 FILLCELL_X1 FILLER_88_1218 ();
 FILLCELL_X8 FILLER_88_1223 ();
 FILLCELL_X4 FILLER_88_1234 ();
 FILLCELL_X2 FILLER_88_1238 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X16 FILLER_89_33 ();
 FILLCELL_X8 FILLER_89_49 ();
 FILLCELL_X4 FILLER_89_57 ();
 FILLCELL_X1 FILLER_89_61 ();
 FILLCELL_X8 FILLER_89_79 ();
 FILLCELL_X4 FILLER_89_87 ();
 FILLCELL_X2 FILLER_89_91 ();
 FILLCELL_X32 FILLER_89_110 ();
 FILLCELL_X4 FILLER_89_149 ();
 FILLCELL_X1 FILLER_89_153 ();
 FILLCELL_X16 FILLER_89_161 ();
 FILLCELL_X8 FILLER_89_177 ();
 FILLCELL_X1 FILLER_89_185 ();
 FILLCELL_X2 FILLER_89_216 ();
 FILLCELL_X1 FILLER_89_218 ();
 FILLCELL_X8 FILLER_89_222 ();
 FILLCELL_X4 FILLER_89_230 ();
 FILLCELL_X2 FILLER_89_234 ();
 FILLCELL_X1 FILLER_89_236 ();
 FILLCELL_X2 FILLER_89_271 ();
 FILLCELL_X4 FILLER_89_280 ();
 FILLCELL_X1 FILLER_89_284 ();
 FILLCELL_X8 FILLER_89_297 ();
 FILLCELL_X8 FILLER_89_336 ();
 FILLCELL_X1 FILLER_89_344 ();
 FILLCELL_X8 FILLER_89_352 ();
 FILLCELL_X32 FILLER_89_367 ();
 FILLCELL_X8 FILLER_89_399 ();
 FILLCELL_X4 FILLER_89_407 ();
 FILLCELL_X1 FILLER_89_411 ();
 FILLCELL_X8 FILLER_89_426 ();
 FILLCELL_X2 FILLER_89_434 ();
 FILLCELL_X32 FILLER_89_443 ();
 FILLCELL_X8 FILLER_89_475 ();
 FILLCELL_X4 FILLER_89_483 ();
 FILLCELL_X2 FILLER_89_504 ();
 FILLCELL_X1 FILLER_89_506 ();
 FILLCELL_X2 FILLER_89_510 ();
 FILLCELL_X2 FILLER_89_518 ();
 FILLCELL_X8 FILLER_89_548 ();
 FILLCELL_X2 FILLER_89_556 ();
 FILLCELL_X1 FILLER_89_558 ();
 FILLCELL_X1 FILLER_89_566 ();
 FILLCELL_X16 FILLER_89_584 ();
 FILLCELL_X2 FILLER_89_600 ();
 FILLCELL_X1 FILLER_89_602 ();
 FILLCELL_X8 FILLER_89_619 ();
 FILLCELL_X4 FILLER_89_627 ();
 FILLCELL_X2 FILLER_89_631 ();
 FILLCELL_X1 FILLER_89_633 ();
 FILLCELL_X1 FILLER_89_661 ();
 FILLCELL_X4 FILLER_89_669 ();
 FILLCELL_X8 FILLER_89_690 ();
 FILLCELL_X2 FILLER_89_705 ();
 FILLCELL_X1 FILLER_89_707 ();
 FILLCELL_X1 FILLER_89_741 ();
 FILLCELL_X1 FILLER_89_762 ();
 FILLCELL_X2 FILLER_89_770 ();
 FILLCELL_X1 FILLER_89_772 ();
 FILLCELL_X1 FILLER_89_801 ();
 FILLCELL_X1 FILLER_89_806 ();
 FILLCELL_X2 FILLER_89_820 ();
 FILLCELL_X1 FILLER_89_829 ();
 FILLCELL_X1 FILLER_89_835 ();
 FILLCELL_X2 FILLER_89_840 ();
 FILLCELL_X1 FILLER_89_842 ();
 FILLCELL_X4 FILLER_89_848 ();
 FILLCELL_X2 FILLER_89_862 ();
 FILLCELL_X1 FILLER_89_899 ();
 FILLCELL_X1 FILLER_89_921 ();
 FILLCELL_X1 FILLER_89_935 ();
 FILLCELL_X2 FILLER_89_960 ();
 FILLCELL_X8 FILLER_89_983 ();
 FILLCELL_X4 FILLER_89_991 ();
 FILLCELL_X2 FILLER_89_995 ();
 FILLCELL_X1 FILLER_89_997 ();
 FILLCELL_X2 FILLER_89_1013 ();
 FILLCELL_X2 FILLER_89_1049 ();
 FILLCELL_X1 FILLER_89_1068 ();
 FILLCELL_X4 FILLER_89_1073 ();
 FILLCELL_X2 FILLER_89_1094 ();
 FILLCELL_X4 FILLER_89_1113 ();
 FILLCELL_X1 FILLER_89_1117 ();
 FILLCELL_X8 FILLER_89_1135 ();
 FILLCELL_X2 FILLER_89_1143 ();
 FILLCELL_X8 FILLER_89_1186 ();
 FILLCELL_X2 FILLER_89_1194 ();
 FILLCELL_X1 FILLER_89_1216 ();
 FILLCELL_X2 FILLER_89_1238 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X8 FILLER_90_65 ();
 FILLCELL_X4 FILLER_90_73 ();
 FILLCELL_X1 FILLER_90_77 ();
 FILLCELL_X16 FILLER_90_85 ();
 FILLCELL_X8 FILLER_90_101 ();
 FILLCELL_X4 FILLER_90_109 ();
 FILLCELL_X1 FILLER_90_113 ();
 FILLCELL_X16 FILLER_90_121 ();
 FILLCELL_X4 FILLER_90_137 ();
 FILLCELL_X1 FILLER_90_148 ();
 FILLCELL_X16 FILLER_90_156 ();
 FILLCELL_X8 FILLER_90_172 ();
 FILLCELL_X4 FILLER_90_180 ();
 FILLCELL_X16 FILLER_90_194 ();
 FILLCELL_X4 FILLER_90_217 ();
 FILLCELL_X2 FILLER_90_221 ();
 FILLCELL_X2 FILLER_90_254 ();
 FILLCELL_X4 FILLER_90_270 ();
 FILLCELL_X1 FILLER_90_274 ();
 FILLCELL_X1 FILLER_90_301 ();
 FILLCELL_X2 FILLER_90_316 ();
 FILLCELL_X1 FILLER_90_325 ();
 FILLCELL_X1 FILLER_90_333 ();
 FILLCELL_X32 FILLER_90_343 ();
 FILLCELL_X32 FILLER_90_375 ();
 FILLCELL_X2 FILLER_90_407 ();
 FILLCELL_X1 FILLER_90_420 ();
 FILLCELL_X1 FILLER_90_438 ();
 FILLCELL_X1 FILLER_90_463 ();
 FILLCELL_X2 FILLER_90_478 ();
 FILLCELL_X1 FILLER_90_480 ();
 FILLCELL_X4 FILLER_90_488 ();
 FILLCELL_X2 FILLER_90_492 ();
 FILLCELL_X1 FILLER_90_494 ();
 FILLCELL_X2 FILLER_90_527 ();
 FILLCELL_X1 FILLER_90_532 ();
 FILLCELL_X2 FILLER_90_542 ();
 FILLCELL_X4 FILLER_90_551 ();
 FILLCELL_X1 FILLER_90_555 ();
 FILLCELL_X4 FILLER_90_580 ();
 FILLCELL_X1 FILLER_90_584 ();
 FILLCELL_X8 FILLER_90_621 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X8 FILLER_90_632 ();
 FILLCELL_X1 FILLER_90_640 ();
 FILLCELL_X8 FILLER_90_670 ();
 FILLCELL_X2 FILLER_90_678 ();
 FILLCELL_X1 FILLER_90_680 ();
 FILLCELL_X8 FILLER_90_698 ();
 FILLCELL_X1 FILLER_90_706 ();
 FILLCELL_X8 FILLER_90_731 ();
 FILLCELL_X8 FILLER_90_744 ();
 FILLCELL_X4 FILLER_90_752 ();
 FILLCELL_X2 FILLER_90_756 ();
 FILLCELL_X4 FILLER_90_796 ();
 FILLCELL_X2 FILLER_90_800 ();
 FILLCELL_X8 FILLER_90_809 ();
 FILLCELL_X4 FILLER_90_817 ();
 FILLCELL_X1 FILLER_90_821 ();
 FILLCELL_X2 FILLER_90_839 ();
 FILLCELL_X1 FILLER_90_841 ();
 FILLCELL_X1 FILLER_90_852 ();
 FILLCELL_X1 FILLER_90_861 ();
 FILLCELL_X2 FILLER_90_876 ();
 FILLCELL_X1 FILLER_90_878 ();
 FILLCELL_X4 FILLER_90_886 ();
 FILLCELL_X2 FILLER_90_897 ();
 FILLCELL_X1 FILLER_90_973 ();
 FILLCELL_X8 FILLER_90_979 ();
 FILLCELL_X1 FILLER_90_987 ();
 FILLCELL_X2 FILLER_90_995 ();
 FILLCELL_X1 FILLER_90_997 ();
 FILLCELL_X16 FILLER_90_1002 ();
 FILLCELL_X4 FILLER_90_1018 ();
 FILLCELL_X2 FILLER_90_1022 ();
 FILLCELL_X1 FILLER_90_1038 ();
 FILLCELL_X1 FILLER_90_1046 ();
 FILLCELL_X1 FILLER_90_1071 ();
 FILLCELL_X2 FILLER_90_1079 ();
 FILLCELL_X1 FILLER_90_1126 ();
 FILLCELL_X2 FILLER_90_1134 ();
 FILLCELL_X2 FILLER_90_1157 ();
 FILLCELL_X8 FILLER_90_1166 ();
 FILLCELL_X2 FILLER_90_1174 ();
 FILLCELL_X8 FILLER_90_1183 ();
 FILLCELL_X4 FILLER_90_1191 ();
 FILLCELL_X1 FILLER_90_1195 ();
 FILLCELL_X1 FILLER_90_1218 ();
 FILLCELL_X1 FILLER_90_1239 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X16 FILLER_91_65 ();
 FILLCELL_X1 FILLER_91_81 ();
 FILLCELL_X8 FILLER_91_120 ();
 FILLCELL_X4 FILLER_91_128 ();
 FILLCELL_X2 FILLER_91_132 ();
 FILLCELL_X2 FILLER_91_158 ();
 FILLCELL_X1 FILLER_91_160 ();
 FILLCELL_X8 FILLER_91_223 ();
 FILLCELL_X4 FILLER_91_231 ();
 FILLCELL_X2 FILLER_91_242 ();
 FILLCELL_X1 FILLER_91_244 ();
 FILLCELL_X32 FILLER_91_262 ();
 FILLCELL_X8 FILLER_91_318 ();
 FILLCELL_X4 FILLER_91_326 ();
 FILLCELL_X1 FILLER_91_330 ();
 FILLCELL_X2 FILLER_91_362 ();
 FILLCELL_X1 FILLER_91_364 ();
 FILLCELL_X8 FILLER_91_382 ();
 FILLCELL_X1 FILLER_91_390 ();
 FILLCELL_X32 FILLER_91_408 ();
 FILLCELL_X16 FILLER_91_440 ();
 FILLCELL_X4 FILLER_91_456 ();
 FILLCELL_X1 FILLER_91_460 ();
 FILLCELL_X2 FILLER_91_468 ();
 FILLCELL_X2 FILLER_91_477 ();
 FILLCELL_X2 FILLER_91_513 ();
 FILLCELL_X8 FILLER_91_522 ();
 FILLCELL_X2 FILLER_91_530 ();
 FILLCELL_X2 FILLER_91_535 ();
 FILLCELL_X2 FILLER_91_555 ();
 FILLCELL_X1 FILLER_91_557 ();
 FILLCELL_X1 FILLER_91_565 ();
 FILLCELL_X16 FILLER_91_573 ();
 FILLCELL_X4 FILLER_91_589 ();
 FILLCELL_X1 FILLER_91_593 ();
 FILLCELL_X4 FILLER_91_632 ();
 FILLCELL_X1 FILLER_91_636 ();
 FILLCELL_X1 FILLER_91_699 ();
 FILLCELL_X2 FILLER_91_707 ();
 FILLCELL_X16 FILLER_91_733 ();
 FILLCELL_X8 FILLER_91_773 ();
 FILLCELL_X4 FILLER_91_781 ();
 FILLCELL_X2 FILLER_91_785 ();
 FILLCELL_X1 FILLER_91_787 ();
 FILLCELL_X16 FILLER_91_812 ();
 FILLCELL_X1 FILLER_91_828 ();
 FILLCELL_X2 FILLER_91_834 ();
 FILLCELL_X2 FILLER_91_856 ();
 FILLCELL_X2 FILLER_91_872 ();
 FILLCELL_X1 FILLER_91_874 ();
 FILLCELL_X2 FILLER_91_891 ();
 FILLCELL_X1 FILLER_91_893 ();
 FILLCELL_X4 FILLER_91_907 ();
 FILLCELL_X4 FILLER_91_916 ();
 FILLCELL_X1 FILLER_91_920 ();
 FILLCELL_X1 FILLER_91_924 ();
 FILLCELL_X1 FILLER_91_930 ();
 FILLCELL_X2 FILLER_91_942 ();
 FILLCELL_X2 FILLER_91_950 ();
 FILLCELL_X2 FILLER_91_956 ();
 FILLCELL_X4 FILLER_91_961 ();
 FILLCELL_X16 FILLER_91_972 ();
 FILLCELL_X8 FILLER_91_988 ();
 FILLCELL_X4 FILLER_91_996 ();
 FILLCELL_X2 FILLER_91_1000 ();
 FILLCELL_X1 FILLER_91_1009 ();
 FILLCELL_X8 FILLER_91_1013 ();
 FILLCELL_X4 FILLER_91_1021 ();
 FILLCELL_X1 FILLER_91_1025 ();
 FILLCELL_X8 FILLER_91_1042 ();
 FILLCELL_X1 FILLER_91_1050 ();
 FILLCELL_X16 FILLER_91_1058 ();
 FILLCELL_X4 FILLER_91_1074 ();
 FILLCELL_X2 FILLER_91_1109 ();
 FILLCELL_X1 FILLER_91_1111 ();
 FILLCELL_X4 FILLER_91_1117 ();
 FILLCELL_X2 FILLER_91_1121 ();
 FILLCELL_X1 FILLER_91_1123 ();
 FILLCELL_X4 FILLER_91_1131 ();
 FILLCELL_X1 FILLER_91_1135 ();
 FILLCELL_X8 FILLER_91_1150 ();
 FILLCELL_X1 FILLER_91_1158 ();
 FILLCELL_X16 FILLER_91_1176 ();
 FILLCELL_X8 FILLER_91_1192 ();
 FILLCELL_X1 FILLER_91_1200 ();
 FILLCELL_X1 FILLER_91_1236 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X4 FILLER_92_33 ();
 FILLCELL_X1 FILLER_92_37 ();
 FILLCELL_X2 FILLER_92_70 ();
 FILLCELL_X1 FILLER_92_72 ();
 FILLCELL_X4 FILLER_92_80 ();
 FILLCELL_X2 FILLER_92_84 ();
 FILLCELL_X8 FILLER_92_93 ();
 FILLCELL_X1 FILLER_92_101 ();
 FILLCELL_X4 FILLER_92_119 ();
 FILLCELL_X2 FILLER_92_123 ();
 FILLCELL_X1 FILLER_92_125 ();
 FILLCELL_X4 FILLER_92_133 ();
 FILLCELL_X1 FILLER_92_137 ();
 FILLCELL_X8 FILLER_92_155 ();
 FILLCELL_X4 FILLER_92_163 ();
 FILLCELL_X2 FILLER_92_167 ();
 FILLCELL_X2 FILLER_92_193 ();
 FILLCELL_X1 FILLER_92_195 ();
 FILLCELL_X1 FILLER_92_203 ();
 FILLCELL_X8 FILLER_92_221 ();
 FILLCELL_X4 FILLER_92_229 ();
 FILLCELL_X4 FILLER_92_240 ();
 FILLCELL_X32 FILLER_92_258 ();
 FILLCELL_X8 FILLER_92_290 ();
 FILLCELL_X4 FILLER_92_305 ();
 FILLCELL_X8 FILLER_92_316 ();
 FILLCELL_X1 FILLER_92_324 ();
 FILLCELL_X2 FILLER_92_332 ();
 FILLCELL_X4 FILLER_92_386 ();
 FILLCELL_X4 FILLER_92_397 ();
 FILLCELL_X2 FILLER_92_401 ();
 FILLCELL_X4 FILLER_92_410 ();
 FILLCELL_X16 FILLER_92_424 ();
 FILLCELL_X8 FILLER_92_440 ();
 FILLCELL_X4 FILLER_92_448 ();
 FILLCELL_X4 FILLER_92_476 ();
 FILLCELL_X1 FILLER_92_480 ();
 FILLCELL_X8 FILLER_92_498 ();
 FILLCELL_X1 FILLER_92_506 ();
 FILLCELL_X4 FILLER_92_514 ();
 FILLCELL_X1 FILLER_92_535 ();
 FILLCELL_X1 FILLER_92_543 ();
 FILLCELL_X2 FILLER_92_551 ();
 FILLCELL_X2 FILLER_92_557 ();
 FILLCELL_X2 FILLER_92_576 ();
 FILLCELL_X1 FILLER_92_578 ();
 FILLCELL_X2 FILLER_92_586 ();
 FILLCELL_X1 FILLER_92_588 ();
 FILLCELL_X2 FILLER_92_606 ();
 FILLCELL_X4 FILLER_92_615 ();
 FILLCELL_X2 FILLER_92_619 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X4 FILLER_92_632 ();
 FILLCELL_X2 FILLER_92_636 ();
 FILLCELL_X16 FILLER_92_662 ();
 FILLCELL_X4 FILLER_92_678 ();
 FILLCELL_X2 FILLER_92_682 ();
 FILLCELL_X16 FILLER_92_701 ();
 FILLCELL_X4 FILLER_92_717 ();
 FILLCELL_X2 FILLER_92_721 ();
 FILLCELL_X1 FILLER_92_723 ();
 FILLCELL_X16 FILLER_92_727 ();
 FILLCELL_X8 FILLER_92_743 ();
 FILLCELL_X2 FILLER_92_774 ();
 FILLCELL_X16 FILLER_92_810 ();
 FILLCELL_X8 FILLER_92_826 ();
 FILLCELL_X4 FILLER_92_834 ();
 FILLCELL_X2 FILLER_92_838 ();
 FILLCELL_X1 FILLER_92_872 ();
 FILLCELL_X4 FILLER_92_906 ();
 FILLCELL_X2 FILLER_92_910 ();
 FILLCELL_X1 FILLER_92_912 ();
 FILLCELL_X2 FILLER_92_951 ();
 FILLCELL_X2 FILLER_92_960 ();
 FILLCELL_X1 FILLER_92_962 ();
 FILLCELL_X2 FILLER_92_968 ();
 FILLCELL_X32 FILLER_92_977 ();
 FILLCELL_X16 FILLER_92_1009 ();
 FILLCELL_X4 FILLER_92_1025 ();
 FILLCELL_X2 FILLER_92_1029 ();
 FILLCELL_X32 FILLER_92_1034 ();
 FILLCELL_X8 FILLER_92_1066 ();
 FILLCELL_X4 FILLER_92_1074 ();
 FILLCELL_X2 FILLER_92_1078 ();
 FILLCELL_X1 FILLER_92_1080 ();
 FILLCELL_X2 FILLER_92_1094 ();
 FILLCELL_X16 FILLER_92_1113 ();
 FILLCELL_X8 FILLER_92_1129 ();
 FILLCELL_X32 FILLER_92_1161 ();
 FILLCELL_X8 FILLER_92_1193 ();
 FILLCELL_X2 FILLER_92_1201 ();
 FILLCELL_X1 FILLER_92_1203 ();
 FILLCELL_X8 FILLER_92_1213 ();
 FILLCELL_X1 FILLER_92_1221 ();
 FILLCELL_X2 FILLER_92_1225 ();
 FILLCELL_X1 FILLER_92_1227 ();
 FILLCELL_X2 FILLER_92_1231 ();
 FILLCELL_X1 FILLER_92_1233 ();
 FILLCELL_X2 FILLER_92_1237 ();
 FILLCELL_X1 FILLER_92_1239 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X4 FILLER_93_57 ();
 FILLCELL_X2 FILLER_93_61 ();
 FILLCELL_X8 FILLER_93_87 ();
 FILLCELL_X2 FILLER_93_95 ();
 FILLCELL_X1 FILLER_93_97 ();
 FILLCELL_X8 FILLER_93_102 ();
 FILLCELL_X4 FILLER_93_110 ();
 FILLCELL_X1 FILLER_93_114 ();
 FILLCELL_X2 FILLER_93_122 ();
 FILLCELL_X1 FILLER_93_124 ();
 FILLCELL_X32 FILLER_93_149 ();
 FILLCELL_X4 FILLER_93_181 ();
 FILLCELL_X1 FILLER_93_185 ();
 FILLCELL_X2 FILLER_93_193 ();
 FILLCELL_X8 FILLER_93_209 ();
 FILLCELL_X2 FILLER_93_217 ();
 FILLCELL_X2 FILLER_93_226 ();
 FILLCELL_X4 FILLER_93_235 ();
 FILLCELL_X16 FILLER_93_246 ();
 FILLCELL_X4 FILLER_93_293 ();
 FILLCELL_X2 FILLER_93_297 ();
 FILLCELL_X1 FILLER_93_299 ();
 FILLCELL_X1 FILLER_93_307 ();
 FILLCELL_X4 FILLER_93_315 ();
 FILLCELL_X2 FILLER_93_319 ();
 FILLCELL_X16 FILLER_93_328 ();
 FILLCELL_X2 FILLER_93_344 ();
 FILLCELL_X16 FILLER_93_381 ();
 FILLCELL_X4 FILLER_93_397 ();
 FILLCELL_X1 FILLER_93_401 ();
 FILLCELL_X1 FILLER_93_419 ();
 FILLCELL_X8 FILLER_93_429 ();
 FILLCELL_X2 FILLER_93_437 ();
 FILLCELL_X16 FILLER_93_444 ();
 FILLCELL_X8 FILLER_93_460 ();
 FILLCELL_X4 FILLER_93_468 ();
 FILLCELL_X2 FILLER_93_486 ();
 FILLCELL_X1 FILLER_93_488 ();
 FILLCELL_X4 FILLER_93_496 ();
 FILLCELL_X2 FILLER_93_509 ();
 FILLCELL_X1 FILLER_93_525 ();
 FILLCELL_X4 FILLER_93_543 ();
 FILLCELL_X1 FILLER_93_547 ();
 FILLCELL_X16 FILLER_93_551 ();
 FILLCELL_X4 FILLER_93_567 ();
 FILLCELL_X4 FILLER_93_578 ();
 FILLCELL_X2 FILLER_93_599 ();
 FILLCELL_X1 FILLER_93_601 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X2 FILLER_93_673 ();
 FILLCELL_X2 FILLER_93_680 ();
 FILLCELL_X2 FILLER_93_689 ();
 FILLCELL_X1 FILLER_93_691 ();
 FILLCELL_X16 FILLER_93_706 ();
 FILLCELL_X4 FILLER_93_722 ();
 FILLCELL_X2 FILLER_93_726 ();
 FILLCELL_X1 FILLER_93_728 ();
 FILLCELL_X2 FILLER_93_761 ();
 FILLCELL_X16 FILLER_93_766 ();
 FILLCELL_X2 FILLER_93_782 ();
 FILLCELL_X1 FILLER_93_784 ();
 FILLCELL_X4 FILLER_93_806 ();
 FILLCELL_X1 FILLER_93_810 ();
 FILLCELL_X8 FILLER_93_828 ();
 FILLCELL_X2 FILLER_93_836 ();
 FILLCELL_X1 FILLER_93_849 ();
 FILLCELL_X2 FILLER_93_862 ();
 FILLCELL_X1 FILLER_93_898 ();
 FILLCELL_X2 FILLER_93_902 ();
 FILLCELL_X2 FILLER_93_946 ();
 FILLCELL_X16 FILLER_93_957 ();
 FILLCELL_X1 FILLER_93_973 ();
 FILLCELL_X1 FILLER_93_984 ();
 FILLCELL_X16 FILLER_93_990 ();
 FILLCELL_X2 FILLER_93_1006 ();
 FILLCELL_X4 FILLER_93_1012 ();
 FILLCELL_X8 FILLER_93_1050 ();
 FILLCELL_X1 FILLER_93_1058 ();
 FILLCELL_X4 FILLER_93_1062 ();
 FILLCELL_X1 FILLER_93_1066 ();
 FILLCELL_X32 FILLER_93_1094 ();
 FILLCELL_X16 FILLER_93_1126 ();
 FILLCELL_X4 FILLER_93_1142 ();
 FILLCELL_X1 FILLER_93_1146 ();
 FILLCELL_X8 FILLER_93_1181 ();
 FILLCELL_X2 FILLER_93_1189 ();
 FILLCELL_X1 FILLER_93_1198 ();
 FILLCELL_X4 FILLER_93_1204 ();
 FILLCELL_X2 FILLER_93_1208 ();
 FILLCELL_X8 FILLER_93_1220 ();
 FILLCELL_X4 FILLER_93_1228 ();
 FILLCELL_X2 FILLER_93_1232 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X16 FILLER_94_33 ();
 FILLCELL_X1 FILLER_94_49 ();
 FILLCELL_X4 FILLER_94_57 ();
 FILLCELL_X2 FILLER_94_61 ();
 FILLCELL_X1 FILLER_94_80 ();
 FILLCELL_X8 FILLER_94_95 ();
 FILLCELL_X1 FILLER_94_103 ();
 FILLCELL_X8 FILLER_94_111 ();
 FILLCELL_X4 FILLER_94_119 ();
 FILLCELL_X1 FILLER_94_123 ();
 FILLCELL_X8 FILLER_94_127 ();
 FILLCELL_X4 FILLER_94_142 ();
 FILLCELL_X2 FILLER_94_146 ();
 FILLCELL_X1 FILLER_94_148 ();
 FILLCELL_X16 FILLER_94_156 ();
 FILLCELL_X4 FILLER_94_172 ();
 FILLCELL_X2 FILLER_94_176 ();
 FILLCELL_X1 FILLER_94_178 ();
 FILLCELL_X4 FILLER_94_186 ();
 FILLCELL_X1 FILLER_94_190 ();
 FILLCELL_X4 FILLER_94_199 ();
 FILLCELL_X2 FILLER_94_203 ();
 FILLCELL_X1 FILLER_94_205 ();
 FILLCELL_X8 FILLER_94_209 ();
 FILLCELL_X4 FILLER_94_224 ();
 FILLCELL_X2 FILLER_94_228 ();
 FILLCELL_X1 FILLER_94_230 ();
 FILLCELL_X4 FILLER_94_245 ();
 FILLCELL_X2 FILLER_94_249 ();
 FILLCELL_X2 FILLER_94_265 ();
 FILLCELL_X1 FILLER_94_267 ();
 FILLCELL_X4 FILLER_94_343 ();
 FILLCELL_X1 FILLER_94_347 ();
 FILLCELL_X2 FILLER_94_362 ();
 FILLCELL_X1 FILLER_94_364 ();
 FILLCELL_X16 FILLER_94_372 ();
 FILLCELL_X8 FILLER_94_388 ();
 FILLCELL_X4 FILLER_94_396 ();
 FILLCELL_X2 FILLER_94_400 ();
 FILLCELL_X1 FILLER_94_402 ();
 FILLCELL_X2 FILLER_94_430 ();
 FILLCELL_X4 FILLER_94_435 ();
 FILLCELL_X4 FILLER_94_465 ();
 FILLCELL_X4 FILLER_94_476 ();
 FILLCELL_X2 FILLER_94_480 ();
 FILLCELL_X1 FILLER_94_506 ();
 FILLCELL_X16 FILLER_94_514 ();
 FILLCELL_X2 FILLER_94_537 ();
 FILLCELL_X4 FILLER_94_546 ();
 FILLCELL_X4 FILLER_94_557 ();
 FILLCELL_X2 FILLER_94_568 ();
 FILLCELL_X1 FILLER_94_570 ();
 FILLCELL_X4 FILLER_94_588 ();
 FILLCELL_X1 FILLER_94_592 ();
 FILLCELL_X8 FILLER_94_617 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X4 FILLER_94_664 ();
 FILLCELL_X2 FILLER_94_668 ();
 FILLCELL_X2 FILLER_94_684 ();
 FILLCELL_X8 FILLER_94_703 ();
 FILLCELL_X4 FILLER_94_711 ();
 FILLCELL_X1 FILLER_94_743 ();
 FILLCELL_X4 FILLER_94_764 ();
 FILLCELL_X1 FILLER_94_768 ();
 FILLCELL_X2 FILLER_94_779 ();
 FILLCELL_X1 FILLER_94_781 ();
 FILLCELL_X4 FILLER_94_789 ();
 FILLCELL_X2 FILLER_94_793 ();
 FILLCELL_X16 FILLER_94_800 ();
 FILLCELL_X8 FILLER_94_816 ();
 FILLCELL_X4 FILLER_94_824 ();
 FILLCELL_X2 FILLER_94_828 ();
 FILLCELL_X2 FILLER_94_846 ();
 FILLCELL_X1 FILLER_94_848 ();
 FILLCELL_X4 FILLER_94_862 ();
 FILLCELL_X1 FILLER_94_866 ();
 FILLCELL_X1 FILLER_94_872 ();
 FILLCELL_X1 FILLER_94_909 ();
 FILLCELL_X4 FILLER_94_931 ();
 FILLCELL_X1 FILLER_94_935 ();
 FILLCELL_X1 FILLER_94_948 ();
 FILLCELL_X8 FILLER_94_953 ();
 FILLCELL_X1 FILLER_94_961 ();
 FILLCELL_X32 FILLER_94_969 ();
 FILLCELL_X16 FILLER_94_1001 ();
 FILLCELL_X2 FILLER_94_1075 ();
 FILLCELL_X16 FILLER_94_1087 ();
 FILLCELL_X1 FILLER_94_1120 ();
 FILLCELL_X8 FILLER_94_1150 ();
 FILLCELL_X4 FILLER_94_1158 ();
 FILLCELL_X2 FILLER_94_1179 ();
 FILLCELL_X1 FILLER_94_1181 ();
 FILLCELL_X1 FILLER_94_1199 ();
 FILLCELL_X2 FILLER_94_1217 ();
 FILLCELL_X2 FILLER_94_1226 ();
 FILLCELL_X2 FILLER_94_1235 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X8 FILLER_95_33 ();
 FILLCELL_X1 FILLER_95_41 ();
 FILLCELL_X1 FILLER_95_70 ();
 FILLCELL_X4 FILLER_95_78 ();
 FILLCELL_X2 FILLER_95_82 ();
 FILLCELL_X4 FILLER_95_125 ();
 FILLCELL_X2 FILLER_95_129 ();
 FILLCELL_X1 FILLER_95_131 ();
 FILLCELL_X1 FILLER_95_139 ();
 FILLCELL_X4 FILLER_95_147 ();
 FILLCELL_X1 FILLER_95_151 ();
 FILLCELL_X4 FILLER_95_159 ();
 FILLCELL_X1 FILLER_95_187 ();
 FILLCELL_X4 FILLER_95_195 ();
 FILLCELL_X16 FILLER_95_206 ();
 FILLCELL_X4 FILLER_95_256 ();
 FILLCELL_X2 FILLER_95_260 ();
 FILLCELL_X4 FILLER_95_290 ();
 FILLCELL_X1 FILLER_95_294 ();
 FILLCELL_X4 FILLER_95_300 ();
 FILLCELL_X2 FILLER_95_304 ();
 FILLCELL_X1 FILLER_95_306 ();
 FILLCELL_X4 FILLER_95_321 ();
 FILLCELL_X2 FILLER_95_325 ();
 FILLCELL_X1 FILLER_95_344 ();
 FILLCELL_X2 FILLER_95_352 ();
 FILLCELL_X16 FILLER_95_378 ();
 FILLCELL_X8 FILLER_95_394 ();
 FILLCELL_X4 FILLER_95_402 ();
 FILLCELL_X4 FILLER_95_413 ();
 FILLCELL_X1 FILLER_95_417 ();
 FILLCELL_X4 FILLER_95_425 ();
 FILLCELL_X4 FILLER_95_434 ();
 FILLCELL_X2 FILLER_95_438 ();
 FILLCELL_X16 FILLER_95_471 ();
 FILLCELL_X8 FILLER_95_494 ();
 FILLCELL_X2 FILLER_95_519 ();
 FILLCELL_X4 FILLER_95_531 ();
 FILLCELL_X2 FILLER_95_535 ();
 FILLCELL_X8 FILLER_95_541 ();
 FILLCELL_X4 FILLER_95_549 ();
 FILLCELL_X1 FILLER_95_553 ();
 FILLCELL_X16 FILLER_95_571 ();
 FILLCELL_X1 FILLER_95_594 ();
 FILLCELL_X32 FILLER_95_612 ();
 FILLCELL_X32 FILLER_95_644 ();
 FILLCELL_X2 FILLER_95_676 ();
 FILLCELL_X16 FILLER_95_685 ();
 FILLCELL_X4 FILLER_95_701 ();
 FILLCELL_X16 FILLER_95_736 ();
 FILLCELL_X8 FILLER_95_752 ();
 FILLCELL_X4 FILLER_95_760 ();
 FILLCELL_X2 FILLER_95_785 ();
 FILLCELL_X32 FILLER_95_804 ();
 FILLCELL_X16 FILLER_95_841 ();
 FILLCELL_X1 FILLER_95_857 ();
 FILLCELL_X2 FILLER_95_874 ();
 FILLCELL_X1 FILLER_95_876 ();
 FILLCELL_X2 FILLER_95_888 ();
 FILLCELL_X16 FILLER_95_926 ();
 FILLCELL_X4 FILLER_95_945 ();
 FILLCELL_X2 FILLER_95_949 ();
 FILLCELL_X2 FILLER_95_990 ();
 FILLCELL_X16 FILLER_95_1003 ();
 FILLCELL_X4 FILLER_95_1019 ();
 FILLCELL_X2 FILLER_95_1023 ();
 FILLCELL_X1 FILLER_95_1025 ();
 FILLCELL_X1 FILLER_95_1040 ();
 FILLCELL_X2 FILLER_95_1048 ();
 FILLCELL_X2 FILLER_95_1057 ();
 FILLCELL_X2 FILLER_95_1076 ();
 FILLCELL_X1 FILLER_95_1078 ();
 FILLCELL_X4 FILLER_95_1096 ();
 FILLCELL_X2 FILLER_95_1117 ();
 FILLCELL_X1 FILLER_95_1119 ();
 FILLCELL_X2 FILLER_95_1189 ();
 FILLCELL_X2 FILLER_95_1198 ();
 FILLCELL_X1 FILLER_95_1207 ();
 FILLCELL_X1 FILLER_95_1239 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X16 FILLER_96_65 ();
 FILLCELL_X8 FILLER_96_81 ();
 FILLCELL_X4 FILLER_96_89 ();
 FILLCELL_X1 FILLER_96_93 ();
 FILLCELL_X4 FILLER_96_101 ();
 FILLCELL_X2 FILLER_96_129 ();
 FILLCELL_X2 FILLER_96_167 ();
 FILLCELL_X1 FILLER_96_169 ();
 FILLCELL_X4 FILLER_96_177 ();
 FILLCELL_X1 FILLER_96_181 ();
 FILLCELL_X2 FILLER_96_199 ();
 FILLCELL_X4 FILLER_96_218 ();
 FILLCELL_X1 FILLER_96_222 ();
 FILLCELL_X4 FILLER_96_247 ();
 FILLCELL_X1 FILLER_96_251 ();
 FILLCELL_X16 FILLER_96_269 ();
 FILLCELL_X4 FILLER_96_285 ();
 FILLCELL_X2 FILLER_96_289 ();
 FILLCELL_X1 FILLER_96_291 ();
 FILLCELL_X4 FILLER_96_323 ();
 FILLCELL_X1 FILLER_96_327 ();
 FILLCELL_X4 FILLER_96_345 ();
 FILLCELL_X1 FILLER_96_349 ();
 FILLCELL_X8 FILLER_96_378 ();
 FILLCELL_X2 FILLER_96_386 ();
 FILLCELL_X1 FILLER_96_388 ();
 FILLCELL_X8 FILLER_96_413 ();
 FILLCELL_X2 FILLER_96_421 ();
 FILLCELL_X1 FILLER_96_423 ();
 FILLCELL_X16 FILLER_96_432 ();
 FILLCELL_X4 FILLER_96_448 ();
 FILLCELL_X1 FILLER_96_452 ();
 FILLCELL_X8 FILLER_96_491 ();
 FILLCELL_X4 FILLER_96_499 ();
 FILLCELL_X8 FILLER_96_517 ();
 FILLCELL_X4 FILLER_96_525 ();
 FILLCELL_X1 FILLER_96_529 ();
 FILLCELL_X16 FILLER_96_551 ();
 FILLCELL_X2 FILLER_96_567 ();
 FILLCELL_X1 FILLER_96_569 ();
 FILLCELL_X8 FILLER_96_584 ();
 FILLCELL_X16 FILLER_96_599 ();
 FILLCELL_X8 FILLER_96_615 ();
 FILLCELL_X1 FILLER_96_623 ();
 FILLCELL_X1 FILLER_96_632 ();
 FILLCELL_X8 FILLER_96_657 ();
 FILLCELL_X4 FILLER_96_665 ();
 FILLCELL_X2 FILLER_96_669 ();
 FILLCELL_X8 FILLER_96_688 ();
 FILLCELL_X4 FILLER_96_696 ();
 FILLCELL_X4 FILLER_96_748 ();
 FILLCELL_X2 FILLER_96_752 ();
 FILLCELL_X2 FILLER_96_778 ();
 FILLCELL_X1 FILLER_96_780 ();
 FILLCELL_X32 FILLER_96_805 ();
 FILLCELL_X4 FILLER_96_837 ();
 FILLCELL_X16 FILLER_96_851 ();
 FILLCELL_X4 FILLER_96_867 ();
 FILLCELL_X2 FILLER_96_871 ();
 FILLCELL_X1 FILLER_96_873 ();
 FILLCELL_X4 FILLER_96_899 ();
 FILLCELL_X4 FILLER_96_909 ();
 FILLCELL_X8 FILLER_96_916 ();
 FILLCELL_X2 FILLER_96_924 ();
 FILLCELL_X8 FILLER_96_947 ();
 FILLCELL_X4 FILLER_96_955 ();
 FILLCELL_X2 FILLER_96_959 ();
 FILLCELL_X8 FILLER_96_991 ();
 FILLCELL_X2 FILLER_96_999 ();
 FILLCELL_X1 FILLER_96_1001 ();
 FILLCELL_X8 FILLER_96_1008 ();
 FILLCELL_X4 FILLER_96_1016 ();
 FILLCELL_X2 FILLER_96_1020 ();
 FILLCELL_X1 FILLER_96_1022 ();
 FILLCELL_X16 FILLER_96_1026 ();
 FILLCELL_X8 FILLER_96_1042 ();
 FILLCELL_X2 FILLER_96_1050 ();
 FILLCELL_X8 FILLER_96_1057 ();
 FILLCELL_X1 FILLER_96_1065 ();
 FILLCELL_X4 FILLER_96_1083 ();
 FILLCELL_X2 FILLER_96_1087 ();
 FILLCELL_X1 FILLER_96_1089 ();
 FILLCELL_X4 FILLER_96_1103 ();
 FILLCELL_X1 FILLER_96_1107 ();
 FILLCELL_X32 FILLER_96_1143 ();
 FILLCELL_X4 FILLER_96_1175 ();
 FILLCELL_X2 FILLER_96_1179 ();
 FILLCELL_X1 FILLER_96_1218 ();
 FILLCELL_X1 FILLER_96_1222 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X16 FILLER_97_33 ();
 FILLCELL_X2 FILLER_97_49 ();
 FILLCELL_X1 FILLER_97_51 ();
 FILLCELL_X8 FILLER_97_86 ();
 FILLCELL_X4 FILLER_97_94 ();
 FILLCELL_X16 FILLER_97_112 ();
 FILLCELL_X1 FILLER_97_142 ();
 FILLCELL_X1 FILLER_97_160 ();
 FILLCELL_X2 FILLER_97_168 ();
 FILLCELL_X1 FILLER_97_174 ();
 FILLCELL_X8 FILLER_97_192 ();
 FILLCELL_X1 FILLER_97_200 ();
 FILLCELL_X32 FILLER_97_218 ();
 FILLCELL_X4 FILLER_97_250 ();
 FILLCELL_X2 FILLER_97_254 ();
 FILLCELL_X32 FILLER_97_263 ();
 FILLCELL_X1 FILLER_97_295 ();
 FILLCELL_X4 FILLER_97_303 ();
 FILLCELL_X2 FILLER_97_307 ();
 FILLCELL_X1 FILLER_97_309 ();
 FILLCELL_X4 FILLER_97_321 ();
 FILLCELL_X1 FILLER_97_357 ();
 FILLCELL_X2 FILLER_97_371 ();
 FILLCELL_X1 FILLER_97_373 ();
 FILLCELL_X8 FILLER_97_378 ();
 FILLCELL_X4 FILLER_97_417 ();
 FILLCELL_X1 FILLER_97_421 ();
 FILLCELL_X16 FILLER_97_429 ();
 FILLCELL_X4 FILLER_97_445 ();
 FILLCELL_X2 FILLER_97_456 ();
 FILLCELL_X2 FILLER_97_482 ();
 FILLCELL_X1 FILLER_97_484 ();
 FILLCELL_X2 FILLER_97_502 ();
 FILLCELL_X1 FILLER_97_504 ();
 FILLCELL_X4 FILLER_97_522 ();
 FILLCELL_X1 FILLER_97_526 ();
 FILLCELL_X4 FILLER_97_551 ();
 FILLCELL_X2 FILLER_97_555 ();
 FILLCELL_X1 FILLER_97_557 ();
 FILLCELL_X1 FILLER_97_575 ();
 FILLCELL_X1 FILLER_97_606 ();
 FILLCELL_X8 FILLER_97_662 ();
 FILLCELL_X4 FILLER_97_670 ();
 FILLCELL_X2 FILLER_97_674 ();
 FILLCELL_X2 FILLER_97_683 ();
 FILLCELL_X1 FILLER_97_685 ();
 FILLCELL_X16 FILLER_97_710 ();
 FILLCELL_X4 FILLER_97_726 ();
 FILLCELL_X8 FILLER_97_743 ();
 FILLCELL_X4 FILLER_97_759 ();
 FILLCELL_X1 FILLER_97_763 ();
 FILLCELL_X2 FILLER_97_781 ();
 FILLCELL_X1 FILLER_97_787 ();
 FILLCELL_X16 FILLER_97_801 ();
 FILLCELL_X1 FILLER_97_817 ();
 FILLCELL_X1 FILLER_97_840 ();
 FILLCELL_X1 FILLER_97_845 ();
 FILLCELL_X8 FILLER_97_878 ();
 FILLCELL_X4 FILLER_97_886 ();
 FILLCELL_X1 FILLER_97_890 ();
 FILLCELL_X16 FILLER_97_911 ();
 FILLCELL_X2 FILLER_97_927 ();
 FILLCELL_X4 FILLER_97_950 ();
 FILLCELL_X2 FILLER_97_954 ();
 FILLCELL_X1 FILLER_97_956 ();
 FILLCELL_X1 FILLER_97_976 ();
 FILLCELL_X1 FILLER_97_982 ();
 FILLCELL_X1 FILLER_97_985 ();
 FILLCELL_X1 FILLER_97_989 ();
 FILLCELL_X2 FILLER_97_1001 ();
 FILLCELL_X1 FILLER_97_1003 ();
 FILLCELL_X16 FILLER_97_1009 ();
 FILLCELL_X2 FILLER_97_1025 ();
 FILLCELL_X16 FILLER_97_1030 ();
 FILLCELL_X8 FILLER_97_1046 ();
 FILLCELL_X2 FILLER_97_1054 ();
 FILLCELL_X16 FILLER_97_1080 ();
 FILLCELL_X32 FILLER_97_1101 ();
 FILLCELL_X2 FILLER_97_1147 ();
 FILLCELL_X2 FILLER_97_1174 ();
 FILLCELL_X1 FILLER_97_1176 ();
 FILLCELL_X1 FILLER_97_1191 ();
 FILLCELL_X4 FILLER_97_1202 ();
 FILLCELL_X1 FILLER_97_1209 ();
 FILLCELL_X2 FILLER_97_1238 ();
 FILLCELL_X16 FILLER_98_1 ();
 FILLCELL_X4 FILLER_98_17 ();
 FILLCELL_X2 FILLER_98_21 ();
 FILLCELL_X4 FILLER_98_26 ();
 FILLCELL_X2 FILLER_98_30 ();
 FILLCELL_X1 FILLER_98_32 ();
 FILLCELL_X16 FILLER_98_40 ();
 FILLCELL_X1 FILLER_98_56 ();
 FILLCELL_X8 FILLER_98_64 ();
 FILLCELL_X16 FILLER_98_86 ();
 FILLCELL_X8 FILLER_98_102 ();
 FILLCELL_X4 FILLER_98_110 ();
 FILLCELL_X8 FILLER_98_121 ();
 FILLCELL_X4 FILLER_98_129 ();
 FILLCELL_X2 FILLER_98_150 ();
 FILLCELL_X16 FILLER_98_159 ();
 FILLCELL_X2 FILLER_98_182 ();
 FILLCELL_X8 FILLER_98_191 ();
 FILLCELL_X1 FILLER_98_199 ();
 FILLCELL_X16 FILLER_98_221 ();
 FILLCELL_X4 FILLER_98_237 ();
 FILLCELL_X2 FILLER_98_241 ();
 FILLCELL_X1 FILLER_98_243 ();
 FILLCELL_X8 FILLER_98_276 ();
 FILLCELL_X4 FILLER_98_284 ();
 FILLCELL_X2 FILLER_98_305 ();
 FILLCELL_X1 FILLER_98_335 ();
 FILLCELL_X1 FILLER_98_342 ();
 FILLCELL_X2 FILLER_98_356 ();
 FILLCELL_X2 FILLER_98_384 ();
 FILLCELL_X1 FILLER_98_386 ();
 FILLCELL_X8 FILLER_98_394 ();
 FILLCELL_X4 FILLER_98_402 ();
 FILLCELL_X2 FILLER_98_406 ();
 FILLCELL_X1 FILLER_98_408 ();
 FILLCELL_X8 FILLER_98_433 ();
 FILLCELL_X4 FILLER_98_441 ();
 FILLCELL_X2 FILLER_98_469 ();
 FILLCELL_X8 FILLER_98_474 ();
 FILLCELL_X1 FILLER_98_487 ();
 FILLCELL_X1 FILLER_98_502 ();
 FILLCELL_X2 FILLER_98_523 ();
 FILLCELL_X1 FILLER_98_525 ();
 FILLCELL_X8 FILLER_98_550 ();
 FILLCELL_X4 FILLER_98_558 ();
 FILLCELL_X1 FILLER_98_562 ();
 FILLCELL_X16 FILLER_98_580 ();
 FILLCELL_X4 FILLER_98_596 ();
 FILLCELL_X2 FILLER_98_600 ();
 FILLCELL_X1 FILLER_98_602 ();
 FILLCELL_X8 FILLER_98_623 ();
 FILLCELL_X1 FILLER_98_632 ();
 FILLCELL_X8 FILLER_98_662 ();
 FILLCELL_X4 FILLER_98_670 ();
 FILLCELL_X1 FILLER_98_706 ();
 FILLCELL_X2 FILLER_98_714 ();
 FILLCELL_X1 FILLER_98_716 ();
 FILLCELL_X1 FILLER_98_722 ();
 FILLCELL_X8 FILLER_98_734 ();
 FILLCELL_X1 FILLER_98_742 ();
 FILLCELL_X32 FILLER_98_773 ();
 FILLCELL_X4 FILLER_98_805 ();
 FILLCELL_X2 FILLER_98_809 ();
 FILLCELL_X1 FILLER_98_811 ();
 FILLCELL_X4 FILLER_98_843 ();
 FILLCELL_X2 FILLER_98_847 ();
 FILLCELL_X1 FILLER_98_849 ();
 FILLCELL_X1 FILLER_98_868 ();
 FILLCELL_X4 FILLER_98_886 ();
 FILLCELL_X1 FILLER_98_911 ();
 FILLCELL_X2 FILLER_98_919 ();
 FILLCELL_X2 FILLER_98_930 ();
 FILLCELL_X8 FILLER_98_958 ();
 FILLCELL_X2 FILLER_98_982 ();
 FILLCELL_X1 FILLER_98_997 ();
 FILLCELL_X4 FILLER_98_1013 ();
 FILLCELL_X2 FILLER_98_1017 ();
 FILLCELL_X1 FILLER_98_1019 ();
 FILLCELL_X16 FILLER_98_1030 ();
 FILLCELL_X8 FILLER_98_1046 ();
 FILLCELL_X4 FILLER_98_1054 ();
 FILLCELL_X2 FILLER_98_1058 ();
 FILLCELL_X1 FILLER_98_1060 ();
 FILLCELL_X16 FILLER_98_1078 ();
 FILLCELL_X4 FILLER_98_1094 ();
 FILLCELL_X2 FILLER_98_1098 ();
 FILLCELL_X16 FILLER_98_1107 ();
 FILLCELL_X1 FILLER_98_1123 ();
 FILLCELL_X8 FILLER_98_1131 ();
 FILLCELL_X4 FILLER_98_1139 ();
 FILLCELL_X1 FILLER_98_1143 ();
 FILLCELL_X8 FILLER_98_1176 ();
 FILLCELL_X1 FILLER_98_1184 ();
 FILLCELL_X4 FILLER_98_1192 ();
 FILLCELL_X2 FILLER_98_1238 ();
 FILLCELL_X16 FILLER_99_1 ();
 FILLCELL_X8 FILLER_99_17 ();
 FILLCELL_X4 FILLER_99_25 ();
 FILLCELL_X2 FILLER_99_46 ();
 FILLCELL_X1 FILLER_99_48 ();
 FILLCELL_X1 FILLER_99_73 ();
 FILLCELL_X16 FILLER_99_81 ();
 FILLCELL_X1 FILLER_99_114 ();
 FILLCELL_X16 FILLER_99_122 ();
 FILLCELL_X4 FILLER_99_138 ();
 FILLCELL_X1 FILLER_99_142 ();
 FILLCELL_X4 FILLER_99_148 ();
 FILLCELL_X2 FILLER_99_152 ();
 FILLCELL_X4 FILLER_99_161 ();
 FILLCELL_X1 FILLER_99_165 ();
 FILLCELL_X32 FILLER_99_173 ();
 FILLCELL_X1 FILLER_99_205 ();
 FILLCELL_X8 FILLER_99_213 ();
 FILLCELL_X4 FILLER_99_221 ();
 FILLCELL_X2 FILLER_99_225 ();
 FILLCELL_X4 FILLER_99_244 ();
 FILLCELL_X8 FILLER_99_276 ();
 FILLCELL_X4 FILLER_99_284 ();
 FILLCELL_X1 FILLER_99_295 ();
 FILLCELL_X1 FILLER_99_310 ();
 FILLCELL_X1 FILLER_99_328 ();
 FILLCELL_X1 FILLER_99_336 ();
 FILLCELL_X1 FILLER_99_349 ();
 FILLCELL_X2 FILLER_99_374 ();
 FILLCELL_X16 FILLER_99_426 ();
 FILLCELL_X8 FILLER_99_442 ();
 FILLCELL_X16 FILLER_99_464 ();
 FILLCELL_X8 FILLER_99_480 ();
 FILLCELL_X4 FILLER_99_492 ();
 FILLCELL_X2 FILLER_99_496 ();
 FILLCELL_X1 FILLER_99_498 ();
 FILLCELL_X1 FILLER_99_530 ();
 FILLCELL_X1 FILLER_99_538 ();
 FILLCELL_X16 FILLER_99_546 ();
 FILLCELL_X8 FILLER_99_562 ();
 FILLCELL_X4 FILLER_99_570 ();
 FILLCELL_X2 FILLER_99_574 ();
 FILLCELL_X1 FILLER_99_576 ();
 FILLCELL_X2 FILLER_99_584 ();
 FILLCELL_X1 FILLER_99_586 ();
 FILLCELL_X32 FILLER_99_604 ();
 FILLCELL_X2 FILLER_99_636 ();
 FILLCELL_X4 FILLER_99_645 ();
 FILLCELL_X1 FILLER_99_649 ();
 FILLCELL_X4 FILLER_99_653 ();
 FILLCELL_X2 FILLER_99_657 ();
 FILLCELL_X1 FILLER_99_659 ();
 FILLCELL_X2 FILLER_99_672 ();
 FILLCELL_X4 FILLER_99_681 ();
 FILLCELL_X4 FILLER_99_692 ();
 FILLCELL_X2 FILLER_99_696 ();
 FILLCELL_X8 FILLER_99_768 ();
 FILLCELL_X4 FILLER_99_776 ();
 FILLCELL_X16 FILLER_99_790 ();
 FILLCELL_X8 FILLER_99_806 ();
 FILLCELL_X4 FILLER_99_814 ();
 FILLCELL_X1 FILLER_99_818 ();
 FILLCELL_X8 FILLER_99_825 ();
 FILLCELL_X1 FILLER_99_833 ();
 FILLCELL_X1 FILLER_99_865 ();
 FILLCELL_X1 FILLER_99_884 ();
 FILLCELL_X1 FILLER_99_896 ();
 FILLCELL_X4 FILLER_99_918 ();
 FILLCELL_X2 FILLER_99_947 ();
 FILLCELL_X16 FILLER_99_960 ();
 FILLCELL_X4 FILLER_99_976 ();
 FILLCELL_X1 FILLER_99_980 ();
 FILLCELL_X4 FILLER_99_984 ();
 FILLCELL_X16 FILLER_99_991 ();
 FILLCELL_X1 FILLER_99_1017 ();
 FILLCELL_X16 FILLER_99_1041 ();
 FILLCELL_X8 FILLER_99_1057 ();
 FILLCELL_X1 FILLER_99_1065 ();
 FILLCELL_X16 FILLER_99_1073 ();
 FILLCELL_X2 FILLER_99_1089 ();
 FILLCELL_X1 FILLER_99_1091 ();
 FILLCELL_X1 FILLER_99_1122 ();
 FILLCELL_X4 FILLER_99_1137 ();
 FILLCELL_X2 FILLER_99_1141 ();
 FILLCELL_X1 FILLER_99_1165 ();
 FILLCELL_X4 FILLER_99_1183 ();
 FILLCELL_X4 FILLER_99_1194 ();
 FILLCELL_X1 FILLER_99_1198 ();
 FILLCELL_X8 FILLER_100_1 ();
 FILLCELL_X4 FILLER_100_9 ();
 FILLCELL_X2 FILLER_100_13 ();
 FILLCELL_X1 FILLER_100_15 ();
 FILLCELL_X4 FILLER_100_40 ();
 FILLCELL_X2 FILLER_100_44 ();
 FILLCELL_X1 FILLER_100_53 ();
 FILLCELL_X2 FILLER_100_61 ();
 FILLCELL_X1 FILLER_100_63 ();
 FILLCELL_X4 FILLER_100_71 ();
 FILLCELL_X1 FILLER_100_75 ();
 FILLCELL_X8 FILLER_100_83 ();
 FILLCELL_X4 FILLER_100_91 ();
 FILLCELL_X8 FILLER_100_126 ();
 FILLCELL_X16 FILLER_100_158 ();
 FILLCELL_X4 FILLER_100_174 ();
 FILLCELL_X4 FILLER_100_192 ();
 FILLCELL_X1 FILLER_100_196 ();
 FILLCELL_X4 FILLER_100_256 ();
 FILLCELL_X2 FILLER_100_260 ();
 FILLCELL_X32 FILLER_100_269 ();
 FILLCELL_X2 FILLER_100_301 ();
 FILLCELL_X1 FILLER_100_303 ();
 FILLCELL_X8 FILLER_100_321 ();
 FILLCELL_X4 FILLER_100_329 ();
 FILLCELL_X2 FILLER_100_333 ();
 FILLCELL_X1 FILLER_100_335 ();
 FILLCELL_X8 FILLER_100_341 ();
 FILLCELL_X1 FILLER_100_349 ();
 FILLCELL_X2 FILLER_100_370 ();
 FILLCELL_X16 FILLER_100_386 ();
 FILLCELL_X2 FILLER_100_402 ();
 FILLCELL_X4 FILLER_100_416 ();
 FILLCELL_X16 FILLER_100_427 ();
 FILLCELL_X2 FILLER_100_443 ();
 FILLCELL_X16 FILLER_100_462 ();
 FILLCELL_X4 FILLER_100_478 ();
 FILLCELL_X2 FILLER_100_482 ();
 FILLCELL_X4 FILLER_100_515 ();
 FILLCELL_X2 FILLER_100_519 ();
 FILLCELL_X4 FILLER_100_526 ();
 FILLCELL_X2 FILLER_100_530 ();
 FILLCELL_X1 FILLER_100_532 ();
 FILLCELL_X8 FILLER_100_550 ();
 FILLCELL_X4 FILLER_100_558 ();
 FILLCELL_X2 FILLER_100_582 ();
 FILLCELL_X4 FILLER_100_604 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X4 FILLER_100_645 ();
 FILLCELL_X4 FILLER_100_666 ();
 FILLCELL_X4 FILLER_100_712 ();
 FILLCELL_X2 FILLER_100_716 ();
 FILLCELL_X2 FILLER_100_725 ();
 FILLCELL_X8 FILLER_100_734 ();
 FILLCELL_X2 FILLER_100_742 ();
 FILLCELL_X1 FILLER_100_758 ();
 FILLCELL_X1 FILLER_100_766 ();
 FILLCELL_X1 FILLER_100_777 ();
 FILLCELL_X16 FILLER_100_787 ();
 FILLCELL_X8 FILLER_100_803 ();
 FILLCELL_X4 FILLER_100_811 ();
 FILLCELL_X4 FILLER_100_845 ();
 FILLCELL_X1 FILLER_100_849 ();
 FILLCELL_X1 FILLER_100_883 ();
 FILLCELL_X1 FILLER_100_894 ();
 FILLCELL_X2 FILLER_100_900 ();
 FILLCELL_X4 FILLER_100_910 ();
 FILLCELL_X16 FILLER_100_926 ();
 FILLCELL_X16 FILLER_100_958 ();
 FILLCELL_X4 FILLER_100_974 ();
 FILLCELL_X2 FILLER_100_978 ();
 FILLCELL_X16 FILLER_100_987 ();
 FILLCELL_X8 FILLER_100_1003 ();
 FILLCELL_X4 FILLER_100_1011 ();
 FILLCELL_X1 FILLER_100_1015 ();
 FILLCELL_X16 FILLER_100_1041 ();
 FILLCELL_X2 FILLER_100_1057 ();
 FILLCELL_X8 FILLER_100_1076 ();
 FILLCELL_X4 FILLER_100_1084 ();
 FILLCELL_X2 FILLER_100_1163 ();
 FILLCELL_X8 FILLER_100_1172 ();
 FILLCELL_X4 FILLER_100_1180 ();
 FILLCELL_X2 FILLER_100_1184 ();
 FILLCELL_X1 FILLER_100_1186 ();
 FILLCELL_X2 FILLER_100_1194 ();
 FILLCELL_X2 FILLER_100_1221 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X8 FILLER_101_33 ();
 FILLCELL_X4 FILLER_101_41 ();
 FILLCELL_X1 FILLER_101_45 ();
 FILLCELL_X8 FILLER_101_63 ();
 FILLCELL_X4 FILLER_101_71 ();
 FILLCELL_X1 FILLER_101_75 ();
 FILLCELL_X4 FILLER_101_107 ();
 FILLCELL_X1 FILLER_101_111 ();
 FILLCELL_X8 FILLER_101_119 ();
 FILLCELL_X2 FILLER_101_127 ();
 FILLCELL_X4 FILLER_101_146 ();
 FILLCELL_X1 FILLER_101_150 ();
 FILLCELL_X1 FILLER_101_168 ();
 FILLCELL_X2 FILLER_101_176 ();
 FILLCELL_X2 FILLER_101_195 ();
 FILLCELL_X1 FILLER_101_197 ();
 FILLCELL_X2 FILLER_101_220 ();
 FILLCELL_X1 FILLER_101_222 ();
 FILLCELL_X8 FILLER_101_232 ();
 FILLCELL_X8 FILLER_101_254 ();
 FILLCELL_X2 FILLER_101_262 ();
 FILLCELL_X32 FILLER_101_274 ();
 FILLCELL_X32 FILLER_101_306 ();
 FILLCELL_X8 FILLER_101_338 ();
 FILLCELL_X1 FILLER_101_346 ();
 FILLCELL_X4 FILLER_101_366 ();
 FILLCELL_X2 FILLER_101_370 ();
 FILLCELL_X8 FILLER_101_375 ();
 FILLCELL_X4 FILLER_101_383 ();
 FILLCELL_X2 FILLER_101_387 ();
 FILLCELL_X4 FILLER_101_394 ();
 FILLCELL_X2 FILLER_101_398 ();
 FILLCELL_X16 FILLER_101_424 ();
 FILLCELL_X2 FILLER_101_440 ();
 FILLCELL_X4 FILLER_101_459 ();
 FILLCELL_X2 FILLER_101_480 ();
 FILLCELL_X16 FILLER_101_499 ();
 FILLCELL_X8 FILLER_101_515 ();
 FILLCELL_X4 FILLER_101_523 ();
 FILLCELL_X1 FILLER_101_527 ();
 FILLCELL_X1 FILLER_101_535 ();
 FILLCELL_X1 FILLER_101_543 ();
 FILLCELL_X8 FILLER_101_551 ();
 FILLCELL_X4 FILLER_101_559 ();
 FILLCELL_X2 FILLER_101_563 ();
 FILLCELL_X4 FILLER_101_568 ();
 FILLCELL_X1 FILLER_101_572 ();
 FILLCELL_X1 FILLER_101_579 ();
 FILLCELL_X16 FILLER_101_586 ();
 FILLCELL_X2 FILLER_101_602 ();
 FILLCELL_X1 FILLER_101_604 ();
 FILLCELL_X1 FILLER_101_612 ();
 FILLCELL_X2 FILLER_101_620 ();
 FILLCELL_X1 FILLER_101_629 ();
 FILLCELL_X2 FILLER_101_664 ();
 FILLCELL_X4 FILLER_101_707 ();
 FILLCELL_X1 FILLER_101_711 ();
 FILLCELL_X8 FILLER_101_753 ();
 FILLCELL_X4 FILLER_101_761 ();
 FILLCELL_X1 FILLER_101_765 ();
 FILLCELL_X1 FILLER_101_776 ();
 FILLCELL_X32 FILLER_101_787 ();
 FILLCELL_X16 FILLER_101_819 ();
 FILLCELL_X8 FILLER_101_835 ();
 FILLCELL_X4 FILLER_101_843 ();
 FILLCELL_X1 FILLER_101_847 ();
 FILLCELL_X2 FILLER_101_851 ();
 FILLCELL_X1 FILLER_101_853 ();
 FILLCELL_X1 FILLER_101_860 ();
 FILLCELL_X1 FILLER_101_868 ();
 FILLCELL_X1 FILLER_101_879 ();
 FILLCELL_X8 FILLER_101_890 ();
 FILLCELL_X2 FILLER_101_898 ();
 FILLCELL_X8 FILLER_101_927 ();
 FILLCELL_X4 FILLER_101_935 ();
 FILLCELL_X2 FILLER_101_939 ();
 FILLCELL_X1 FILLER_101_941 ();
 FILLCELL_X4 FILLER_101_949 ();
 FILLCELL_X16 FILLER_101_967 ();
 FILLCELL_X2 FILLER_101_983 ();
 FILLCELL_X4 FILLER_101_1017 ();
 FILLCELL_X16 FILLER_101_1030 ();
 FILLCELL_X8 FILLER_101_1046 ();
 FILLCELL_X2 FILLER_101_1054 ();
 FILLCELL_X1 FILLER_101_1056 ();
 FILLCELL_X1 FILLER_101_1081 ();
 FILLCELL_X4 FILLER_101_1091 ();
 FILLCELL_X2 FILLER_101_1138 ();
 FILLCELL_X1 FILLER_101_1147 ();
 FILLCELL_X2 FILLER_101_1155 ();
 FILLCELL_X1 FILLER_101_1157 ();
 FILLCELL_X4 FILLER_101_1182 ();
 FILLCELL_X2 FILLER_101_1186 ();
 FILLCELL_X1 FILLER_101_1188 ();
 FILLCELL_X1 FILLER_101_1229 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X8 FILLER_102_33 ();
 FILLCELL_X4 FILLER_102_41 ();
 FILLCELL_X2 FILLER_102_45 ();
 FILLCELL_X4 FILLER_102_64 ();
 FILLCELL_X1 FILLER_102_75 ();
 FILLCELL_X4 FILLER_102_83 ();
 FILLCELL_X4 FILLER_102_94 ();
 FILLCELL_X1 FILLER_102_98 ();
 FILLCELL_X4 FILLER_102_106 ();
 FILLCELL_X1 FILLER_102_110 ();
 FILLCELL_X4 FILLER_102_118 ();
 FILLCELL_X2 FILLER_102_122 ();
 FILLCELL_X1 FILLER_102_124 ();
 FILLCELL_X2 FILLER_102_139 ();
 FILLCELL_X1 FILLER_102_141 ();
 FILLCELL_X4 FILLER_102_149 ();
 FILLCELL_X2 FILLER_102_153 ();
 FILLCELL_X4 FILLER_102_162 ();
 FILLCELL_X2 FILLER_102_166 ();
 FILLCELL_X4 FILLER_102_175 ();
 FILLCELL_X2 FILLER_102_196 ();
 FILLCELL_X16 FILLER_102_217 ();
 FILLCELL_X2 FILLER_102_233 ();
 FILLCELL_X4 FILLER_102_259 ();
 FILLCELL_X2 FILLER_102_263 ();
 FILLCELL_X1 FILLER_102_265 ();
 FILLCELL_X16 FILLER_102_280 ();
 FILLCELL_X2 FILLER_102_296 ();
 FILLCELL_X1 FILLER_102_298 ();
 FILLCELL_X1 FILLER_102_306 ();
 FILLCELL_X1 FILLER_102_314 ();
 FILLCELL_X2 FILLER_102_343 ();
 FILLCELL_X8 FILLER_102_391 ();
 FILLCELL_X2 FILLER_102_399 ();
 FILLCELL_X8 FILLER_102_405 ();
 FILLCELL_X8 FILLER_102_430 ();
 FILLCELL_X2 FILLER_102_438 ();
 FILLCELL_X1 FILLER_102_440 ();
 FILLCELL_X4 FILLER_102_448 ();
 FILLCELL_X1 FILLER_102_452 ();
 FILLCELL_X4 FILLER_102_467 ();
 FILLCELL_X4 FILLER_102_475 ();
 FILLCELL_X2 FILLER_102_479 ();
 FILLCELL_X1 FILLER_102_481 ();
 FILLCELL_X8 FILLER_102_496 ();
 FILLCELL_X2 FILLER_102_504 ();
 FILLCELL_X4 FILLER_102_526 ();
 FILLCELL_X8 FILLER_102_547 ();
 FILLCELL_X4 FILLER_102_555 ();
 FILLCELL_X1 FILLER_102_559 ();
 FILLCELL_X16 FILLER_102_585 ();
 FILLCELL_X4 FILLER_102_601 ();
 FILLCELL_X2 FILLER_102_605 ();
 FILLCELL_X8 FILLER_102_632 ();
 FILLCELL_X2 FILLER_102_640 ();
 FILLCELL_X4 FILLER_102_656 ();
 FILLCELL_X4 FILLER_102_697 ();
 FILLCELL_X32 FILLER_102_714 ();
 FILLCELL_X16 FILLER_102_746 ();
 FILLCELL_X2 FILLER_102_762 ();
 FILLCELL_X32 FILLER_102_789 ();
 FILLCELL_X16 FILLER_102_821 ();
 FILLCELL_X8 FILLER_102_837 ();
 FILLCELL_X2 FILLER_102_845 ();
 FILLCELL_X1 FILLER_102_847 ();
 FILLCELL_X8 FILLER_102_859 ();
 FILLCELL_X4 FILLER_102_867 ();
 FILLCELL_X2 FILLER_102_871 ();
 FILLCELL_X1 FILLER_102_873 ();
 FILLCELL_X2 FILLER_102_877 ();
 FILLCELL_X4 FILLER_102_881 ();
 FILLCELL_X8 FILLER_102_888 ();
 FILLCELL_X2 FILLER_102_896 ();
 FILLCELL_X2 FILLER_102_904 ();
 FILLCELL_X1 FILLER_102_906 ();
 FILLCELL_X8 FILLER_102_934 ();
 FILLCELL_X4 FILLER_102_946 ();
 FILLCELL_X2 FILLER_102_950 ();
 FILLCELL_X4 FILLER_102_959 ();
 FILLCELL_X2 FILLER_102_963 ();
 FILLCELL_X2 FILLER_102_967 ();
 FILLCELL_X2 FILLER_102_971 ();
 FILLCELL_X2 FILLER_102_980 ();
 FILLCELL_X1 FILLER_102_989 ();
 FILLCELL_X1 FILLER_102_992 ();
 FILLCELL_X1 FILLER_102_999 ();
 FILLCELL_X1 FILLER_102_1010 ();
 FILLCELL_X8 FILLER_102_1015 ();
 FILLCELL_X4 FILLER_102_1023 ();
 FILLCELL_X1 FILLER_102_1027 ();
 FILLCELL_X16 FILLER_102_1037 ();
 FILLCELL_X8 FILLER_102_1053 ();
 FILLCELL_X1 FILLER_102_1061 ();
 FILLCELL_X4 FILLER_102_1083 ();
 FILLCELL_X32 FILLER_102_1092 ();
 FILLCELL_X2 FILLER_102_1124 ();
 FILLCELL_X1 FILLER_102_1126 ();
 FILLCELL_X32 FILLER_102_1132 ();
 FILLCELL_X32 FILLER_102_1164 ();
 FILLCELL_X8 FILLER_102_1196 ();
 FILLCELL_X1 FILLER_102_1204 ();
 FILLCELL_X1 FILLER_102_1208 ();
 FILLCELL_X4 FILLER_102_1212 ();
 FILLCELL_X2 FILLER_102_1222 ();
 FILLCELL_X1 FILLER_102_1231 ();
 FILLCELL_X2 FILLER_102_1238 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X4 FILLER_103_33 ();
 FILLCELL_X8 FILLER_103_41 ();
 FILLCELL_X2 FILLER_103_49 ();
 FILLCELL_X8 FILLER_103_58 ();
 FILLCELL_X2 FILLER_103_66 ();
 FILLCELL_X8 FILLER_103_85 ();
 FILLCELL_X4 FILLER_103_93 ();
 FILLCELL_X2 FILLER_103_97 ();
 FILLCELL_X8 FILLER_103_116 ();
 FILLCELL_X4 FILLER_103_141 ();
 FILLCELL_X4 FILLER_103_152 ();
 FILLCELL_X2 FILLER_103_156 ();
 FILLCELL_X1 FILLER_103_158 ();
 FILLCELL_X2 FILLER_103_176 ();
 FILLCELL_X1 FILLER_103_178 ();
 FILLCELL_X4 FILLER_103_186 ();
 FILLCELL_X2 FILLER_103_190 ();
 FILLCELL_X1 FILLER_103_192 ();
 FILLCELL_X1 FILLER_103_200 ();
 FILLCELL_X16 FILLER_103_213 ();
 FILLCELL_X4 FILLER_103_229 ();
 FILLCELL_X2 FILLER_103_233 ();
 FILLCELL_X1 FILLER_103_235 ();
 FILLCELL_X1 FILLER_103_277 ();
 FILLCELL_X8 FILLER_103_292 ();
 FILLCELL_X8 FILLER_103_341 ();
 FILLCELL_X2 FILLER_103_349 ();
 FILLCELL_X4 FILLER_103_369 ();
 FILLCELL_X2 FILLER_103_403 ();
 FILLCELL_X16 FILLER_103_422 ();
 FILLCELL_X8 FILLER_103_438 ();
 FILLCELL_X4 FILLER_103_446 ();
 FILLCELL_X2 FILLER_103_457 ();
 FILLCELL_X1 FILLER_103_459 ();
 FILLCELL_X16 FILLER_103_495 ();
 FILLCELL_X8 FILLER_103_511 ();
 FILLCELL_X2 FILLER_103_519 ();
 FILLCELL_X1 FILLER_103_521 ();
 FILLCELL_X16 FILLER_103_535 ();
 FILLCELL_X1 FILLER_103_551 ();
 FILLCELL_X1 FILLER_103_569 ();
 FILLCELL_X1 FILLER_103_574 ();
 FILLCELL_X32 FILLER_103_588 ();
 FILLCELL_X4 FILLER_103_620 ();
 FILLCELL_X2 FILLER_103_624 ();
 FILLCELL_X1 FILLER_103_626 ();
 FILLCELL_X8 FILLER_103_631 ();
 FILLCELL_X4 FILLER_103_639 ();
 FILLCELL_X1 FILLER_103_643 ();
 FILLCELL_X8 FILLER_103_700 ();
 FILLCELL_X1 FILLER_103_708 ();
 FILLCELL_X2 FILLER_103_733 ();
 FILLCELL_X1 FILLER_103_735 ();
 FILLCELL_X16 FILLER_103_753 ();
 FILLCELL_X1 FILLER_103_769 ();
 FILLCELL_X1 FILLER_103_774 ();
 FILLCELL_X8 FILLER_103_800 ();
 FILLCELL_X4 FILLER_103_808 ();
 FILLCELL_X2 FILLER_103_812 ();
 FILLCELL_X32 FILLER_103_824 ();
 FILLCELL_X16 FILLER_103_870 ();
 FILLCELL_X4 FILLER_103_886 ();
 FILLCELL_X2 FILLER_103_901 ();
 FILLCELL_X1 FILLER_103_912 ();
 FILLCELL_X2 FILLER_103_924 ();
 FILLCELL_X2 FILLER_103_939 ();
 FILLCELL_X2 FILLER_103_958 ();
 FILLCELL_X4 FILLER_103_980 ();
 FILLCELL_X16 FILLER_103_1003 ();
 FILLCELL_X8 FILLER_103_1019 ();
 FILLCELL_X2 FILLER_103_1027 ();
 FILLCELL_X1 FILLER_103_1029 ();
 FILLCELL_X16 FILLER_103_1037 ();
 FILLCELL_X2 FILLER_103_1053 ();
 FILLCELL_X1 FILLER_103_1055 ();
 FILLCELL_X2 FILLER_103_1059 ();
 FILLCELL_X1 FILLER_103_1061 ();
 FILLCELL_X16 FILLER_103_1086 ();
 FILLCELL_X8 FILLER_103_1102 ();
 FILLCELL_X4 FILLER_103_1110 ();
 FILLCELL_X1 FILLER_103_1114 ();
 FILLCELL_X4 FILLER_103_1128 ();
 FILLCELL_X2 FILLER_103_1132 ();
 FILLCELL_X1 FILLER_103_1151 ();
 FILLCELL_X16 FILLER_103_1156 ();
 FILLCELL_X2 FILLER_103_1172 ();
 FILLCELL_X1 FILLER_103_1174 ();
 FILLCELL_X2 FILLER_103_1192 ();
 FILLCELL_X4 FILLER_103_1218 ();
 FILLCELL_X16 FILLER_104_1 ();
 FILLCELL_X8 FILLER_104_20 ();
 FILLCELL_X2 FILLER_104_28 ();
 FILLCELL_X1 FILLER_104_30 ();
 FILLCELL_X1 FILLER_104_48 ();
 FILLCELL_X8 FILLER_104_66 ();
 FILLCELL_X4 FILLER_104_74 ();
 FILLCELL_X1 FILLER_104_78 ();
 FILLCELL_X16 FILLER_104_89 ();
 FILLCELL_X1 FILLER_104_105 ();
 FILLCELL_X4 FILLER_104_110 ();
 FILLCELL_X32 FILLER_104_121 ();
 FILLCELL_X16 FILLER_104_153 ();
 FILLCELL_X8 FILLER_104_169 ();
 FILLCELL_X4 FILLER_104_177 ();
 FILLCELL_X1 FILLER_104_181 ();
 FILLCELL_X8 FILLER_104_189 ();
 FILLCELL_X1 FILLER_104_197 ();
 FILLCELL_X8 FILLER_104_205 ();
 FILLCELL_X1 FILLER_104_213 ();
 FILLCELL_X16 FILLER_104_217 ();
 FILLCELL_X8 FILLER_104_233 ();
 FILLCELL_X2 FILLER_104_241 ();
 FILLCELL_X16 FILLER_104_250 ();
 FILLCELL_X8 FILLER_104_266 ();
 FILLCELL_X1 FILLER_104_274 ();
 FILLCELL_X8 FILLER_104_292 ();
 FILLCELL_X2 FILLER_104_300 ();
 FILLCELL_X4 FILLER_104_319 ();
 FILLCELL_X32 FILLER_104_330 ();
 FILLCELL_X8 FILLER_104_366 ();
 FILLCELL_X2 FILLER_104_374 ();
 FILLCELL_X1 FILLER_104_376 ();
 FILLCELL_X8 FILLER_104_394 ();
 FILLCELL_X4 FILLER_104_402 ();
 FILLCELL_X1 FILLER_104_413 ();
 FILLCELL_X1 FILLER_104_421 ();
 FILLCELL_X8 FILLER_104_429 ();
 FILLCELL_X4 FILLER_104_437 ();
 FILLCELL_X2 FILLER_104_441 ();
 FILLCELL_X1 FILLER_104_443 ();
 FILLCELL_X4 FILLER_104_461 ();
 FILLCELL_X4 FILLER_104_472 ();
 FILLCELL_X2 FILLER_104_476 ();
 FILLCELL_X1 FILLER_104_478 ();
 FILLCELL_X16 FILLER_104_486 ();
 FILLCELL_X2 FILLER_104_502 ();
 FILLCELL_X2 FILLER_104_508 ();
 FILLCELL_X1 FILLER_104_510 ();
 FILLCELL_X16 FILLER_104_518 ();
 FILLCELL_X4 FILLER_104_534 ();
 FILLCELL_X2 FILLER_104_538 ();
 FILLCELL_X2 FILLER_104_558 ();
 FILLCELL_X8 FILLER_104_581 ();
 FILLCELL_X16 FILLER_104_606 ();
 FILLCELL_X8 FILLER_104_622 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X2 FILLER_104_632 ();
 FILLCELL_X1 FILLER_104_634 ();
 FILLCELL_X4 FILLER_104_652 ();
 FILLCELL_X1 FILLER_104_656 ();
 FILLCELL_X2 FILLER_104_713 ();
 FILLCELL_X4 FILLER_104_732 ();
 FILLCELL_X4 FILLER_104_743 ();
 FILLCELL_X2 FILLER_104_747 ();
 FILLCELL_X1 FILLER_104_749 ();
 FILLCELL_X4 FILLER_104_757 ();
 FILLCELL_X1 FILLER_104_761 ();
 FILLCELL_X2 FILLER_104_766 ();
 FILLCELL_X1 FILLER_104_779 ();
 FILLCELL_X16 FILLER_104_790 ();
 FILLCELL_X4 FILLER_104_806 ();
 FILLCELL_X1 FILLER_104_810 ();
 FILLCELL_X32 FILLER_104_821 ();
 FILLCELL_X1 FILLER_104_853 ();
 FILLCELL_X1 FILLER_104_863 ();
 FILLCELL_X4 FILLER_104_873 ();
 FILLCELL_X4 FILLER_104_884 ();
 FILLCELL_X1 FILLER_104_923 ();
 FILLCELL_X4 FILLER_104_930 ();
 FILLCELL_X1 FILLER_104_934 ();
 FILLCELL_X8 FILLER_104_942 ();
 FILLCELL_X4 FILLER_104_950 ();
 FILLCELL_X4 FILLER_104_989 ();
 FILLCELL_X1 FILLER_104_993 ();
 FILLCELL_X8 FILLER_104_1016 ();
 FILLCELL_X4 FILLER_104_1024 ();
 FILLCELL_X2 FILLER_104_1028 ();
 FILLCELL_X1 FILLER_104_1030 ();
 FILLCELL_X16 FILLER_104_1039 ();
 FILLCELL_X1 FILLER_104_1055 ();
 FILLCELL_X8 FILLER_104_1059 ();
 FILLCELL_X8 FILLER_104_1091 ();
 FILLCELL_X2 FILLER_104_1099 ();
 FILLCELL_X8 FILLER_104_1125 ();
 FILLCELL_X4 FILLER_104_1157 ();
 FILLCELL_X1 FILLER_104_1185 ();
 FILLCELL_X2 FILLER_104_1193 ();
 FILLCELL_X2 FILLER_104_1202 ();
 FILLCELL_X4 FILLER_104_1209 ();
 FILLCELL_X2 FILLER_104_1227 ();
 FILLCELL_X1 FILLER_104_1229 ();
 FILLCELL_X2 FILLER_104_1233 ();
 FILLCELL_X1 FILLER_104_1235 ();
 FILLCELL_X16 FILLER_105_1 ();
 FILLCELL_X8 FILLER_105_17 ();
 FILLCELL_X2 FILLER_105_25 ();
 FILLCELL_X1 FILLER_105_71 ();
 FILLCELL_X4 FILLER_105_89 ();
 FILLCELL_X2 FILLER_105_93 ();
 FILLCELL_X1 FILLER_105_95 ();
 FILLCELL_X1 FILLER_105_110 ();
 FILLCELL_X4 FILLER_105_118 ();
 FILLCELL_X1 FILLER_105_122 ();
 FILLCELL_X8 FILLER_105_130 ();
 FILLCELL_X1 FILLER_105_138 ();
 FILLCELL_X2 FILLER_105_146 ();
 FILLCELL_X1 FILLER_105_148 ();
 FILLCELL_X8 FILLER_105_163 ();
 FILLCELL_X4 FILLER_105_171 ();
 FILLCELL_X2 FILLER_105_175 ();
 FILLCELL_X16 FILLER_105_199 ();
 FILLCELL_X4 FILLER_105_215 ();
 FILLCELL_X2 FILLER_105_219 ();
 FILLCELL_X2 FILLER_105_228 ();
 FILLCELL_X1 FILLER_105_230 ();
 FILLCELL_X4 FILLER_105_238 ();
 FILLCELL_X2 FILLER_105_242 ();
 FILLCELL_X4 FILLER_105_261 ();
 FILLCELL_X2 FILLER_105_265 ();
 FILLCELL_X1 FILLER_105_291 ();
 FILLCELL_X16 FILLER_105_297 ();
 FILLCELL_X8 FILLER_105_313 ();
 FILLCELL_X2 FILLER_105_321 ();
 FILLCELL_X1 FILLER_105_323 ();
 FILLCELL_X32 FILLER_105_341 ();
 FILLCELL_X32 FILLER_105_373 ();
 FILLCELL_X8 FILLER_105_405 ();
 FILLCELL_X2 FILLER_105_413 ();
 FILLCELL_X4 FILLER_105_485 ();
 FILLCELL_X2 FILLER_105_522 ();
 FILLCELL_X1 FILLER_105_524 ();
 FILLCELL_X8 FILLER_105_536 ();
 FILLCELL_X4 FILLER_105_544 ();
 FILLCELL_X1 FILLER_105_548 ();
 FILLCELL_X1 FILLER_105_552 ();
 FILLCELL_X8 FILLER_105_570 ();
 FILLCELL_X4 FILLER_105_578 ();
 FILLCELL_X2 FILLER_105_582 ();
 FILLCELL_X1 FILLER_105_584 ();
 FILLCELL_X8 FILLER_105_616 ();
 FILLCELL_X4 FILLER_105_624 ();
 FILLCELL_X2 FILLER_105_628 ();
 FILLCELL_X4 FILLER_105_654 ();
 FILLCELL_X2 FILLER_105_658 ();
 FILLCELL_X1 FILLER_105_667 ();
 FILLCELL_X2 FILLER_105_675 ();
 FILLCELL_X1 FILLER_105_677 ();
 FILLCELL_X4 FILLER_105_689 ();
 FILLCELL_X2 FILLER_105_693 ();
 FILLCELL_X1 FILLER_105_729 ();
 FILLCELL_X2 FILLER_105_759 ();
 FILLCELL_X16 FILLER_105_783 ();
 FILLCELL_X4 FILLER_105_799 ();
 FILLCELL_X16 FILLER_105_822 ();
 FILLCELL_X8 FILLER_105_838 ();
 FILLCELL_X2 FILLER_105_846 ();
 FILLCELL_X1 FILLER_105_855 ();
 FILLCELL_X2 FILLER_105_865 ();
 FILLCELL_X4 FILLER_105_878 ();
 FILLCELL_X2 FILLER_105_882 ();
 FILLCELL_X1 FILLER_105_884 ();
 FILLCELL_X4 FILLER_105_887 ();
 FILLCELL_X1 FILLER_105_902 ();
 FILLCELL_X1 FILLER_105_923 ();
 FILLCELL_X1 FILLER_105_933 ();
 FILLCELL_X8 FILLER_105_939 ();
 FILLCELL_X2 FILLER_105_950 ();
 FILLCELL_X1 FILLER_105_952 ();
 FILLCELL_X4 FILLER_105_984 ();
 FILLCELL_X2 FILLER_105_988 ();
 FILLCELL_X2 FILLER_105_1000 ();
 FILLCELL_X1 FILLER_105_1002 ();
 FILLCELL_X8 FILLER_105_1007 ();
 FILLCELL_X2 FILLER_105_1015 ();
 FILLCELL_X1 FILLER_105_1017 ();
 FILLCELL_X1 FILLER_105_1028 ();
 FILLCELL_X32 FILLER_105_1047 ();
 FILLCELL_X16 FILLER_105_1079 ();
 FILLCELL_X1 FILLER_105_1095 ();
 FILLCELL_X8 FILLER_105_1127 ();
 FILLCELL_X2 FILLER_105_1149 ();
 FILLCELL_X2 FILLER_105_1165 ();
 FILLCELL_X1 FILLER_105_1181 ();
 FILLCELL_X2 FILLER_105_1213 ();
 FILLCELL_X2 FILLER_105_1232 ();
 FILLCELL_X2 FILLER_105_1237 ();
 FILLCELL_X1 FILLER_105_1239 ();
 FILLCELL_X16 FILLER_106_1 ();
 FILLCELL_X8 FILLER_106_17 ();
 FILLCELL_X4 FILLER_106_25 ();
 FILLCELL_X1 FILLER_106_50 ();
 FILLCELL_X2 FILLER_106_56 ();
 FILLCELL_X1 FILLER_106_65 ();
 FILLCELL_X4 FILLER_106_80 ();
 FILLCELL_X2 FILLER_106_91 ();
 FILLCELL_X1 FILLER_106_115 ();
 FILLCELL_X2 FILLER_106_123 ();
 FILLCELL_X2 FILLER_106_142 ();
 FILLCELL_X2 FILLER_106_161 ();
 FILLCELL_X16 FILLER_106_201 ();
 FILLCELL_X1 FILLER_106_217 ();
 FILLCELL_X4 FILLER_106_235 ();
 FILLCELL_X2 FILLER_106_239 ();
 FILLCELL_X8 FILLER_106_248 ();
 FILLCELL_X1 FILLER_106_263 ();
 FILLCELL_X4 FILLER_106_271 ();
 FILLCELL_X8 FILLER_106_299 ();
 FILLCELL_X16 FILLER_106_324 ();
 FILLCELL_X4 FILLER_106_340 ();
 FILLCELL_X4 FILLER_106_351 ();
 FILLCELL_X2 FILLER_106_355 ();
 FILLCELL_X1 FILLER_106_357 ();
 FILLCELL_X16 FILLER_106_365 ();
 FILLCELL_X4 FILLER_106_381 ();
 FILLCELL_X2 FILLER_106_385 ();
 FILLCELL_X2 FILLER_106_404 ();
 FILLCELL_X1 FILLER_106_406 ();
 FILLCELL_X1 FILLER_106_414 ();
 FILLCELL_X4 FILLER_106_446 ();
 FILLCELL_X16 FILLER_106_454 ();
 FILLCELL_X8 FILLER_106_470 ();
 FILLCELL_X4 FILLER_106_478 ();
 FILLCELL_X2 FILLER_106_482 ();
 FILLCELL_X1 FILLER_106_484 ();
 FILLCELL_X1 FILLER_106_492 ();
 FILLCELL_X2 FILLER_106_496 ();
 FILLCELL_X2 FILLER_106_505 ();
 FILLCELL_X4 FILLER_106_517 ();
 FILLCELL_X2 FILLER_106_545 ();
 FILLCELL_X16 FILLER_106_560 ();
 FILLCELL_X8 FILLER_106_576 ();
 FILLCELL_X2 FILLER_106_584 ();
 FILLCELL_X1 FILLER_106_586 ();
 FILLCELL_X4 FILLER_106_592 ();
 FILLCELL_X1 FILLER_106_596 ();
 FILLCELL_X8 FILLER_106_621 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X16 FILLER_106_652 ();
 FILLCELL_X1 FILLER_106_668 ();
 FILLCELL_X4 FILLER_106_726 ();
 FILLCELL_X1 FILLER_106_730 ();
 FILLCELL_X8 FILLER_106_734 ();
 FILLCELL_X2 FILLER_106_742 ();
 FILLCELL_X16 FILLER_106_780 ();
 FILLCELL_X4 FILLER_106_796 ();
 FILLCELL_X2 FILLER_106_800 ();
 FILLCELL_X16 FILLER_106_828 ();
 FILLCELL_X8 FILLER_106_844 ();
 FILLCELL_X4 FILLER_106_852 ();
 FILLCELL_X2 FILLER_106_856 ();
 FILLCELL_X16 FILLER_106_876 ();
 FILLCELL_X1 FILLER_106_913 ();
 FILLCELL_X1 FILLER_106_927 ();
 FILLCELL_X1 FILLER_106_931 ();
 FILLCELL_X4 FILLER_106_951 ();
 FILLCELL_X1 FILLER_106_955 ();
 FILLCELL_X2 FILLER_106_960 ();
 FILLCELL_X1 FILLER_106_965 ();
 FILLCELL_X1 FILLER_106_971 ();
 FILLCELL_X8 FILLER_106_974 ();
 FILLCELL_X2 FILLER_106_982 ();
 FILLCELL_X1 FILLER_106_984 ();
 FILLCELL_X8 FILLER_106_1007 ();
 FILLCELL_X1 FILLER_106_1015 ();
 FILLCELL_X16 FILLER_106_1032 ();
 FILLCELL_X8 FILLER_106_1048 ();
 FILLCELL_X4 FILLER_106_1056 ();
 FILLCELL_X8 FILLER_106_1062 ();
 FILLCELL_X1 FILLER_106_1070 ();
 FILLCELL_X32 FILLER_106_1074 ();
 FILLCELL_X8 FILLER_106_1106 ();
 FILLCELL_X2 FILLER_106_1114 ();
 FILLCELL_X1 FILLER_106_1116 ();
 FILLCELL_X4 FILLER_106_1124 ();
 FILLCELL_X2 FILLER_106_1141 ();
 FILLCELL_X1 FILLER_106_1143 ();
 FILLCELL_X2 FILLER_106_1151 ();
 FILLCELL_X8 FILLER_106_1192 ();
 FILLCELL_X2 FILLER_106_1200 ();
 FILLCELL_X1 FILLER_106_1202 ();
 FILLCELL_X1 FILLER_106_1219 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X16 FILLER_107_33 ();
 FILLCELL_X8 FILLER_107_49 ();
 FILLCELL_X1 FILLER_107_64 ();
 FILLCELL_X2 FILLER_107_82 ();
 FILLCELL_X2 FILLER_107_91 ();
 FILLCELL_X2 FILLER_107_100 ();
 FILLCELL_X1 FILLER_107_119 ();
 FILLCELL_X4 FILLER_107_146 ();
 FILLCELL_X2 FILLER_107_150 ();
 FILLCELL_X1 FILLER_107_169 ();
 FILLCELL_X1 FILLER_107_177 ();
 FILLCELL_X2 FILLER_107_195 ();
 FILLCELL_X1 FILLER_107_204 ();
 FILLCELL_X2 FILLER_107_222 ();
 FILLCELL_X4 FILLER_107_241 ();
 FILLCELL_X1 FILLER_107_245 ();
 FILLCELL_X4 FILLER_107_274 ();
 FILLCELL_X4 FILLER_107_285 ();
 FILLCELL_X2 FILLER_107_289 ();
 FILLCELL_X2 FILLER_107_329 ();
 FILLCELL_X1 FILLER_107_331 ();
 FILLCELL_X2 FILLER_107_346 ();
 FILLCELL_X1 FILLER_107_357 ();
 FILLCELL_X16 FILLER_107_365 ();
 FILLCELL_X1 FILLER_107_381 ();
 FILLCELL_X8 FILLER_107_415 ();
 FILLCELL_X1 FILLER_107_423 ();
 FILLCELL_X4 FILLER_107_453 ();
 FILLCELL_X2 FILLER_107_457 ();
 FILLCELL_X2 FILLER_107_483 ();
 FILLCELL_X1 FILLER_107_485 ();
 FILLCELL_X4 FILLER_107_493 ();
 FILLCELL_X1 FILLER_107_497 ();
 FILLCELL_X2 FILLER_107_515 ();
 FILLCELL_X2 FILLER_107_524 ();
 FILLCELL_X4 FILLER_107_543 ();
 FILLCELL_X1 FILLER_107_547 ();
 FILLCELL_X4 FILLER_107_562 ();
 FILLCELL_X2 FILLER_107_573 ();
 FILLCELL_X16 FILLER_107_582 ();
 FILLCELL_X4 FILLER_107_598 ();
 FILLCELL_X2 FILLER_107_616 ();
 FILLCELL_X1 FILLER_107_618 ();
 FILLCELL_X4 FILLER_107_626 ();
 FILLCELL_X2 FILLER_107_630 ();
 FILLCELL_X1 FILLER_107_632 ();
 FILLCELL_X8 FILLER_107_637 ();
 FILLCELL_X4 FILLER_107_658 ();
 FILLCELL_X2 FILLER_107_662 ();
 FILLCELL_X2 FILLER_107_695 ();
 FILLCELL_X1 FILLER_107_697 ();
 FILLCELL_X8 FILLER_107_702 ();
 FILLCELL_X2 FILLER_107_710 ();
 FILLCELL_X2 FILLER_107_740 ();
 FILLCELL_X1 FILLER_107_742 ();
 FILLCELL_X8 FILLER_107_747 ();
 FILLCELL_X1 FILLER_107_755 ();
 FILLCELL_X8 FILLER_107_760 ();
 FILLCELL_X4 FILLER_107_768 ();
 FILLCELL_X32 FILLER_107_774 ();
 FILLCELL_X2 FILLER_107_806 ();
 FILLCELL_X1 FILLER_107_808 ();
 FILLCELL_X2 FILLER_107_821 ();
 FILLCELL_X1 FILLER_107_823 ();
 FILLCELL_X2 FILLER_107_833 ();
 FILLCELL_X1 FILLER_107_835 ();
 FILLCELL_X8 FILLER_107_845 ();
 FILLCELL_X2 FILLER_107_853 ();
 FILLCELL_X1 FILLER_107_855 ();
 FILLCELL_X4 FILLER_107_859 ();
 FILLCELL_X2 FILLER_107_863 ();
 FILLCELL_X4 FILLER_107_882 ();
 FILLCELL_X2 FILLER_107_886 ();
 FILLCELL_X1 FILLER_107_888 ();
 FILLCELL_X4 FILLER_107_900 ();
 FILLCELL_X2 FILLER_107_904 ();
 FILLCELL_X1 FILLER_107_906 ();
 FILLCELL_X1 FILLER_107_910 ();
 FILLCELL_X1 FILLER_107_914 ();
 FILLCELL_X1 FILLER_107_922 ();
 FILLCELL_X2 FILLER_107_947 ();
 FILLCELL_X1 FILLER_107_949 ();
 FILLCELL_X16 FILLER_107_955 ();
 FILLCELL_X8 FILLER_107_971 ();
 FILLCELL_X4 FILLER_107_979 ();
 FILLCELL_X1 FILLER_107_983 ();
 FILLCELL_X2 FILLER_107_1003 ();
 FILLCELL_X1 FILLER_107_1016 ();
 FILLCELL_X8 FILLER_107_1020 ();
 FILLCELL_X8 FILLER_107_1044 ();
 FILLCELL_X4 FILLER_107_1052 ();
 FILLCELL_X32 FILLER_107_1068 ();
 FILLCELL_X4 FILLER_107_1100 ();
 FILLCELL_X2 FILLER_107_1128 ();
 FILLCELL_X1 FILLER_107_1130 ();
 FILLCELL_X16 FILLER_107_1155 ();
 FILLCELL_X1 FILLER_107_1171 ();
 FILLCELL_X8 FILLER_107_1179 ();
 FILLCELL_X2 FILLER_107_1187 ();
 FILLCELL_X4 FILLER_107_1227 ();
 FILLCELL_X2 FILLER_107_1231 ();
 FILLCELL_X1 FILLER_107_1236 ();
 FILLCELL_X16 FILLER_108_1 ();
 FILLCELL_X2 FILLER_108_17 ();
 FILLCELL_X1 FILLER_108_19 ();
 FILLCELL_X2 FILLER_108_44 ();
 FILLCELL_X32 FILLER_108_53 ();
 FILLCELL_X16 FILLER_108_85 ();
 FILLCELL_X2 FILLER_108_101 ();
 FILLCELL_X1 FILLER_108_103 ();
 FILLCELL_X16 FILLER_108_107 ();
 FILLCELL_X8 FILLER_108_123 ();
 FILLCELL_X4 FILLER_108_131 ();
 FILLCELL_X1 FILLER_108_135 ();
 FILLCELL_X4 FILLER_108_143 ();
 FILLCELL_X1 FILLER_108_147 ();
 FILLCELL_X8 FILLER_108_183 ();
 FILLCELL_X2 FILLER_108_191 ();
 FILLCELL_X2 FILLER_108_200 ();
 FILLCELL_X1 FILLER_108_202 ();
 FILLCELL_X8 FILLER_108_210 ();
 FILLCELL_X4 FILLER_108_218 ();
 FILLCELL_X1 FILLER_108_222 ();
 FILLCELL_X8 FILLER_108_230 ();
 FILLCELL_X4 FILLER_108_238 ();
 FILLCELL_X4 FILLER_108_247 ();
 FILLCELL_X2 FILLER_108_251 ();
 FILLCELL_X1 FILLER_108_253 ();
 FILLCELL_X2 FILLER_108_261 ();
 FILLCELL_X1 FILLER_108_263 ();
 FILLCELL_X16 FILLER_108_281 ();
 FILLCELL_X8 FILLER_108_297 ();
 FILLCELL_X4 FILLER_108_305 ();
 FILLCELL_X2 FILLER_108_309 ();
 FILLCELL_X4 FILLER_108_325 ();
 FILLCELL_X2 FILLER_108_329 ();
 FILLCELL_X1 FILLER_108_331 ();
 FILLCELL_X2 FILLER_108_349 ();
 FILLCELL_X8 FILLER_108_382 ();
 FILLCELL_X1 FILLER_108_390 ();
 FILLCELL_X32 FILLER_108_414 ();
 FILLCELL_X32 FILLER_108_446 ();
 FILLCELL_X8 FILLER_108_478 ();
 FILLCELL_X2 FILLER_108_486 ();
 FILLCELL_X8 FILLER_108_505 ();
 FILLCELL_X4 FILLER_108_513 ();
 FILLCELL_X8 FILLER_108_524 ();
 FILLCELL_X8 FILLER_108_540 ();
 FILLCELL_X1 FILLER_108_548 ();
 FILLCELL_X8 FILLER_108_552 ();
 FILLCELL_X4 FILLER_108_560 ();
 FILLCELL_X1 FILLER_108_588 ();
 FILLCELL_X4 FILLER_108_605 ();
 FILLCELL_X1 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_627 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X16 FILLER_108_664 ();
 FILLCELL_X8 FILLER_108_680 ();
 FILLCELL_X4 FILLER_108_691 ();
 FILLCELL_X1 FILLER_108_695 ();
 FILLCELL_X8 FILLER_108_701 ();
 FILLCELL_X4 FILLER_108_709 ();
 FILLCELL_X2 FILLER_108_730 ();
 FILLCELL_X2 FILLER_108_739 ();
 FILLCELL_X1 FILLER_108_741 ();
 FILLCELL_X2 FILLER_108_749 ();
 FILLCELL_X1 FILLER_108_751 ();
 FILLCELL_X16 FILLER_108_776 ();
 FILLCELL_X8 FILLER_108_792 ();
 FILLCELL_X4 FILLER_108_800 ();
 FILLCELL_X1 FILLER_108_804 ();
 FILLCELL_X32 FILLER_108_827 ();
 FILLCELL_X16 FILLER_108_859 ();
 FILLCELL_X2 FILLER_108_875 ();
 FILLCELL_X1 FILLER_108_877 ();
 FILLCELL_X16 FILLER_108_882 ();
 FILLCELL_X4 FILLER_108_898 ();
 FILLCELL_X1 FILLER_108_902 ();
 FILLCELL_X4 FILLER_108_916 ();
 FILLCELL_X4 FILLER_108_926 ();
 FILLCELL_X1 FILLER_108_930 ();
 FILLCELL_X8 FILLER_108_938 ();
 FILLCELL_X8 FILLER_108_950 ();
 FILLCELL_X2 FILLER_108_958 ();
 FILLCELL_X1 FILLER_108_960 ();
 FILLCELL_X2 FILLER_108_965 ();
 FILLCELL_X1 FILLER_108_967 ();
 FILLCELL_X8 FILLER_108_973 ();
 FILLCELL_X2 FILLER_108_1009 ();
 FILLCELL_X1 FILLER_108_1014 ();
 FILLCELL_X4 FILLER_108_1024 ();
 FILLCELL_X2 FILLER_108_1028 ();
 FILLCELL_X2 FILLER_108_1039 ();
 FILLCELL_X1 FILLER_108_1058 ();
 FILLCELL_X16 FILLER_108_1072 ();
 FILLCELL_X8 FILLER_108_1088 ();
 FILLCELL_X4 FILLER_108_1096 ();
 FILLCELL_X2 FILLER_108_1100 ();
 FILLCELL_X1 FILLER_108_1119 ();
 FILLCELL_X4 FILLER_108_1127 ();
 FILLCELL_X1 FILLER_108_1131 ();
 FILLCELL_X32 FILLER_108_1156 ();
 FILLCELL_X2 FILLER_108_1188 ();
 FILLCELL_X1 FILLER_108_1190 ();
 FILLCELL_X1 FILLER_108_1215 ();
 FILLCELL_X1 FILLER_108_1236 ();
 FILLCELL_X16 FILLER_109_1 ();
 FILLCELL_X8 FILLER_109_17 ();
 FILLCELL_X4 FILLER_109_25 ();
 FILLCELL_X2 FILLER_109_29 ();
 FILLCELL_X1 FILLER_109_31 ();
 FILLCELL_X32 FILLER_109_56 ();
 FILLCELL_X32 FILLER_109_88 ();
 FILLCELL_X32 FILLER_109_120 ();
 FILLCELL_X8 FILLER_109_152 ();
 FILLCELL_X4 FILLER_109_160 ();
 FILLCELL_X1 FILLER_109_164 ();
 FILLCELL_X32 FILLER_109_168 ();
 FILLCELL_X32 FILLER_109_200 ();
 FILLCELL_X16 FILLER_109_232 ();
 FILLCELL_X4 FILLER_109_248 ();
 FILLCELL_X2 FILLER_109_252 ();
 FILLCELL_X8 FILLER_109_285 ();
 FILLCELL_X2 FILLER_109_293 ();
 FILLCELL_X1 FILLER_109_295 ();
 FILLCELL_X1 FILLER_109_320 ();
 FILLCELL_X2 FILLER_109_328 ();
 FILLCELL_X8 FILLER_109_335 ();
 FILLCELL_X2 FILLER_109_343 ();
 FILLCELL_X2 FILLER_109_352 ();
 FILLCELL_X32 FILLER_109_361 ();
 FILLCELL_X4 FILLER_109_410 ();
 FILLCELL_X16 FILLER_109_418 ();
 FILLCELL_X8 FILLER_109_434 ();
 FILLCELL_X1 FILLER_109_442 ();
 FILLCELL_X4 FILLER_109_474 ();
 FILLCELL_X8 FILLER_109_493 ();
 FILLCELL_X2 FILLER_109_501 ();
 FILLCELL_X8 FILLER_109_514 ();
 FILLCELL_X1 FILLER_109_522 ();
 FILLCELL_X16 FILLER_109_540 ();
 FILLCELL_X1 FILLER_109_556 ();
 FILLCELL_X32 FILLER_109_591 ();
 FILLCELL_X8 FILLER_109_623 ();
 FILLCELL_X4 FILLER_109_631 ();
 FILLCELL_X1 FILLER_109_635 ();
 FILLCELL_X8 FILLER_109_640 ();
 FILLCELL_X2 FILLER_109_687 ();
 FILLCELL_X4 FILLER_109_714 ();
 FILLCELL_X2 FILLER_109_718 ();
 FILLCELL_X4 FILLER_109_727 ();
 FILLCELL_X2 FILLER_109_731 ();
 FILLCELL_X1 FILLER_109_733 ();
 FILLCELL_X32 FILLER_109_758 ();
 FILLCELL_X32 FILLER_109_790 ();
 FILLCELL_X32 FILLER_109_822 ();
 FILLCELL_X4 FILLER_109_854 ();
 FILLCELL_X1 FILLER_109_858 ();
 FILLCELL_X16 FILLER_109_879 ();
 FILLCELL_X8 FILLER_109_895 ();
 FILLCELL_X4 FILLER_109_919 ();
 FILLCELL_X1 FILLER_109_923 ();
 FILLCELL_X16 FILLER_109_927 ();
 FILLCELL_X2 FILLER_109_946 ();
 FILLCELL_X1 FILLER_109_948 ();
 FILLCELL_X1 FILLER_109_956 ();
 FILLCELL_X8 FILLER_109_1019 ();
 FILLCELL_X2 FILLER_109_1027 ();
 FILLCELL_X16 FILLER_109_1086 ();
 FILLCELL_X4 FILLER_109_1102 ();
 FILLCELL_X1 FILLER_109_1106 ();
 FILLCELL_X2 FILLER_109_1133 ();
 FILLCELL_X32 FILLER_109_1142 ();
 FILLCELL_X2 FILLER_109_1174 ();
 FILLCELL_X1 FILLER_109_1176 ();
 FILLCELL_X1 FILLER_109_1201 ();
 FILLCELL_X1 FILLER_109_1209 ();
 FILLCELL_X2 FILLER_109_1227 ();
 FILLCELL_X1 FILLER_109_1229 ();
 FILLCELL_X2 FILLER_109_1233 ();
 FILLCELL_X1 FILLER_109_1235 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X16 FILLER_110_33 ();
 FILLCELL_X8 FILLER_110_49 ();
 FILLCELL_X2 FILLER_110_74 ();
 FILLCELL_X1 FILLER_110_76 ();
 FILLCELL_X1 FILLER_110_101 ();
 FILLCELL_X4 FILLER_110_119 ();
 FILLCELL_X2 FILLER_110_123 ();
 FILLCELL_X16 FILLER_110_142 ();
 FILLCELL_X4 FILLER_110_158 ();
 FILLCELL_X2 FILLER_110_162 ();
 FILLCELL_X32 FILLER_110_195 ();
 FILLCELL_X32 FILLER_110_227 ();
 FILLCELL_X16 FILLER_110_259 ();
 FILLCELL_X2 FILLER_110_275 ();
 FILLCELL_X1 FILLER_110_277 ();
 FILLCELL_X8 FILLER_110_295 ();
 FILLCELL_X4 FILLER_110_303 ();
 FILLCELL_X1 FILLER_110_307 ();
 FILLCELL_X16 FILLER_110_315 ();
 FILLCELL_X4 FILLER_110_331 ();
 FILLCELL_X1 FILLER_110_335 ();
 FILLCELL_X2 FILLER_110_353 ();
 FILLCELL_X1 FILLER_110_355 ();
 FILLCELL_X32 FILLER_110_373 ();
 FILLCELL_X8 FILLER_110_405 ();
 FILLCELL_X4 FILLER_110_413 ();
 FILLCELL_X2 FILLER_110_417 ();
 FILLCELL_X16 FILLER_110_433 ();
 FILLCELL_X2 FILLER_110_449 ();
 FILLCELL_X8 FILLER_110_458 ();
 FILLCELL_X2 FILLER_110_466 ();
 FILLCELL_X4 FILLER_110_475 ();
 FILLCELL_X2 FILLER_110_479 ();
 FILLCELL_X1 FILLER_110_481 ();
 FILLCELL_X2 FILLER_110_489 ();
 FILLCELL_X8 FILLER_110_512 ();
 FILLCELL_X2 FILLER_110_520 ();
 FILLCELL_X8 FILLER_110_546 ();
 FILLCELL_X2 FILLER_110_554 ();
 FILLCELL_X1 FILLER_110_556 ();
 FILLCELL_X1 FILLER_110_564 ();
 FILLCELL_X16 FILLER_110_589 ();
 FILLCELL_X2 FILLER_110_612 ();
 FILLCELL_X2 FILLER_110_621 ();
 FILLCELL_X1 FILLER_110_630 ();
 FILLCELL_X1 FILLER_110_632 ();
 FILLCELL_X2 FILLER_110_646 ();
 FILLCELL_X4 FILLER_110_679 ();
 FILLCELL_X2 FILLER_110_683 ();
 FILLCELL_X4 FILLER_110_716 ();
 FILLCELL_X2 FILLER_110_720 ();
 FILLCELL_X1 FILLER_110_722 ();
 FILLCELL_X16 FILLER_110_747 ();
 FILLCELL_X8 FILLER_110_763 ();
 FILLCELL_X2 FILLER_110_771 ();
 FILLCELL_X32 FILLER_110_776 ();
 FILLCELL_X16 FILLER_110_808 ();
 FILLCELL_X8 FILLER_110_824 ();
 FILLCELL_X2 FILLER_110_832 ();
 FILLCELL_X8 FILLER_110_837 ();
 FILLCELL_X4 FILLER_110_845 ();
 FILLCELL_X8 FILLER_110_873 ();
 FILLCELL_X2 FILLER_110_881 ();
 FILLCELL_X2 FILLER_110_898 ();
 FILLCELL_X4 FILLER_110_938 ();
 FILLCELL_X2 FILLER_110_942 ();
 FILLCELL_X16 FILLER_110_1002 ();
 FILLCELL_X4 FILLER_110_1018 ();
 FILLCELL_X1 FILLER_110_1022 ();
 FILLCELL_X2 FILLER_110_1047 ();
 FILLCELL_X1 FILLER_110_1049 ();
 FILLCELL_X2 FILLER_110_1064 ();
 FILLCELL_X16 FILLER_110_1088 ();
 FILLCELL_X2 FILLER_110_1104 ();
 FILLCELL_X16 FILLER_110_1154 ();
 FILLCELL_X8 FILLER_110_1170 ();
 FILLCELL_X4 FILLER_110_1178 ();
 FILLCELL_X2 FILLER_110_1182 ();
 FILLCELL_X2 FILLER_110_1198 ();
 FILLCELL_X2 FILLER_110_1217 ();
 FILLCELL_X2 FILLER_110_1222 ();
 FILLCELL_X1 FILLER_110_1224 ();
 FILLCELL_X8 FILLER_110_1228 ();
 FILLCELL_X4 FILLER_110_1236 ();
 FILLCELL_X32 FILLER_111_5 ();
 FILLCELL_X8 FILLER_111_37 ();
 FILLCELL_X1 FILLER_111_45 ();
 FILLCELL_X4 FILLER_111_63 ();
 FILLCELL_X2 FILLER_111_67 ();
 FILLCELL_X1 FILLER_111_69 ();
 FILLCELL_X4 FILLER_111_77 ();
 FILLCELL_X4 FILLER_111_95 ();
 FILLCELL_X1 FILLER_111_99 ();
 FILLCELL_X8 FILLER_111_117 ();
 FILLCELL_X8 FILLER_111_149 ();
 FILLCELL_X2 FILLER_111_157 ();
 FILLCELL_X1 FILLER_111_159 ();
 FILLCELL_X2 FILLER_111_177 ();
 FILLCELL_X1 FILLER_111_179 ();
 FILLCELL_X16 FILLER_111_211 ();
 FILLCELL_X8 FILLER_111_227 ();
 FILLCELL_X4 FILLER_111_259 ();
 FILLCELL_X2 FILLER_111_263 ();
 FILLCELL_X1 FILLER_111_265 ();
 FILLCELL_X4 FILLER_111_273 ();
 FILLCELL_X2 FILLER_111_277 ();
 FILLCELL_X1 FILLER_111_279 ();
 FILLCELL_X16 FILLER_111_285 ();
 FILLCELL_X4 FILLER_111_301 ();
 FILLCELL_X2 FILLER_111_305 ();
 FILLCELL_X32 FILLER_111_331 ();
 FILLCELL_X8 FILLER_111_387 ();
 FILLCELL_X4 FILLER_111_395 ();
 FILLCELL_X8 FILLER_111_406 ();
 FILLCELL_X1 FILLER_111_414 ();
 FILLCELL_X4 FILLER_111_432 ();
 FILLCELL_X1 FILLER_111_436 ();
 FILLCELL_X1 FILLER_111_445 ();
 FILLCELL_X2 FILLER_111_463 ();
 FILLCELL_X1 FILLER_111_465 ();
 FILLCELL_X8 FILLER_111_493 ();
 FILLCELL_X4 FILLER_111_501 ();
 FILLCELL_X2 FILLER_111_505 ();
 FILLCELL_X2 FILLER_111_521 ();
 FILLCELL_X1 FILLER_111_523 ();
 FILLCELL_X16 FILLER_111_548 ();
 FILLCELL_X8 FILLER_111_564 ();
 FILLCELL_X1 FILLER_111_572 ();
 FILLCELL_X16 FILLER_111_580 ();
 FILLCELL_X4 FILLER_111_596 ();
 FILLCELL_X1 FILLER_111_617 ();
 FILLCELL_X1 FILLER_111_635 ();
 FILLCELL_X2 FILLER_111_667 ();
 FILLCELL_X1 FILLER_111_669 ();
 FILLCELL_X16 FILLER_111_704 ();
 FILLCELL_X8 FILLER_111_720 ();
 FILLCELL_X1 FILLER_111_728 ();
 FILLCELL_X1 FILLER_111_736 ();
 FILLCELL_X32 FILLER_111_744 ();
 FILLCELL_X32 FILLER_111_776 ();
 FILLCELL_X2 FILLER_111_808 ();
 FILLCELL_X2 FILLER_111_817 ();
 FILLCELL_X1 FILLER_111_819 ();
 FILLCELL_X1 FILLER_111_827 ();
 FILLCELL_X2 FILLER_111_841 ();
 FILLCELL_X1 FILLER_111_843 ();
 FILLCELL_X1 FILLER_111_856 ();
 FILLCELL_X2 FILLER_111_866 ();
 FILLCELL_X1 FILLER_111_886 ();
 FILLCELL_X2 FILLER_111_898 ();
 FILLCELL_X1 FILLER_111_900 ();
 FILLCELL_X2 FILLER_111_929 ();
 FILLCELL_X2 FILLER_111_938 ();
 FILLCELL_X1 FILLER_111_946 ();
 FILLCELL_X1 FILLER_111_953 ();
 FILLCELL_X1 FILLER_111_976 ();
 FILLCELL_X1 FILLER_111_1005 ();
 FILLCELL_X4 FILLER_111_1010 ();
 FILLCELL_X2 FILLER_111_1014 ();
 FILLCELL_X1 FILLER_111_1016 ();
 FILLCELL_X1 FILLER_111_1020 ();
 FILLCELL_X1 FILLER_111_1066 ();
 FILLCELL_X1 FILLER_111_1080 ();
 FILLCELL_X8 FILLER_111_1087 ();
 FILLCELL_X1 FILLER_111_1095 ();
 FILLCELL_X8 FILLER_111_1101 ();
 FILLCELL_X2 FILLER_111_1109 ();
 FILLCELL_X1 FILLER_111_1111 ();
 FILLCELL_X16 FILLER_111_1156 ();
 FILLCELL_X2 FILLER_111_1172 ();
 FILLCELL_X4 FILLER_111_1225 ();
 FILLCELL_X1 FILLER_111_1236 ();
 FILLCELL_X16 FILLER_112_1 ();
 FILLCELL_X4 FILLER_112_17 ();
 FILLCELL_X8 FILLER_112_38 ();
 FILLCELL_X1 FILLER_112_46 ();
 FILLCELL_X32 FILLER_112_59 ();
 FILLCELL_X4 FILLER_112_91 ();
 FILLCELL_X1 FILLER_112_95 ();
 FILLCELL_X2 FILLER_112_103 ();
 FILLCELL_X2 FILLER_112_122 ();
 FILLCELL_X1 FILLER_112_124 ();
 FILLCELL_X1 FILLER_112_132 ();
 FILLCELL_X2 FILLER_112_140 ();
 FILLCELL_X1 FILLER_112_142 ();
 FILLCELL_X2 FILLER_112_155 ();
 FILLCELL_X2 FILLER_112_181 ();
 FILLCELL_X1 FILLER_112_190 ();
 FILLCELL_X4 FILLER_112_225 ();
 FILLCELL_X2 FILLER_112_229 ();
 FILLCELL_X1 FILLER_112_231 ();
 FILLCELL_X8 FILLER_112_249 ();
 FILLCELL_X4 FILLER_112_257 ();
 FILLCELL_X1 FILLER_112_261 ();
 FILLCELL_X4 FILLER_112_296 ();
 FILLCELL_X4 FILLER_112_307 ();
 FILLCELL_X8 FILLER_112_335 ();
 FILLCELL_X1 FILLER_112_343 ();
 FILLCELL_X8 FILLER_112_351 ();
 FILLCELL_X1 FILLER_112_359 ();
 FILLCELL_X2 FILLER_112_371 ();
 FILLCELL_X1 FILLER_112_373 ();
 FILLCELL_X4 FILLER_112_391 ();
 FILLCELL_X1 FILLER_112_412 ();
 FILLCELL_X4 FILLER_112_444 ();
 FILLCELL_X1 FILLER_112_448 ();
 FILLCELL_X8 FILLER_112_456 ();
 FILLCELL_X4 FILLER_112_464 ();
 FILLCELL_X1 FILLER_112_485 ();
 FILLCELL_X2 FILLER_112_525 ();
 FILLCELL_X1 FILLER_112_527 ();
 FILLCELL_X8 FILLER_112_535 ();
 FILLCELL_X4 FILLER_112_543 ();
 FILLCELL_X2 FILLER_112_547 ();
 FILLCELL_X4 FILLER_112_574 ();
 FILLCELL_X2 FILLER_112_578 ();
 FILLCELL_X1 FILLER_112_580 ();
 FILLCELL_X16 FILLER_112_586 ();
 FILLCELL_X2 FILLER_112_602 ();
 FILLCELL_X8 FILLER_112_611 ();
 FILLCELL_X2 FILLER_112_619 ();
 FILLCELL_X2 FILLER_112_628 ();
 FILLCELL_X1 FILLER_112_630 ();
 FILLCELL_X32 FILLER_112_639 ();
 FILLCELL_X8 FILLER_112_671 ();
 FILLCELL_X1 FILLER_112_679 ();
 FILLCELL_X4 FILLER_112_711 ();
 FILLCELL_X2 FILLER_112_722 ();
 FILLCELL_X1 FILLER_112_724 ();
 FILLCELL_X8 FILLER_112_744 ();
 FILLCELL_X4 FILLER_112_752 ();
 FILLCELL_X4 FILLER_112_781 ();
 FILLCELL_X1 FILLER_112_785 ();
 FILLCELL_X4 FILLER_112_798 ();
 FILLCELL_X2 FILLER_112_802 ();
 FILLCELL_X2 FILLER_112_811 ();
 FILLCELL_X1 FILLER_112_813 ();
 FILLCELL_X2 FILLER_112_820 ();
 FILLCELL_X2 FILLER_112_832 ();
 FILLCELL_X1 FILLER_112_834 ();
 FILLCELL_X2 FILLER_112_849 ();
 FILLCELL_X2 FILLER_112_867 ();
 FILLCELL_X16 FILLER_112_891 ();
 FILLCELL_X1 FILLER_112_907 ();
 FILLCELL_X1 FILLER_112_921 ();
 FILLCELL_X1 FILLER_112_925 ();
 FILLCELL_X1 FILLER_112_939 ();
 FILLCELL_X1 FILLER_112_945 ();
 FILLCELL_X8 FILLER_112_973 ();
 FILLCELL_X2 FILLER_112_981 ();
 FILLCELL_X4 FILLER_112_1017 ();
 FILLCELL_X2 FILLER_112_1021 ();
 FILLCELL_X1 FILLER_112_1023 ();
 FILLCELL_X4 FILLER_112_1036 ();
 FILLCELL_X1 FILLER_112_1047 ();
 FILLCELL_X8 FILLER_112_1052 ();
 FILLCELL_X4 FILLER_112_1069 ();
 FILLCELL_X1 FILLER_112_1073 ();
 FILLCELL_X32 FILLER_112_1092 ();
 FILLCELL_X4 FILLER_112_1129 ();
 FILLCELL_X1 FILLER_112_1133 ();
 FILLCELL_X16 FILLER_112_1138 ();
 FILLCELL_X8 FILLER_112_1154 ();
 FILLCELL_X4 FILLER_112_1162 ();
 FILLCELL_X2 FILLER_112_1238 ();
 FILLCELL_X2 FILLER_113_1 ();
 FILLCELL_X4 FILLER_113_34 ();
 FILLCELL_X32 FILLER_113_71 ();
 FILLCELL_X4 FILLER_113_103 ();
 FILLCELL_X4 FILLER_113_114 ();
 FILLCELL_X4 FILLER_113_130 ();
 FILLCELL_X2 FILLER_113_134 ();
 FILLCELL_X1 FILLER_113_136 ();
 FILLCELL_X1 FILLER_113_168 ();
 FILLCELL_X8 FILLER_113_176 ();
 FILLCELL_X1 FILLER_113_184 ();
 FILLCELL_X8 FILLER_113_192 ();
 FILLCELL_X16 FILLER_113_214 ();
 FILLCELL_X4 FILLER_113_230 ();
 FILLCELL_X1 FILLER_113_234 ();
 FILLCELL_X4 FILLER_113_249 ();
 FILLCELL_X2 FILLER_113_253 ();
 FILLCELL_X4 FILLER_113_293 ();
 FILLCELL_X16 FILLER_113_321 ();
 FILLCELL_X4 FILLER_113_337 ();
 FILLCELL_X1 FILLER_113_341 ();
 FILLCELL_X16 FILLER_113_373 ();
 FILLCELL_X16 FILLER_113_393 ();
 FILLCELL_X8 FILLER_113_409 ();
 FILLCELL_X4 FILLER_113_417 ();
 FILLCELL_X16 FILLER_113_445 ();
 FILLCELL_X4 FILLER_113_461 ();
 FILLCELL_X2 FILLER_113_465 ();
 FILLCELL_X1 FILLER_113_467 ();
 FILLCELL_X8 FILLER_113_479 ();
 FILLCELL_X4 FILLER_113_487 ();
 FILLCELL_X8 FILLER_113_498 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X16 FILLER_113_545 ();
 FILLCELL_X4 FILLER_113_561 ();
 FILLCELL_X1 FILLER_113_565 ();
 FILLCELL_X1 FILLER_113_573 ();
 FILLCELL_X8 FILLER_113_593 ();
 FILLCELL_X16 FILLER_113_618 ();
 FILLCELL_X8 FILLER_113_634 ();
 FILLCELL_X4 FILLER_113_642 ();
 FILLCELL_X2 FILLER_113_646 ();
 FILLCELL_X8 FILLER_113_655 ();
 FILLCELL_X4 FILLER_113_663 ();
 FILLCELL_X4 FILLER_113_716 ();
 FILLCELL_X2 FILLER_113_720 ();
 FILLCELL_X4 FILLER_113_753 ();
 FILLCELL_X1 FILLER_113_785 ();
 FILLCELL_X8 FILLER_113_802 ();
 FILLCELL_X1 FILLER_113_827 ();
 FILLCELL_X2 FILLER_113_835 ();
 FILLCELL_X2 FILLER_113_844 ();
 FILLCELL_X1 FILLER_113_846 ();
 FILLCELL_X1 FILLER_113_857 ();
 FILLCELL_X2 FILLER_113_875 ();
 FILLCELL_X16 FILLER_113_881 ();
 FILLCELL_X8 FILLER_113_897 ();
 FILLCELL_X1 FILLER_113_905 ();
 FILLCELL_X2 FILLER_113_913 ();
 FILLCELL_X1 FILLER_113_915 ();
 FILLCELL_X1 FILLER_113_919 ();
 FILLCELL_X4 FILLER_113_944 ();
 FILLCELL_X1 FILLER_113_959 ();
 FILLCELL_X1 FILLER_113_973 ();
 FILLCELL_X1 FILLER_113_986 ();
 FILLCELL_X1 FILLER_113_998 ();
 FILLCELL_X1 FILLER_113_1012 ();
 FILLCELL_X8 FILLER_113_1019 ();
 FILLCELL_X4 FILLER_113_1027 ();
 FILLCELL_X32 FILLER_113_1055 ();
 FILLCELL_X16 FILLER_113_1087 ();
 FILLCELL_X8 FILLER_113_1103 ();
 FILLCELL_X4 FILLER_113_1111 ();
 FILLCELL_X2 FILLER_113_1115 ();
 FILLCELL_X1 FILLER_113_1117 ();
 FILLCELL_X4 FILLER_113_1138 ();
 FILLCELL_X8 FILLER_113_1159 ();
 FILLCELL_X4 FILLER_113_1167 ();
 FILLCELL_X2 FILLER_113_1171 ();
 FILLCELL_X1 FILLER_113_1239 ();
 FILLCELL_X2 FILLER_114_1 ();
 FILLCELL_X2 FILLER_114_27 ();
 FILLCELL_X1 FILLER_114_29 ();
 FILLCELL_X4 FILLER_114_37 ();
 FILLCELL_X1 FILLER_114_41 ();
 FILLCELL_X8 FILLER_114_63 ();
 FILLCELL_X8 FILLER_114_99 ();
 FILLCELL_X2 FILLER_114_107 ();
 FILLCELL_X1 FILLER_114_109 ();
 FILLCELL_X8 FILLER_114_117 ();
 FILLCELL_X1 FILLER_114_125 ();
 FILLCELL_X4 FILLER_114_140 ();
 FILLCELL_X2 FILLER_114_144 ();
 FILLCELL_X1 FILLER_114_146 ();
 FILLCELL_X2 FILLER_114_154 ();
 FILLCELL_X8 FILLER_114_180 ();
 FILLCELL_X8 FILLER_114_209 ();
 FILLCELL_X4 FILLER_114_217 ();
 FILLCELL_X2 FILLER_114_228 ();
 FILLCELL_X1 FILLER_114_230 ();
 FILLCELL_X8 FILLER_114_238 ();
 FILLCELL_X1 FILLER_114_246 ();
 FILLCELL_X16 FILLER_114_261 ();
 FILLCELL_X2 FILLER_114_277 ();
 FILLCELL_X1 FILLER_114_279 ();
 FILLCELL_X8 FILLER_114_291 ();
 FILLCELL_X1 FILLER_114_299 ();
 FILLCELL_X2 FILLER_114_314 ();
 FILLCELL_X8 FILLER_114_323 ();
 FILLCELL_X4 FILLER_114_331 ();
 FILLCELL_X1 FILLER_114_335 ();
 FILLCELL_X2 FILLER_114_343 ();
 FILLCELL_X4 FILLER_114_390 ();
 FILLCELL_X2 FILLER_114_394 ();
 FILLCELL_X1 FILLER_114_396 ();
 FILLCELL_X8 FILLER_114_404 ();
 FILLCELL_X4 FILLER_114_412 ();
 FILLCELL_X1 FILLER_114_416 ();
 FILLCELL_X4 FILLER_114_441 ();
 FILLCELL_X2 FILLER_114_445 ();
 FILLCELL_X1 FILLER_114_447 ();
 FILLCELL_X1 FILLER_114_477 ();
 FILLCELL_X4 FILLER_114_485 ();
 FILLCELL_X2 FILLER_114_489 ();
 FILLCELL_X16 FILLER_114_539 ();
 FILLCELL_X16 FILLER_114_586 ();
 FILLCELL_X2 FILLER_114_602 ();
 FILLCELL_X1 FILLER_114_604 ();
 FILLCELL_X8 FILLER_114_619 ();
 FILLCELL_X4 FILLER_114_627 ();
 FILLCELL_X8 FILLER_114_632 ();
 FILLCELL_X4 FILLER_114_640 ();
 FILLCELL_X4 FILLER_114_668 ();
 FILLCELL_X2 FILLER_114_672 ();
 FILLCELL_X1 FILLER_114_674 ();
 FILLCELL_X2 FILLER_114_689 ();
 FILLCELL_X8 FILLER_114_712 ();
 FILLCELL_X1 FILLER_114_720 ();
 FILLCELL_X8 FILLER_114_745 ();
 FILLCELL_X2 FILLER_114_753 ();
 FILLCELL_X1 FILLER_114_755 ();
 FILLCELL_X8 FILLER_114_775 ();
 FILLCELL_X8 FILLER_114_812 ();
 FILLCELL_X2 FILLER_114_820 ();
 FILLCELL_X1 FILLER_114_822 ();
 FILLCELL_X2 FILLER_114_836 ();
 FILLCELL_X1 FILLER_114_838 ();
 FILLCELL_X4 FILLER_114_846 ();
 FILLCELL_X2 FILLER_114_871 ();
 FILLCELL_X4 FILLER_114_877 ();
 FILLCELL_X2 FILLER_114_881 ();
 FILLCELL_X1 FILLER_114_883 ();
 FILLCELL_X1 FILLER_114_895 ();
 FILLCELL_X4 FILLER_114_905 ();
 FILLCELL_X4 FILLER_114_934 ();
 FILLCELL_X1 FILLER_114_938 ();
 FILLCELL_X1 FILLER_114_943 ();
 FILLCELL_X8 FILLER_114_962 ();
 FILLCELL_X2 FILLER_114_970 ();
 FILLCELL_X1 FILLER_114_999 ();
 FILLCELL_X4 FILLER_114_1011 ();
 FILLCELL_X8 FILLER_114_1019 ();
 FILLCELL_X2 FILLER_114_1027 ();
 FILLCELL_X2 FILLER_114_1033 ();
 FILLCELL_X32 FILLER_114_1043 ();
 FILLCELL_X16 FILLER_114_1075 ();
 FILLCELL_X8 FILLER_114_1091 ();
 FILLCELL_X4 FILLER_114_1099 ();
 FILLCELL_X1 FILLER_114_1103 ();
 FILLCELL_X1 FILLER_114_1135 ();
 FILLCELL_X4 FILLER_114_1143 ();
 FILLCELL_X1 FILLER_114_1147 ();
 FILLCELL_X2 FILLER_114_1155 ();
 FILLCELL_X1 FILLER_114_1157 ();
 FILLCELL_X2 FILLER_114_1170 ();
 FILLCELL_X2 FILLER_114_1179 ();
 FILLCELL_X1 FILLER_114_1181 ();
 FILLCELL_X1 FILLER_114_1199 ();
 FILLCELL_X1 FILLER_114_1234 ();
 FILLCELL_X1 FILLER_114_1239 ();
 FILLCELL_X16 FILLER_115_1 ();
 FILLCELL_X4 FILLER_115_17 ();
 FILLCELL_X8 FILLER_115_45 ();
 FILLCELL_X4 FILLER_115_53 ();
 FILLCELL_X2 FILLER_115_57 ();
 FILLCELL_X1 FILLER_115_59 ();
 FILLCELL_X4 FILLER_115_77 ();
 FILLCELL_X2 FILLER_115_81 ();
 FILLCELL_X8 FILLER_115_90 ();
 FILLCELL_X2 FILLER_115_98 ();
 FILLCELL_X2 FILLER_115_107 ();
 FILLCELL_X1 FILLER_115_109 ();
 FILLCELL_X4 FILLER_115_134 ();
 FILLCELL_X2 FILLER_115_138 ();
 FILLCELL_X8 FILLER_115_149 ();
 FILLCELL_X2 FILLER_115_157 ();
 FILLCELL_X8 FILLER_115_166 ();
 FILLCELL_X4 FILLER_115_174 ();
 FILLCELL_X1 FILLER_115_178 ();
 FILLCELL_X4 FILLER_115_186 ();
 FILLCELL_X1 FILLER_115_213 ();
 FILLCELL_X1 FILLER_115_231 ();
 FILLCELL_X2 FILLER_115_239 ();
 FILLCELL_X2 FILLER_115_248 ();
 FILLCELL_X1 FILLER_115_250 ();
 FILLCELL_X32 FILLER_115_275 ();
 FILLCELL_X16 FILLER_115_307 ();
 FILLCELL_X8 FILLER_115_323 ();
 FILLCELL_X2 FILLER_115_331 ();
 FILLCELL_X1 FILLER_115_333 ();
 FILLCELL_X4 FILLER_115_341 ();
 FILLCELL_X4 FILLER_115_352 ();
 FILLCELL_X32 FILLER_115_366 ();
 FILLCELL_X32 FILLER_115_398 ();
 FILLCELL_X4 FILLER_115_430 ();
 FILLCELL_X2 FILLER_115_434 ();
 FILLCELL_X8 FILLER_115_443 ();
 FILLCELL_X2 FILLER_115_451 ();
 FILLCELL_X1 FILLER_115_453 ();
 FILLCELL_X1 FILLER_115_461 ();
 FILLCELL_X2 FILLER_115_479 ();
 FILLCELL_X2 FILLER_115_486 ();
 FILLCELL_X2 FILLER_115_495 ();
 FILLCELL_X1 FILLER_115_497 ();
 FILLCELL_X8 FILLER_115_515 ();
 FILLCELL_X4 FILLER_115_523 ();
 FILLCELL_X2 FILLER_115_527 ();
 FILLCELL_X1 FILLER_115_529 ();
 FILLCELL_X8 FILLER_115_537 ();
 FILLCELL_X2 FILLER_115_545 ();
 FILLCELL_X1 FILLER_115_564 ();
 FILLCELL_X1 FILLER_115_572 ();
 FILLCELL_X1 FILLER_115_590 ();
 FILLCELL_X2 FILLER_115_598 ();
 FILLCELL_X1 FILLER_115_617 ();
 FILLCELL_X2 FILLER_115_625 ();
 FILLCELL_X1 FILLER_115_627 ();
 FILLCELL_X4 FILLER_115_641 ();
 FILLCELL_X1 FILLER_115_645 ();
 FILLCELL_X2 FILLER_115_663 ();
 FILLCELL_X2 FILLER_115_678 ();
 FILLCELL_X4 FILLER_115_711 ();
 FILLCELL_X1 FILLER_115_715 ();
 FILLCELL_X32 FILLER_115_718 ();
 FILLCELL_X4 FILLER_115_750 ();
 FILLCELL_X2 FILLER_115_754 ();
 FILLCELL_X4 FILLER_115_761 ();
 FILLCELL_X2 FILLER_115_765 ();
 FILLCELL_X1 FILLER_115_767 ();
 FILLCELL_X2 FILLER_115_775 ();
 FILLCELL_X4 FILLER_115_779 ();
 FILLCELL_X2 FILLER_115_783 ();
 FILLCELL_X1 FILLER_115_788 ();
 FILLCELL_X1 FILLER_115_795 ();
 FILLCELL_X4 FILLER_115_800 ();
 FILLCELL_X2 FILLER_115_806 ();
 FILLCELL_X1 FILLER_115_808 ();
 FILLCELL_X16 FILLER_115_811 ();
 FILLCELL_X4 FILLER_115_827 ();
 FILLCELL_X2 FILLER_115_831 ();
 FILLCELL_X1 FILLER_115_833 ();
 FILLCELL_X16 FILLER_115_870 ();
 FILLCELL_X1 FILLER_115_886 ();
 FILLCELL_X4 FILLER_115_892 ();
 FILLCELL_X1 FILLER_115_904 ();
 FILLCELL_X8 FILLER_115_937 ();
 FILLCELL_X4 FILLER_115_945 ();
 FILLCELL_X8 FILLER_115_952 ();
 FILLCELL_X4 FILLER_115_960 ();
 FILLCELL_X2 FILLER_115_964 ();
 FILLCELL_X2 FILLER_115_971 ();
 FILLCELL_X1 FILLER_115_973 ();
 FILLCELL_X2 FILLER_115_977 ();
 FILLCELL_X4 FILLER_115_993 ();
 FILLCELL_X1 FILLER_115_997 ();
 FILLCELL_X1 FILLER_115_1007 ();
 FILLCELL_X2 FILLER_115_1014 ();
 FILLCELL_X4 FILLER_115_1021 ();
 FILLCELL_X1 FILLER_115_1037 ();
 FILLCELL_X1 FILLER_115_1048 ();
 FILLCELL_X1 FILLER_115_1051 ();
 FILLCELL_X1 FILLER_115_1072 ();
 FILLCELL_X4 FILLER_115_1075 ();
 FILLCELL_X2 FILLER_115_1081 ();
 FILLCELL_X8 FILLER_115_1093 ();
 FILLCELL_X2 FILLER_115_1101 ();
 FILLCELL_X1 FILLER_115_1120 ();
 FILLCELL_X1 FILLER_115_1130 ();
 FILLCELL_X8 FILLER_115_1138 ();
 FILLCELL_X2 FILLER_115_1146 ();
 FILLCELL_X1 FILLER_115_1165 ();
 FILLCELL_X2 FILLER_115_1170 ();
 FILLCELL_X1 FILLER_115_1172 ();
 FILLCELL_X2 FILLER_115_1180 ();
 FILLCELL_X1 FILLER_115_1182 ();
 FILLCELL_X2 FILLER_115_1200 ();
 FILLCELL_X1 FILLER_116_1 ();
 FILLCELL_X8 FILLER_116_5 ();
 FILLCELL_X4 FILLER_116_13 ();
 FILLCELL_X16 FILLER_116_21 ();
 FILLCELL_X8 FILLER_116_37 ();
 FILLCELL_X4 FILLER_116_45 ();
 FILLCELL_X2 FILLER_116_49 ();
 FILLCELL_X1 FILLER_116_51 ();
 FILLCELL_X8 FILLER_116_63 ();
 FILLCELL_X1 FILLER_116_95 ();
 FILLCELL_X1 FILLER_116_113 ();
 FILLCELL_X1 FILLER_116_131 ();
 FILLCELL_X8 FILLER_116_139 ();
 FILLCELL_X2 FILLER_116_147 ();
 FILLCELL_X8 FILLER_116_184 ();
 FILLCELL_X4 FILLER_116_192 ();
 FILLCELL_X1 FILLER_116_196 ();
 FILLCELL_X2 FILLER_116_204 ();
 FILLCELL_X4 FILLER_116_223 ();
 FILLCELL_X1 FILLER_116_251 ();
 FILLCELL_X1 FILLER_116_259 ();
 FILLCELL_X1 FILLER_116_267 ();
 FILLCELL_X2 FILLER_116_275 ();
 FILLCELL_X16 FILLER_116_284 ();
 FILLCELL_X4 FILLER_116_300 ();
 FILLCELL_X16 FILLER_116_321 ();
 FILLCELL_X16 FILLER_116_354 ();
 FILLCELL_X8 FILLER_116_370 ();
 FILLCELL_X4 FILLER_116_378 ();
 FILLCELL_X2 FILLER_116_382 ();
 FILLCELL_X32 FILLER_116_401 ();
 FILLCELL_X8 FILLER_116_433 ();
 FILLCELL_X4 FILLER_116_441 ();
 FILLCELL_X2 FILLER_116_445 ();
 FILLCELL_X16 FILLER_116_452 ();
 FILLCELL_X1 FILLER_116_468 ();
 FILLCELL_X4 FILLER_116_493 ();
 FILLCELL_X2 FILLER_116_497 ();
 FILLCELL_X1 FILLER_116_499 ();
 FILLCELL_X4 FILLER_116_505 ();
 FILLCELL_X1 FILLER_116_513 ();
 FILLCELL_X8 FILLER_116_523 ();
 FILLCELL_X8 FILLER_116_548 ();
 FILLCELL_X4 FILLER_116_556 ();
 FILLCELL_X1 FILLER_116_560 ();
 FILLCELL_X8 FILLER_116_578 ();
 FILLCELL_X4 FILLER_116_586 ();
 FILLCELL_X1 FILLER_116_607 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X2 FILLER_116_632 ();
 FILLCELL_X1 FILLER_116_634 ();
 FILLCELL_X4 FILLER_116_670 ();
 FILLCELL_X32 FILLER_116_727 ();
 FILLCELL_X2 FILLER_116_759 ();
 FILLCELL_X1 FILLER_116_761 ();
 FILLCELL_X4 FILLER_116_787 ();
 FILLCELL_X2 FILLER_116_791 ();
 FILLCELL_X8 FILLER_116_795 ();
 FILLCELL_X1 FILLER_116_803 ();
 FILLCELL_X16 FILLER_116_807 ();
 FILLCELL_X8 FILLER_116_823 ();
 FILLCELL_X4 FILLER_116_831 ();
 FILLCELL_X1 FILLER_116_835 ();
 FILLCELL_X1 FILLER_116_842 ();
 FILLCELL_X1 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_864 ();
 FILLCELL_X2 FILLER_116_896 ();
 FILLCELL_X1 FILLER_116_901 ();
 FILLCELL_X1 FILLER_116_922 ();
 FILLCELL_X4 FILLER_116_942 ();
 FILLCELL_X1 FILLER_116_946 ();
 FILLCELL_X2 FILLER_116_966 ();
 FILLCELL_X4 FILLER_116_982 ();
 FILLCELL_X4 FILLER_116_1020 ();
 FILLCELL_X2 FILLER_116_1038 ();
 FILLCELL_X4 FILLER_116_1057 ();
 FILLCELL_X1 FILLER_116_1065 ();
 FILLCELL_X1 FILLER_116_1070 ();
 FILLCELL_X1 FILLER_116_1075 ();
 FILLCELL_X8 FILLER_116_1092 ();
 FILLCELL_X2 FILLER_116_1117 ();
 FILLCELL_X1 FILLER_116_1119 ();
 FILLCELL_X2 FILLER_116_1127 ();
 FILLCELL_X1 FILLER_116_1153 ();
 FILLCELL_X1 FILLER_116_1167 ();
 FILLCELL_X1 FILLER_116_1175 ();
 FILLCELL_X16 FILLER_117_1 ();
 FILLCELL_X2 FILLER_117_17 ();
 FILLCELL_X1 FILLER_117_19 ();
 FILLCELL_X32 FILLER_117_25 ();
 FILLCELL_X1 FILLER_117_57 ();
 FILLCELL_X16 FILLER_117_75 ();
 FILLCELL_X8 FILLER_117_91 ();
 FILLCELL_X4 FILLER_117_99 ();
 FILLCELL_X2 FILLER_117_103 ();
 FILLCELL_X1 FILLER_117_105 ();
 FILLCELL_X16 FILLER_117_137 ();
 FILLCELL_X8 FILLER_117_153 ();
 FILLCELL_X1 FILLER_117_161 ();
 FILLCELL_X4 FILLER_117_203 ();
 FILLCELL_X1 FILLER_117_207 ();
 FILLCELL_X16 FILLER_117_225 ();
 FILLCELL_X4 FILLER_117_241 ();
 FILLCELL_X16 FILLER_117_252 ();
 FILLCELL_X2 FILLER_117_268 ();
 FILLCELL_X8 FILLER_117_287 ();
 FILLCELL_X4 FILLER_117_295 ();
 FILLCELL_X2 FILLER_117_299 ();
 FILLCELL_X1 FILLER_117_301 ();
 FILLCELL_X4 FILLER_117_317 ();
 FILLCELL_X2 FILLER_117_321 ();
 FILLCELL_X1 FILLER_117_323 ();
 FILLCELL_X1 FILLER_117_338 ();
 FILLCELL_X16 FILLER_117_346 ();
 FILLCELL_X1 FILLER_117_362 ();
 FILLCELL_X2 FILLER_117_408 ();
 FILLCELL_X1 FILLER_117_410 ();
 FILLCELL_X1 FILLER_117_445 ();
 FILLCELL_X1 FILLER_117_456 ();
 FILLCELL_X1 FILLER_117_464 ();
 FILLCELL_X2 FILLER_117_472 ();
 FILLCELL_X1 FILLER_117_487 ();
 FILLCELL_X2 FILLER_117_505 ();
 FILLCELL_X32 FILLER_117_527 ();
 FILLCELL_X8 FILLER_117_559 ();
 FILLCELL_X16 FILLER_117_574 ();
 FILLCELL_X2 FILLER_117_590 ();
 FILLCELL_X1 FILLER_117_592 ();
 FILLCELL_X8 FILLER_117_624 ();
 FILLCELL_X4 FILLER_117_632 ();
 FILLCELL_X2 FILLER_117_636 ();
 FILLCELL_X1 FILLER_117_662 ();
 FILLCELL_X1 FILLER_117_687 ();
 FILLCELL_X1 FILLER_117_695 ();
 FILLCELL_X8 FILLER_117_703 ();
 FILLCELL_X4 FILLER_117_711 ();
 FILLCELL_X1 FILLER_117_715 ();
 FILLCELL_X1 FILLER_117_744 ();
 FILLCELL_X1 FILLER_117_798 ();
 FILLCELL_X4 FILLER_117_826 ();
 FILLCELL_X1 FILLER_117_830 ();
 FILLCELL_X4 FILLER_117_834 ();
 FILLCELL_X1 FILLER_117_838 ();
 FILLCELL_X2 FILLER_117_851 ();
 FILLCELL_X2 FILLER_117_869 ();
 FILLCELL_X4 FILLER_117_880 ();
 FILLCELL_X1 FILLER_117_884 ();
 FILLCELL_X1 FILLER_117_889 ();
 FILLCELL_X2 FILLER_117_900 ();
 FILLCELL_X8 FILLER_117_907 ();
 FILLCELL_X2 FILLER_117_919 ();
 FILLCELL_X2 FILLER_117_928 ();
 FILLCELL_X8 FILLER_117_934 ();
 FILLCELL_X1 FILLER_117_942 ();
 FILLCELL_X4 FILLER_117_974 ();
 FILLCELL_X2 FILLER_117_978 ();
 FILLCELL_X1 FILLER_117_980 ();
 FILLCELL_X8 FILLER_117_990 ();
 FILLCELL_X2 FILLER_117_1021 ();
 FILLCELL_X1 FILLER_117_1023 ();
 FILLCELL_X16 FILLER_117_1031 ();
 FILLCELL_X1 FILLER_117_1062 ();
 FILLCELL_X1 FILLER_117_1066 ();
 FILLCELL_X2 FILLER_117_1076 ();
 FILLCELL_X16 FILLER_117_1097 ();
 FILLCELL_X1 FILLER_117_1113 ();
 FILLCELL_X32 FILLER_117_1121 ();
 FILLCELL_X16 FILLER_117_1153 ();
 FILLCELL_X2 FILLER_117_1169 ();
 FILLCELL_X1 FILLER_117_1171 ();
 FILLCELL_X4 FILLER_117_1189 ();
 FILLCELL_X1 FILLER_117_1193 ();
 FILLCELL_X4 FILLER_118_1 ();
 FILLCELL_X2 FILLER_118_29 ();
 FILLCELL_X4 FILLER_118_72 ();
 FILLCELL_X1 FILLER_118_76 ();
 FILLCELL_X32 FILLER_118_84 ();
 FILLCELL_X32 FILLER_118_116 ();
 FILLCELL_X32 FILLER_118_148 ();
 FILLCELL_X16 FILLER_118_180 ();
 FILLCELL_X8 FILLER_118_196 ();
 FILLCELL_X8 FILLER_118_211 ();
 FILLCELL_X4 FILLER_118_219 ();
 FILLCELL_X2 FILLER_118_223 ();
 FILLCELL_X1 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_233 ();
 FILLCELL_X4 FILLER_118_265 ();
 FILLCELL_X2 FILLER_118_324 ();
 FILLCELL_X8 FILLER_118_357 ();
 FILLCELL_X4 FILLER_118_365 ();
 FILLCELL_X2 FILLER_118_369 ();
 FILLCELL_X1 FILLER_118_371 ();
 FILLCELL_X16 FILLER_118_403 ();
 FILLCELL_X1 FILLER_118_419 ();
 FILLCELL_X8 FILLER_118_444 ();
 FILLCELL_X1 FILLER_118_452 ();
 FILLCELL_X16 FILLER_118_470 ();
 FILLCELL_X1 FILLER_118_486 ();
 FILLCELL_X8 FILLER_118_494 ();
 FILLCELL_X2 FILLER_118_502 ();
 FILLCELL_X2 FILLER_118_518 ();
 FILLCELL_X1 FILLER_118_527 ();
 FILLCELL_X16 FILLER_118_545 ();
 FILLCELL_X8 FILLER_118_561 ();
 FILLCELL_X4 FILLER_118_569 ();
 FILLCELL_X1 FILLER_118_573 ();
 FILLCELL_X16 FILLER_118_579 ();
 FILLCELL_X8 FILLER_118_595 ();
 FILLCELL_X4 FILLER_118_603 ();
 FILLCELL_X2 FILLER_118_607 ();
 FILLCELL_X8 FILLER_118_614 ();
 FILLCELL_X4 FILLER_118_627 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X16 FILLER_118_696 ();
 FILLCELL_X4 FILLER_118_712 ();
 FILLCELL_X1 FILLER_118_716 ();
 FILLCELL_X4 FILLER_118_719 ();
 FILLCELL_X1 FILLER_118_723 ();
 FILLCELL_X8 FILLER_118_740 ();
 FILLCELL_X4 FILLER_118_748 ();
 FILLCELL_X2 FILLER_118_752 ();
 FILLCELL_X1 FILLER_118_754 ();
 FILLCELL_X2 FILLER_118_783 ();
 FILLCELL_X1 FILLER_118_828 ();
 FILLCELL_X2 FILLER_118_846 ();
 FILLCELL_X1 FILLER_118_848 ();
 FILLCELL_X1 FILLER_118_856 ();
 FILLCELL_X1 FILLER_118_870 ();
 FILLCELL_X1 FILLER_118_874 ();
 FILLCELL_X4 FILLER_118_879 ();
 FILLCELL_X16 FILLER_118_890 ();
 FILLCELL_X4 FILLER_118_906 ();
 FILLCELL_X2 FILLER_118_910 ();
 FILLCELL_X4 FILLER_118_923 ();
 FILLCELL_X2 FILLER_118_931 ();
 FILLCELL_X1 FILLER_118_933 ();
 FILLCELL_X2 FILLER_118_937 ();
 FILLCELL_X1 FILLER_118_939 ();
 FILLCELL_X8 FILLER_118_978 ();
 FILLCELL_X1 FILLER_118_986 ();
 FILLCELL_X2 FILLER_118_1018 ();
 FILLCELL_X8 FILLER_118_1024 ();
 FILLCELL_X16 FILLER_118_1037 ();
 FILLCELL_X4 FILLER_118_1053 ();
 FILLCELL_X2 FILLER_118_1057 ();
 FILLCELL_X32 FILLER_118_1092 ();
 FILLCELL_X1 FILLER_118_1124 ();
 FILLCELL_X8 FILLER_118_1142 ();
 FILLCELL_X4 FILLER_118_1150 ();
 FILLCELL_X2 FILLER_118_1154 ();
 FILLCELL_X1 FILLER_118_1188 ();
 FILLCELL_X2 FILLER_118_1238 ();
 FILLCELL_X4 FILLER_119_1 ();
 FILLCELL_X2 FILLER_119_39 ();
 FILLCELL_X1 FILLER_119_41 ();
 FILLCELL_X8 FILLER_119_49 ();
 FILLCELL_X2 FILLER_119_57 ();
 FILLCELL_X2 FILLER_119_90 ();
 FILLCELL_X1 FILLER_119_92 ();
 FILLCELL_X4 FILLER_119_110 ();
 FILLCELL_X1 FILLER_119_114 ();
 FILLCELL_X2 FILLER_119_132 ();
 FILLCELL_X1 FILLER_119_134 ();
 FILLCELL_X4 FILLER_119_142 ();
 FILLCELL_X2 FILLER_119_146 ();
 FILLCELL_X1 FILLER_119_148 ();
 FILLCELL_X16 FILLER_119_173 ();
 FILLCELL_X4 FILLER_119_189 ();
 FILLCELL_X2 FILLER_119_193 ();
 FILLCELL_X16 FILLER_119_216 ();
 FILLCELL_X1 FILLER_119_232 ();
 FILLCELL_X4 FILLER_119_250 ();
 FILLCELL_X8 FILLER_119_261 ();
 FILLCELL_X4 FILLER_119_331 ();
 FILLCELL_X4 FILLER_119_365 ();
 FILLCELL_X2 FILLER_119_369 ();
 FILLCELL_X1 FILLER_119_371 ();
 FILLCELL_X8 FILLER_119_396 ();
 FILLCELL_X2 FILLER_119_404 ();
 FILLCELL_X1 FILLER_119_451 ();
 FILLCELL_X1 FILLER_119_466 ();
 FILLCELL_X8 FILLER_119_498 ();
 FILLCELL_X2 FILLER_119_506 ();
 FILLCELL_X1 FILLER_119_508 ();
 FILLCELL_X1 FILLER_119_516 ();
 FILLCELL_X8 FILLER_119_541 ();
 FILLCELL_X4 FILLER_119_549 ();
 FILLCELL_X4 FILLER_119_560 ();
 FILLCELL_X2 FILLER_119_564 ();
 FILLCELL_X2 FILLER_119_573 ();
 FILLCELL_X8 FILLER_119_599 ();
 FILLCELL_X1 FILLER_119_607 ();
 FILLCELL_X4 FILLER_119_622 ();
 FILLCELL_X8 FILLER_119_639 ();
 FILLCELL_X32 FILLER_119_659 ();
 FILLCELL_X16 FILLER_119_699 ();
 FILLCELL_X8 FILLER_119_715 ();
 FILLCELL_X4 FILLER_119_723 ();
 FILLCELL_X2 FILLER_119_727 ();
 FILLCELL_X1 FILLER_119_729 ();
 FILLCELL_X2 FILLER_119_781 ();
 FILLCELL_X2 FILLER_119_809 ();
 FILLCELL_X1 FILLER_119_811 ();
 FILLCELL_X4 FILLER_119_815 ();
 FILLCELL_X2 FILLER_119_822 ();
 FILLCELL_X8 FILLER_119_827 ();
 FILLCELL_X2 FILLER_119_845 ();
 FILLCELL_X1 FILLER_119_847 ();
 FILLCELL_X1 FILLER_119_864 ();
 FILLCELL_X16 FILLER_119_868 ();
 FILLCELL_X4 FILLER_119_889 ();
 FILLCELL_X16 FILLER_119_897 ();
 FILLCELL_X4 FILLER_119_933 ();
 FILLCELL_X2 FILLER_119_937 ();
 FILLCELL_X2 FILLER_119_944 ();
 FILLCELL_X1 FILLER_119_957 ();
 FILLCELL_X1 FILLER_119_969 ();
 FILLCELL_X2 FILLER_119_972 ();
 FILLCELL_X2 FILLER_119_985 ();
 FILLCELL_X4 FILLER_119_1007 ();
 FILLCELL_X2 FILLER_119_1018 ();
 FILLCELL_X1 FILLER_119_1033 ();
 FILLCELL_X16 FILLER_119_1038 ();
 FILLCELL_X4 FILLER_119_1054 ();
 FILLCELL_X2 FILLER_119_1058 ();
 FILLCELL_X4 FILLER_119_1064 ();
 FILLCELL_X2 FILLER_119_1068 ();
 FILLCELL_X1 FILLER_119_1070 ();
 FILLCELL_X32 FILLER_119_1074 ();
 FILLCELL_X1 FILLER_119_1106 ();
 FILLCELL_X2 FILLER_119_1143 ();
 FILLCELL_X1 FILLER_120_4 ();
 FILLCELL_X4 FILLER_120_19 ();
 FILLCELL_X2 FILLER_120_23 ();
 FILLCELL_X2 FILLER_120_46 ();
 FILLCELL_X8 FILLER_120_52 ();
 FILLCELL_X2 FILLER_120_60 ();
 FILLCELL_X8 FILLER_120_67 ();
 FILLCELL_X2 FILLER_120_75 ();
 FILLCELL_X1 FILLER_120_77 ();
 FILLCELL_X4 FILLER_120_99 ();
 FILLCELL_X2 FILLER_120_103 ();
 FILLCELL_X2 FILLER_120_136 ();
 FILLCELL_X2 FILLER_120_147 ();
 FILLCELL_X8 FILLER_120_163 ();
 FILLCELL_X2 FILLER_120_171 ();
 FILLCELL_X2 FILLER_120_198 ();
 FILLCELL_X4 FILLER_120_224 ();
 FILLCELL_X2 FILLER_120_228 ();
 FILLCELL_X16 FILLER_120_261 ();
 FILLCELL_X4 FILLER_120_277 ();
 FILLCELL_X1 FILLER_120_288 ();
 FILLCELL_X16 FILLER_120_317 ();
 FILLCELL_X2 FILLER_120_340 ();
 FILLCELL_X32 FILLER_120_366 ();
 FILLCELL_X32 FILLER_120_398 ();
 FILLCELL_X8 FILLER_120_430 ();
 FILLCELL_X4 FILLER_120_438 ();
 FILLCELL_X2 FILLER_120_459 ();
 FILLCELL_X16 FILLER_120_478 ();
 FILLCELL_X8 FILLER_120_494 ();
 FILLCELL_X2 FILLER_120_502 ();
 FILLCELL_X1 FILLER_120_504 ();
 FILLCELL_X16 FILLER_120_520 ();
 FILLCELL_X8 FILLER_120_536 ();
 FILLCELL_X2 FILLER_120_544 ();
 FILLCELL_X1 FILLER_120_546 ();
 FILLCELL_X2 FILLER_120_597 ();
 FILLCELL_X1 FILLER_120_599 ();
 FILLCELL_X4 FILLER_120_624 ();
 FILLCELL_X2 FILLER_120_628 ();
 FILLCELL_X1 FILLER_120_630 ();
 FILLCELL_X2 FILLER_120_632 ();
 FILLCELL_X8 FILLER_120_667 ();
 FILLCELL_X2 FILLER_120_675 ();
 FILLCELL_X1 FILLER_120_677 ();
 FILLCELL_X4 FILLER_120_709 ();
 FILLCELL_X1 FILLER_120_713 ();
 FILLCELL_X2 FILLER_120_751 ();
 FILLCELL_X1 FILLER_120_753 ();
 FILLCELL_X4 FILLER_120_777 ();
 FILLCELL_X2 FILLER_120_781 ();
 FILLCELL_X1 FILLER_120_783 ();
 FILLCELL_X1 FILLER_120_789 ();
 FILLCELL_X4 FILLER_120_793 ();
 FILLCELL_X4 FILLER_120_799 ();
 FILLCELL_X2 FILLER_120_803 ();
 FILLCELL_X4 FILLER_120_808 ();
 FILLCELL_X1 FILLER_120_812 ();
 FILLCELL_X16 FILLER_120_819 ();
 FILLCELL_X8 FILLER_120_835 ();
 FILLCELL_X4 FILLER_120_843 ();
 FILLCELL_X4 FILLER_120_852 ();
 FILLCELL_X4 FILLER_120_888 ();
 FILLCELL_X2 FILLER_120_892 ();
 FILLCELL_X1 FILLER_120_894 ();
 FILLCELL_X4 FILLER_120_906 ();
 FILLCELL_X8 FILLER_120_949 ();
 FILLCELL_X4 FILLER_120_957 ();
 FILLCELL_X1 FILLER_120_961 ();
 FILLCELL_X1 FILLER_120_972 ();
 FILLCELL_X1 FILLER_120_984 ();
 FILLCELL_X2 FILLER_120_994 ();
 FILLCELL_X4 FILLER_120_1011 ();
 FILLCELL_X2 FILLER_120_1015 ();
 FILLCELL_X1 FILLER_120_1017 ();
 FILLCELL_X32 FILLER_120_1022 ();
 FILLCELL_X1 FILLER_120_1054 ();
 FILLCELL_X1 FILLER_120_1068 ();
 FILLCELL_X2 FILLER_120_1076 ();
 FILLCELL_X32 FILLER_120_1083 ();
 FILLCELL_X4 FILLER_120_1115 ();
 FILLCELL_X1 FILLER_120_1119 ();
 FILLCELL_X1 FILLER_120_1150 ();
 FILLCELL_X2 FILLER_120_1158 ();
 FILLCELL_X2 FILLER_120_1169 ();
 FILLCELL_X2 FILLER_120_1178 ();
 FILLCELL_X4 FILLER_120_1197 ();
 FILLCELL_X1 FILLER_120_1201 ();
 FILLCELL_X2 FILLER_120_1216 ();
 FILLCELL_X2 FILLER_120_1238 ();
 FILLCELL_X4 FILLER_121_1 ();
 FILLCELL_X1 FILLER_121_5 ();
 FILLCELL_X2 FILLER_121_23 ();
 FILLCELL_X1 FILLER_121_25 ();
 FILLCELL_X1 FILLER_121_33 ();
 FILLCELL_X1 FILLER_121_41 ();
 FILLCELL_X1 FILLER_121_49 ();
 FILLCELL_X2 FILLER_121_67 ();
 FILLCELL_X8 FILLER_121_76 ();
 FILLCELL_X8 FILLER_121_108 ();
 FILLCELL_X4 FILLER_121_116 ();
 FILLCELL_X1 FILLER_121_120 ();
 FILLCELL_X1 FILLER_121_135 ();
 FILLCELL_X16 FILLER_121_143 ();
 FILLCELL_X8 FILLER_121_159 ();
 FILLCELL_X4 FILLER_121_167 ();
 FILLCELL_X1 FILLER_121_171 ();
 FILLCELL_X8 FILLER_121_189 ();
 FILLCELL_X4 FILLER_121_197 ();
 FILLCELL_X4 FILLER_121_262 ();
 FILLCELL_X1 FILLER_121_266 ();
 FILLCELL_X1 FILLER_121_291 ();
 FILLCELL_X2 FILLER_121_309 ();
 FILLCELL_X1 FILLER_121_311 ();
 FILLCELL_X32 FILLER_121_336 ();
 FILLCELL_X8 FILLER_121_368 ();
 FILLCELL_X4 FILLER_121_376 ();
 FILLCELL_X2 FILLER_121_380 ();
 FILLCELL_X1 FILLER_121_382 ();
 FILLCELL_X32 FILLER_121_390 ();
 FILLCELL_X8 FILLER_121_422 ();
 FILLCELL_X4 FILLER_121_430 ();
 FILLCELL_X2 FILLER_121_441 ();
 FILLCELL_X1 FILLER_121_443 ();
 FILLCELL_X4 FILLER_121_451 ();
 FILLCELL_X1 FILLER_121_455 ();
 FILLCELL_X8 FILLER_121_463 ();
 FILLCELL_X4 FILLER_121_471 ();
 FILLCELL_X2 FILLER_121_482 ();
 FILLCELL_X4 FILLER_121_491 ();
 FILLCELL_X1 FILLER_121_495 ();
 FILLCELL_X1 FILLER_121_503 ();
 FILLCELL_X16 FILLER_121_511 ();
 FILLCELL_X4 FILLER_121_527 ();
 FILLCELL_X1 FILLER_121_531 ();
 FILLCELL_X8 FILLER_121_537 ();
 FILLCELL_X1 FILLER_121_545 ();
 FILLCELL_X2 FILLER_121_563 ();
 FILLCELL_X2 FILLER_121_572 ();
 FILLCELL_X4 FILLER_121_581 ();
 FILLCELL_X2 FILLER_121_602 ();
 FILLCELL_X1 FILLER_121_621 ();
 FILLCELL_X2 FILLER_121_639 ();
 FILLCELL_X2 FILLER_121_648 ();
 FILLCELL_X2 FILLER_121_667 ();
 FILLCELL_X1 FILLER_121_669 ();
 FILLCELL_X16 FILLER_121_713 ();
 FILLCELL_X8 FILLER_121_729 ();
 FILLCELL_X4 FILLER_121_737 ();
 FILLCELL_X1 FILLER_121_741 ();
 FILLCELL_X16 FILLER_121_756 ();
 FILLCELL_X2 FILLER_121_772 ();
 FILLCELL_X1 FILLER_121_774 ();
 FILLCELL_X16 FILLER_121_779 ();
 FILLCELL_X8 FILLER_121_795 ();
 FILLCELL_X1 FILLER_121_803 ();
 FILLCELL_X4 FILLER_121_809 ();
 FILLCELL_X2 FILLER_121_813 ();
 FILLCELL_X1 FILLER_121_824 ();
 FILLCELL_X4 FILLER_121_828 ();
 FILLCELL_X4 FILLER_121_841 ();
 FILLCELL_X2 FILLER_121_845 ();
 FILLCELL_X1 FILLER_121_854 ();
 FILLCELL_X4 FILLER_121_859 ();
 FILLCELL_X2 FILLER_121_863 ();
 FILLCELL_X2 FILLER_121_880 ();
 FILLCELL_X4 FILLER_121_887 ();
 FILLCELL_X1 FILLER_121_891 ();
 FILLCELL_X4 FILLER_121_906 ();
 FILLCELL_X1 FILLER_121_910 ();
 FILLCELL_X8 FILLER_121_933 ();
 FILLCELL_X2 FILLER_121_941 ();
 FILLCELL_X2 FILLER_121_949 ();
 FILLCELL_X1 FILLER_121_951 ();
 FILLCELL_X2 FILLER_121_959 ();
 FILLCELL_X1 FILLER_121_961 ();
 FILLCELL_X4 FILLER_121_965 ();
 FILLCELL_X2 FILLER_121_969 ();
 FILLCELL_X1 FILLER_121_971 ();
 FILLCELL_X8 FILLER_121_974 ();
 FILLCELL_X4 FILLER_121_982 ();
 FILLCELL_X1 FILLER_121_986 ();
 FILLCELL_X1 FILLER_121_1001 ();
 FILLCELL_X4 FILLER_121_1008 ();
 FILLCELL_X4 FILLER_121_1028 ();
 FILLCELL_X2 FILLER_121_1039 ();
 FILLCELL_X2 FILLER_121_1046 ();
 FILLCELL_X1 FILLER_121_1065 ();
 FILLCELL_X2 FILLER_121_1074 ();
 FILLCELL_X1 FILLER_121_1079 ();
 FILLCELL_X8 FILLER_121_1083 ();
 FILLCELL_X4 FILLER_121_1091 ();
 FILLCELL_X2 FILLER_121_1095 ();
 FILLCELL_X1 FILLER_121_1097 ();
 FILLCELL_X16 FILLER_121_1109 ();
 FILLCELL_X2 FILLER_121_1125 ();
 FILLCELL_X1 FILLER_121_1127 ();
 FILLCELL_X2 FILLER_121_1152 ();
 FILLCELL_X1 FILLER_121_1154 ();
 FILLCELL_X2 FILLER_121_1179 ();
 FILLCELL_X2 FILLER_121_1188 ();
 FILLCELL_X2 FILLER_121_1207 ();
 FILLCELL_X2 FILLER_121_1226 ();
 FILLCELL_X16 FILLER_122_1 ();
 FILLCELL_X1 FILLER_122_17 ();
 FILLCELL_X4 FILLER_122_42 ();
 FILLCELL_X2 FILLER_122_46 ();
 FILLCELL_X1 FILLER_122_48 ();
 FILLCELL_X32 FILLER_122_73 ();
 FILLCELL_X32 FILLER_122_105 ();
 FILLCELL_X16 FILLER_122_137 ();
 FILLCELL_X8 FILLER_122_153 ();
 FILLCELL_X4 FILLER_122_161 ();
 FILLCELL_X2 FILLER_122_165 ();
 FILLCELL_X2 FILLER_122_181 ();
 FILLCELL_X1 FILLER_122_183 ();
 FILLCELL_X4 FILLER_122_208 ();
 FILLCELL_X1 FILLER_122_212 ();
 FILLCELL_X4 FILLER_122_220 ();
 FILLCELL_X4 FILLER_122_231 ();
 FILLCELL_X2 FILLER_122_235 ();
 FILLCELL_X32 FILLER_122_240 ();
 FILLCELL_X16 FILLER_122_272 ();
 FILLCELL_X4 FILLER_122_288 ();
 FILLCELL_X1 FILLER_122_292 ();
 FILLCELL_X8 FILLER_122_300 ();
 FILLCELL_X4 FILLER_122_308 ();
 FILLCELL_X16 FILLER_122_319 ();
 FILLCELL_X4 FILLER_122_335 ();
 FILLCELL_X8 FILLER_122_346 ();
 FILLCELL_X2 FILLER_122_354 ();
 FILLCELL_X1 FILLER_122_356 ();
 FILLCELL_X1 FILLER_122_365 ();
 FILLCELL_X32 FILLER_122_400 ();
 FILLCELL_X1 FILLER_122_432 ();
 FILLCELL_X2 FILLER_122_450 ();
 FILLCELL_X1 FILLER_122_452 ();
 FILLCELL_X1 FILLER_122_474 ();
 FILLCELL_X4 FILLER_122_492 ();
 FILLCELL_X2 FILLER_122_496 ();
 FILLCELL_X32 FILLER_122_522 ();
 FILLCELL_X8 FILLER_122_554 ();
 FILLCELL_X16 FILLER_122_569 ();
 FILLCELL_X4 FILLER_122_585 ();
 FILLCELL_X8 FILLER_122_620 ();
 FILLCELL_X2 FILLER_122_628 ();
 FILLCELL_X1 FILLER_122_630 ();
 FILLCELL_X2 FILLER_122_632 ();
 FILLCELL_X2 FILLER_122_641 ();
 FILLCELL_X1 FILLER_122_643 ();
 FILLCELL_X4 FILLER_122_696 ();
 FILLCELL_X2 FILLER_122_700 ();
 FILLCELL_X1 FILLER_122_702 ();
 FILLCELL_X2 FILLER_122_707 ();
 FILLCELL_X2 FILLER_122_721 ();
 FILLCELL_X16 FILLER_122_736 ();
 FILLCELL_X4 FILLER_122_752 ();
 FILLCELL_X2 FILLER_122_756 ();
 FILLCELL_X1 FILLER_122_758 ();
 FILLCELL_X4 FILLER_122_793 ();
 FILLCELL_X2 FILLER_122_797 ();
 FILLCELL_X1 FILLER_122_833 ();
 FILLCELL_X16 FILLER_122_854 ();
 FILLCELL_X4 FILLER_122_870 ();
 FILLCELL_X1 FILLER_122_874 ();
 FILLCELL_X2 FILLER_122_882 ();
 FILLCELL_X2 FILLER_122_887 ();
 FILLCELL_X1 FILLER_122_889 ();
 FILLCELL_X4 FILLER_122_900 ();
 FILLCELL_X2 FILLER_122_916 ();
 FILLCELL_X4 FILLER_122_922 ();
 FILLCELL_X1 FILLER_122_926 ();
 FILLCELL_X1 FILLER_122_930 ();
 FILLCELL_X1 FILLER_122_938 ();
 FILLCELL_X2 FILLER_122_953 ();
 FILLCELL_X4 FILLER_122_970 ();
 FILLCELL_X2 FILLER_122_987 ();
 FILLCELL_X16 FILLER_122_1004 ();
 FILLCELL_X4 FILLER_122_1020 ();
 FILLCELL_X4 FILLER_122_1037 ();
 FILLCELL_X1 FILLER_122_1046 ();
 FILLCELL_X1 FILLER_122_1053 ();
 FILLCELL_X1 FILLER_122_1060 ();
 FILLCELL_X2 FILLER_122_1067 ();
 FILLCELL_X4 FILLER_122_1076 ();
 FILLCELL_X1 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1084 ();
 FILLCELL_X8 FILLER_122_1116 ();
 FILLCELL_X4 FILLER_122_1124 ();
 FILLCELL_X2 FILLER_122_1128 ();
 FILLCELL_X4 FILLER_122_1147 ();
 FILLCELL_X2 FILLER_122_1151 ();
 FILLCELL_X1 FILLER_122_1153 ();
 FILLCELL_X8 FILLER_122_1170 ();
 FILLCELL_X4 FILLER_122_1178 ();
 FILLCELL_X2 FILLER_122_1182 ();
 FILLCELL_X1 FILLER_122_1224 ();
 FILLCELL_X4 FILLER_122_1236 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X16 FILLER_123_33 ();
 FILLCELL_X4 FILLER_123_49 ();
 FILLCELL_X32 FILLER_123_60 ();
 FILLCELL_X8 FILLER_123_92 ();
 FILLCELL_X4 FILLER_123_100 ();
 FILLCELL_X2 FILLER_123_104 ();
 FILLCELL_X1 FILLER_123_106 ();
 FILLCELL_X8 FILLER_123_124 ();
 FILLCELL_X4 FILLER_123_132 ();
 FILLCELL_X2 FILLER_123_136 ();
 FILLCELL_X32 FILLER_123_143 ();
 FILLCELL_X2 FILLER_123_175 ();
 FILLCELL_X16 FILLER_123_184 ();
 FILLCELL_X8 FILLER_123_200 ();
 FILLCELL_X4 FILLER_123_208 ();
 FILLCELL_X2 FILLER_123_212 ();
 FILLCELL_X16 FILLER_123_221 ();
 FILLCELL_X2 FILLER_123_237 ();
 FILLCELL_X1 FILLER_123_239 ();
 FILLCELL_X32 FILLER_123_247 ();
 FILLCELL_X32 FILLER_123_279 ();
 FILLCELL_X1 FILLER_123_311 ();
 FILLCELL_X2 FILLER_123_329 ();
 FILLCELL_X8 FILLER_123_355 ();
 FILLCELL_X2 FILLER_123_363 ();
 FILLCELL_X1 FILLER_123_365 ();
 FILLCELL_X4 FILLER_123_407 ();
 FILLCELL_X32 FILLER_123_432 ();
 FILLCELL_X16 FILLER_123_464 ();
 FILLCELL_X4 FILLER_123_480 ();
 FILLCELL_X2 FILLER_123_484 ();
 FILLCELL_X1 FILLER_123_486 ();
 FILLCELL_X32 FILLER_123_521 ();
 FILLCELL_X32 FILLER_123_553 ();
 FILLCELL_X32 FILLER_123_585 ();
 FILLCELL_X16 FILLER_123_617 ();
 FILLCELL_X8 FILLER_123_633 ();
 FILLCELL_X4 FILLER_123_641 ();
 FILLCELL_X2 FILLER_123_645 ();
 FILLCELL_X1 FILLER_123_647 ();
 FILLCELL_X1 FILLER_123_655 ();
 FILLCELL_X16 FILLER_123_670 ();
 FILLCELL_X1 FILLER_123_699 ();
 FILLCELL_X4 FILLER_123_713 ();
 FILLCELL_X4 FILLER_123_749 ();
 FILLCELL_X2 FILLER_123_753 ();
 FILLCELL_X1 FILLER_123_762 ();
 FILLCELL_X2 FILLER_123_771 ();
 FILLCELL_X1 FILLER_123_773 ();
 FILLCELL_X8 FILLER_123_781 ();
 FILLCELL_X2 FILLER_123_789 ();
 FILLCELL_X1 FILLER_123_791 ();
 FILLCELL_X1 FILLER_123_831 ();
 FILLCELL_X32 FILLER_123_846 ();
 FILLCELL_X8 FILLER_123_878 ();
 FILLCELL_X4 FILLER_123_886 ();
 FILLCELL_X1 FILLER_123_890 ();
 FILLCELL_X4 FILLER_123_904 ();
 FILLCELL_X2 FILLER_123_908 ();
 FILLCELL_X1 FILLER_123_910 ();
 FILLCELL_X1 FILLER_123_918 ();
 FILLCELL_X4 FILLER_123_943 ();
 FILLCELL_X1 FILLER_123_947 ();
 FILLCELL_X1 FILLER_123_959 ();
 FILLCELL_X8 FILLER_123_967 ();
 FILLCELL_X1 FILLER_123_993 ();
 FILLCELL_X8 FILLER_123_1005 ();
 FILLCELL_X1 FILLER_123_1013 ();
 FILLCELL_X1 FILLER_123_1068 ();
 FILLCELL_X4 FILLER_123_1083 ();
 FILLCELL_X2 FILLER_123_1087 ();
 FILLCELL_X1 FILLER_123_1089 ();
 FILLCELL_X32 FILLER_123_1092 ();
 FILLCELL_X16 FILLER_123_1124 ();
 FILLCELL_X2 FILLER_123_1140 ();
 FILLCELL_X1 FILLER_123_1142 ();
 FILLCELL_X2 FILLER_123_1167 ();
 FILLCELL_X1 FILLER_123_1169 ();
 FILLCELL_X4 FILLER_123_1177 ();
 FILLCELL_X2 FILLER_123_1181 ();
 FILLCELL_X8 FILLER_123_1190 ();
 FILLCELL_X1 FILLER_123_1198 ();
 FILLCELL_X8 FILLER_123_1206 ();
 FILLCELL_X4 FILLER_123_1214 ();
 FILLCELL_X2 FILLER_123_1228 ();
 FILLCELL_X1 FILLER_123_1230 ();
 FILLCELL_X4 FILLER_123_1234 ();
 FILLCELL_X2 FILLER_123_1238 ();
 FILLCELL_X16 FILLER_124_1 ();
 FILLCELL_X8 FILLER_124_17 ();
 FILLCELL_X32 FILLER_124_49 ();
 FILLCELL_X2 FILLER_124_81 ();
 FILLCELL_X1 FILLER_124_83 ();
 FILLCELL_X2 FILLER_124_115 ();
 FILLCELL_X1 FILLER_124_117 ();
 FILLCELL_X8 FILLER_124_125 ();
 FILLCELL_X2 FILLER_124_133 ();
 FILLCELL_X1 FILLER_124_135 ();
 FILLCELL_X16 FILLER_124_174 ();
 FILLCELL_X2 FILLER_124_190 ();
 FILLCELL_X8 FILLER_124_209 ();
 FILLCELL_X2 FILLER_124_241 ();
 FILLCELL_X4 FILLER_124_250 ();
 FILLCELL_X1 FILLER_124_254 ();
 FILLCELL_X16 FILLER_124_269 ();
 FILLCELL_X1 FILLER_124_285 ();
 FILLCELL_X8 FILLER_124_310 ();
 FILLCELL_X2 FILLER_124_318 ();
 FILLCELL_X1 FILLER_124_320 ();
 FILLCELL_X2 FILLER_124_328 ();
 FILLCELL_X1 FILLER_124_330 ();
 FILLCELL_X1 FILLER_124_348 ();
 FILLCELL_X8 FILLER_124_356 ();
 FILLCELL_X4 FILLER_124_364 ();
 FILLCELL_X1 FILLER_124_408 ();
 FILLCELL_X16 FILLER_124_423 ();
 FILLCELL_X4 FILLER_124_439 ();
 FILLCELL_X1 FILLER_124_443 ();
 FILLCELL_X32 FILLER_124_468 ();
 FILLCELL_X2 FILLER_124_500 ();
 FILLCELL_X16 FILLER_124_509 ();
 FILLCELL_X8 FILLER_124_525 ();
 FILLCELL_X2 FILLER_124_533 ();
 FILLCELL_X4 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_566 ();
 FILLCELL_X8 FILLER_124_598 ();
 FILLCELL_X2 FILLER_124_606 ();
 FILLCELL_X1 FILLER_124_615 ();
 FILLCELL_X8 FILLER_124_623 ();
 FILLCELL_X16 FILLER_124_632 ();
 FILLCELL_X4 FILLER_124_648 ();
 FILLCELL_X16 FILLER_124_666 ();
 FILLCELL_X8 FILLER_124_686 ();
 FILLCELL_X4 FILLER_124_694 ();
 FILLCELL_X2 FILLER_124_698 ();
 FILLCELL_X1 FILLER_124_709 ();
 FILLCELL_X8 FILLER_124_713 ();
 FILLCELL_X8 FILLER_124_740 ();
 FILLCELL_X8 FILLER_124_784 ();
 FILLCELL_X4 FILLER_124_792 ();
 FILLCELL_X1 FILLER_124_796 ();
 FILLCELL_X4 FILLER_124_800 ();
 FILLCELL_X2 FILLER_124_804 ();
 FILLCELL_X1 FILLER_124_845 ();
 FILLCELL_X1 FILLER_124_852 ();
 FILLCELL_X8 FILLER_124_857 ();
 FILLCELL_X2 FILLER_124_865 ();
 FILLCELL_X16 FILLER_124_886 ();
 FILLCELL_X4 FILLER_124_902 ();
 FILLCELL_X2 FILLER_124_932 ();
 FILLCELL_X8 FILLER_124_961 ();
 FILLCELL_X4 FILLER_124_969 ();
 FILLCELL_X1 FILLER_124_1012 ();
 FILLCELL_X1 FILLER_124_1018 ();
 FILLCELL_X1 FILLER_124_1030 ();
 FILLCELL_X2 FILLER_124_1036 ();
 FILLCELL_X2 FILLER_124_1044 ();
 FILLCELL_X2 FILLER_124_1051 ();
 FILLCELL_X1 FILLER_124_1053 ();
 FILLCELL_X8 FILLER_124_1060 ();
 FILLCELL_X1 FILLER_124_1068 ();
 FILLCELL_X4 FILLER_124_1072 ();
 FILLCELL_X1 FILLER_124_1076 ();
 FILLCELL_X4 FILLER_124_1083 ();
 FILLCELL_X32 FILLER_124_1104 ();
 FILLCELL_X2 FILLER_124_1136 ();
 FILLCELL_X1 FILLER_124_1162 ();
 FILLCELL_X2 FILLER_124_1204 ();
 FILLCELL_X1 FILLER_124_1206 ();
 FILLCELL_X2 FILLER_124_1210 ();
 FILLCELL_X4 FILLER_124_1236 ();
 FILLCELL_X16 FILLER_125_1 ();
 FILLCELL_X2 FILLER_125_17 ();
 FILLCELL_X16 FILLER_125_43 ();
 FILLCELL_X8 FILLER_125_59 ();
 FILLCELL_X2 FILLER_125_67 ();
 FILLCELL_X1 FILLER_125_69 ();
 FILLCELL_X8 FILLER_125_94 ();
 FILLCELL_X2 FILLER_125_102 ();
 FILLCELL_X4 FILLER_125_133 ();
 FILLCELL_X1 FILLER_125_137 ();
 FILLCELL_X16 FILLER_125_162 ();
 FILLCELL_X4 FILLER_125_178 ();
 FILLCELL_X4 FILLER_125_213 ();
 FILLCELL_X1 FILLER_125_217 ();
 FILLCELL_X2 FILLER_125_242 ();
 FILLCELL_X2 FILLER_125_261 ();
 FILLCELL_X1 FILLER_125_263 ();
 FILLCELL_X8 FILLER_125_273 ();
 FILLCELL_X2 FILLER_125_281 ();
 FILLCELL_X1 FILLER_125_283 ();
 FILLCELL_X8 FILLER_125_298 ();
 FILLCELL_X2 FILLER_125_306 ();
 FILLCELL_X8 FILLER_125_339 ();
 FILLCELL_X4 FILLER_125_347 ();
 FILLCELL_X32 FILLER_125_360 ();
 FILLCELL_X16 FILLER_125_392 ();
 FILLCELL_X2 FILLER_125_408 ();
 FILLCELL_X1 FILLER_125_410 ();
 FILLCELL_X8 FILLER_125_435 ();
 FILLCELL_X4 FILLER_125_452 ();
 FILLCELL_X1 FILLER_125_456 ();
 FILLCELL_X32 FILLER_125_474 ();
 FILLCELL_X32 FILLER_125_506 ();
 FILLCELL_X8 FILLER_125_538 ();
 FILLCELL_X4 FILLER_125_546 ();
 FILLCELL_X2 FILLER_125_550 ();
 FILLCELL_X8 FILLER_125_593 ();
 FILLCELL_X1 FILLER_125_601 ();
 FILLCELL_X1 FILLER_125_633 ();
 FILLCELL_X8 FILLER_125_643 ();
 FILLCELL_X2 FILLER_125_651 ();
 FILLCELL_X8 FILLER_125_688 ();
 FILLCELL_X2 FILLER_125_700 ();
 FILLCELL_X16 FILLER_125_712 ();
 FILLCELL_X2 FILLER_125_728 ();
 FILLCELL_X1 FILLER_125_744 ();
 FILLCELL_X1 FILLER_125_750 ();
 FILLCELL_X2 FILLER_125_756 ();
 FILLCELL_X2 FILLER_125_762 ();
 FILLCELL_X1 FILLER_125_770 ();
 FILLCELL_X32 FILLER_125_797 ();
 FILLCELL_X4 FILLER_125_829 ();
 FILLCELL_X2 FILLER_125_833 ();
 FILLCELL_X8 FILLER_125_862 ();
 FILLCELL_X4 FILLER_125_870 ();
 FILLCELL_X2 FILLER_125_874 ();
 FILLCELL_X4 FILLER_125_900 ();
 FILLCELL_X4 FILLER_125_909 ();
 FILLCELL_X2 FILLER_125_913 ();
 FILLCELL_X1 FILLER_125_915 ();
 FILLCELL_X4 FILLER_125_921 ();
 FILLCELL_X1 FILLER_125_925 ();
 FILLCELL_X4 FILLER_125_928 ();
 FILLCELL_X1 FILLER_125_932 ();
 FILLCELL_X4 FILLER_125_942 ();
 FILLCELL_X1 FILLER_125_946 ();
 FILLCELL_X4 FILLER_125_953 ();
 FILLCELL_X16 FILLER_125_961 ();
 FILLCELL_X2 FILLER_125_977 ();
 FILLCELL_X1 FILLER_125_979 ();
 FILLCELL_X2 FILLER_125_991 ();
 FILLCELL_X2 FILLER_125_1004 ();
 FILLCELL_X1 FILLER_125_1018 ();
 FILLCELL_X2 FILLER_125_1062 ();
 FILLCELL_X1 FILLER_125_1064 ();
 FILLCELL_X1 FILLER_125_1076 ();
 FILLCELL_X4 FILLER_125_1080 ();
 FILLCELL_X2 FILLER_125_1084 ();
 FILLCELL_X2 FILLER_125_1090 ();
 FILLCELL_X16 FILLER_125_1125 ();
 FILLCELL_X8 FILLER_125_1141 ();
 FILLCELL_X4 FILLER_125_1149 ();
 FILLCELL_X2 FILLER_125_1153 ();
 FILLCELL_X32 FILLER_125_1160 ();
 FILLCELL_X4 FILLER_125_1192 ();
 FILLCELL_X2 FILLER_125_1196 ();
 FILLCELL_X4 FILLER_126_1 ();
 FILLCELL_X4 FILLER_126_22 ();
 FILLCELL_X4 FILLER_126_33 ();
 FILLCELL_X2 FILLER_126_37 ();
 FILLCELL_X2 FILLER_126_46 ();
 FILLCELL_X2 FILLER_126_55 ();
 FILLCELL_X1 FILLER_126_57 ();
 FILLCELL_X8 FILLER_126_63 ();
 FILLCELL_X2 FILLER_126_85 ();
 FILLCELL_X1 FILLER_126_111 ();
 FILLCELL_X2 FILLER_126_119 ();
 FILLCELL_X2 FILLER_126_128 ();
 FILLCELL_X1 FILLER_126_130 ();
 FILLCELL_X4 FILLER_126_147 ();
 FILLCELL_X2 FILLER_126_151 ();
 FILLCELL_X1 FILLER_126_153 ();
 FILLCELL_X8 FILLER_126_161 ();
 FILLCELL_X1 FILLER_126_169 ();
 FILLCELL_X16 FILLER_126_177 ();
 FILLCELL_X2 FILLER_126_193 ();
 FILLCELL_X1 FILLER_126_195 ();
 FILLCELL_X8 FILLER_126_203 ();
 FILLCELL_X4 FILLER_126_211 ();
 FILLCELL_X2 FILLER_126_215 ();
 FILLCELL_X8 FILLER_126_224 ();
 FILLCELL_X4 FILLER_126_232 ();
 FILLCELL_X2 FILLER_126_236 ();
 FILLCELL_X1 FILLER_126_252 ();
 FILLCELL_X4 FILLER_126_260 ();
 FILLCELL_X1 FILLER_126_264 ();
 FILLCELL_X32 FILLER_126_290 ();
 FILLCELL_X8 FILLER_126_322 ();
 FILLCELL_X4 FILLER_126_330 ();
 FILLCELL_X1 FILLER_126_334 ();
 FILLCELL_X2 FILLER_126_356 ();
 FILLCELL_X1 FILLER_126_358 ();
 FILLCELL_X2 FILLER_126_368 ();
 FILLCELL_X1 FILLER_126_377 ();
 FILLCELL_X16 FILLER_126_394 ();
 FILLCELL_X1 FILLER_126_410 ();
 FILLCELL_X8 FILLER_126_425 ();
 FILLCELL_X4 FILLER_126_438 ();
 FILLCELL_X1 FILLER_126_442 ();
 FILLCELL_X4 FILLER_126_450 ();
 FILLCELL_X2 FILLER_126_454 ();
 FILLCELL_X32 FILLER_126_477 ();
 FILLCELL_X32 FILLER_126_509 ();
 FILLCELL_X8 FILLER_126_541 ();
 FILLCELL_X2 FILLER_126_549 ();
 FILLCELL_X2 FILLER_126_575 ();
 FILLCELL_X2 FILLER_126_580 ();
 FILLCELL_X4 FILLER_126_591 ();
 FILLCELL_X1 FILLER_126_595 ();
 FILLCELL_X1 FILLER_126_630 ();
 FILLCELL_X16 FILLER_126_632 ();
 FILLCELL_X4 FILLER_126_648 ();
 FILLCELL_X2 FILLER_126_652 ();
 FILLCELL_X4 FILLER_126_680 ();
 FILLCELL_X1 FILLER_126_684 ();
 FILLCELL_X16 FILLER_126_711 ();
 FILLCELL_X4 FILLER_126_727 ();
 FILLCELL_X2 FILLER_126_731 ();
 FILLCELL_X1 FILLER_126_733 ();
 FILLCELL_X16 FILLER_126_744 ();
 FILLCELL_X8 FILLER_126_760 ();
 FILLCELL_X4 FILLER_126_768 ();
 FILLCELL_X1 FILLER_126_772 ();
 FILLCELL_X2 FILLER_126_791 ();
 FILLCELL_X1 FILLER_126_793 ();
 FILLCELL_X4 FILLER_126_829 ();
 FILLCELL_X2 FILLER_126_833 ();
 FILLCELL_X1 FILLER_126_835 ();
 FILLCELL_X2 FILLER_126_852 ();
 FILLCELL_X1 FILLER_126_854 ();
 FILLCELL_X4 FILLER_126_862 ();
 FILLCELL_X8 FILLER_126_874 ();
 FILLCELL_X2 FILLER_126_887 ();
 FILLCELL_X8 FILLER_126_906 ();
 FILLCELL_X4 FILLER_126_932 ();
 FILLCELL_X8 FILLER_126_943 ();
 FILLCELL_X4 FILLER_126_951 ();
 FILLCELL_X1 FILLER_126_955 ();
 FILLCELL_X2 FILLER_126_964 ();
 FILLCELL_X1 FILLER_126_966 ();
 FILLCELL_X4 FILLER_126_975 ();
 FILLCELL_X2 FILLER_126_979 ();
 FILLCELL_X8 FILLER_126_992 ();
 FILLCELL_X4 FILLER_126_1000 ();
 FILLCELL_X1 FILLER_126_1004 ();
 FILLCELL_X2 FILLER_126_1009 ();
 FILLCELL_X2 FILLER_126_1026 ();
 FILLCELL_X2 FILLER_126_1033 ();
 FILLCELL_X2 FILLER_126_1039 ();
 FILLCELL_X1 FILLER_126_1041 ();
 FILLCELL_X1 FILLER_126_1048 ();
 FILLCELL_X8 FILLER_126_1074 ();
 FILLCELL_X2 FILLER_126_1082 ();
 FILLCELL_X1 FILLER_126_1084 ();
 FILLCELL_X4 FILLER_126_1092 ();
 FILLCELL_X2 FILLER_126_1108 ();
 FILLCELL_X1 FILLER_126_1114 ();
 FILLCELL_X16 FILLER_126_1118 ();
 FILLCELL_X4 FILLER_126_1134 ();
 FILLCELL_X4 FILLER_126_1193 ();
 FILLCELL_X1 FILLER_126_1197 ();
 FILLCELL_X1 FILLER_126_1239 ();
 FILLCELL_X1 FILLER_127_1 ();
 FILLCELL_X16 FILLER_127_29 ();
 FILLCELL_X4 FILLER_127_45 ();
 FILLCELL_X2 FILLER_127_49 ();
 FILLCELL_X2 FILLER_127_75 ();
 FILLCELL_X1 FILLER_127_77 ();
 FILLCELL_X2 FILLER_127_85 ();
 FILLCELL_X8 FILLER_127_94 ();
 FILLCELL_X4 FILLER_127_102 ();
 FILLCELL_X2 FILLER_127_126 ();
 FILLCELL_X1 FILLER_127_128 ();
 FILLCELL_X8 FILLER_127_136 ();
 FILLCELL_X2 FILLER_127_144 ();
 FILLCELL_X4 FILLER_127_185 ();
 FILLCELL_X2 FILLER_127_189 ();
 FILLCELL_X8 FILLER_127_222 ();
 FILLCELL_X4 FILLER_127_230 ();
 FILLCELL_X1 FILLER_127_234 ();
 FILLCELL_X16 FILLER_127_259 ();
 FILLCELL_X4 FILLER_127_275 ();
 FILLCELL_X1 FILLER_127_279 ();
 FILLCELL_X1 FILLER_127_287 ();
 FILLCELL_X1 FILLER_127_305 ();
 FILLCELL_X1 FILLER_127_320 ();
 FILLCELL_X8 FILLER_127_349 ();
 FILLCELL_X4 FILLER_127_357 ();
 FILLCELL_X2 FILLER_127_361 ();
 FILLCELL_X4 FILLER_127_397 ();
 FILLCELL_X2 FILLER_127_401 ();
 FILLCELL_X8 FILLER_127_427 ();
 FILLCELL_X1 FILLER_127_435 ();
 FILLCELL_X2 FILLER_127_443 ();
 FILLCELL_X1 FILLER_127_445 ();
 FILLCELL_X32 FILLER_127_470 ();
 FILLCELL_X16 FILLER_127_502 ();
 FILLCELL_X8 FILLER_127_518 ();
 FILLCELL_X4 FILLER_127_526 ();
 FILLCELL_X2 FILLER_127_530 ();
 FILLCELL_X8 FILLER_127_541 ();
 FILLCELL_X2 FILLER_127_549 ();
 FILLCELL_X1 FILLER_127_585 ();
 FILLCELL_X16 FILLER_127_590 ();
 FILLCELL_X8 FILLER_127_630 ();
 FILLCELL_X4 FILLER_127_638 ();
 FILLCELL_X2 FILLER_127_642 ();
 FILLCELL_X1 FILLER_127_644 ();
 FILLCELL_X1 FILLER_127_680 ();
 FILLCELL_X16 FILLER_127_734 ();
 FILLCELL_X1 FILLER_127_750 ();
 FILLCELL_X4 FILLER_127_758 ();
 FILLCELL_X2 FILLER_127_762 ();
 FILLCELL_X1 FILLER_127_764 ();
 FILLCELL_X32 FILLER_127_780 ();
 FILLCELL_X4 FILLER_127_812 ();
 FILLCELL_X2 FILLER_127_816 ();
 FILLCELL_X1 FILLER_127_818 ();
 FILLCELL_X16 FILLER_127_821 ();
 FILLCELL_X2 FILLER_127_840 ();
 FILLCELL_X1 FILLER_127_842 ();
 FILLCELL_X8 FILLER_127_863 ();
 FILLCELL_X1 FILLER_127_883 ();
 FILLCELL_X2 FILLER_127_888 ();
 FILLCELL_X4 FILLER_127_895 ();
 FILLCELL_X1 FILLER_127_899 ();
 FILLCELL_X16 FILLER_127_905 ();
 FILLCELL_X1 FILLER_127_925 ();
 FILLCELL_X4 FILLER_127_929 ();
 FILLCELL_X2 FILLER_127_933 ();
 FILLCELL_X1 FILLER_127_935 ();
 FILLCELL_X8 FILLER_127_940 ();
 FILLCELL_X4 FILLER_127_948 ();
 FILLCELL_X2 FILLER_127_952 ();
 FILLCELL_X1 FILLER_127_973 ();
 FILLCELL_X4 FILLER_127_978 ();
 FILLCELL_X8 FILLER_127_988 ();
 FILLCELL_X4 FILLER_127_996 ();
 FILLCELL_X2 FILLER_127_1000 ();
 FILLCELL_X4 FILLER_127_1007 ();
 FILLCELL_X2 FILLER_127_1015 ();
 FILLCELL_X1 FILLER_127_1024 ();
 FILLCELL_X4 FILLER_127_1033 ();
 FILLCELL_X1 FILLER_127_1037 ();
 FILLCELL_X1 FILLER_127_1042 ();
 FILLCELL_X4 FILLER_127_1046 ();
 FILLCELL_X8 FILLER_127_1054 ();
 FILLCELL_X2 FILLER_127_1062 ();
 FILLCELL_X1 FILLER_127_1064 ();
 FILLCELL_X16 FILLER_127_1074 ();
 FILLCELL_X2 FILLER_127_1090 ();
 FILLCELL_X8 FILLER_127_1095 ();
 FILLCELL_X2 FILLER_127_1103 ();
 FILLCELL_X4 FILLER_127_1134 ();
 FILLCELL_X2 FILLER_127_1138 ();
 FILLCELL_X1 FILLER_127_1140 ();
 FILLCELL_X4 FILLER_127_1158 ();
 FILLCELL_X1 FILLER_127_1162 ();
 FILLCELL_X4 FILLER_127_1204 ();
 FILLCELL_X1 FILLER_127_1227 ();
 FILLCELL_X2 FILLER_128_1 ();
 FILLCELL_X1 FILLER_128_3 ();
 FILLCELL_X4 FILLER_128_11 ();
 FILLCELL_X2 FILLER_128_15 ();
 FILLCELL_X8 FILLER_128_24 ();
 FILLCELL_X2 FILLER_128_32 ();
 FILLCELL_X1 FILLER_128_34 ();
 FILLCELL_X1 FILLER_128_59 ();
 FILLCELL_X16 FILLER_128_84 ();
 FILLCELL_X4 FILLER_128_100 ();
 FILLCELL_X2 FILLER_128_104 ();
 FILLCELL_X1 FILLER_128_106 ();
 FILLCELL_X2 FILLER_128_138 ();
 FILLCELL_X1 FILLER_128_140 ();
 FILLCELL_X1 FILLER_128_150 ();
 FILLCELL_X2 FILLER_128_184 ();
 FILLCELL_X8 FILLER_128_195 ();
 FILLCELL_X4 FILLER_128_203 ();
 FILLCELL_X1 FILLER_128_207 ();
 FILLCELL_X32 FILLER_128_232 ();
 FILLCELL_X16 FILLER_128_264 ();
 FILLCELL_X4 FILLER_128_280 ();
 FILLCELL_X1 FILLER_128_284 ();
 FILLCELL_X8 FILLER_128_360 ();
 FILLCELL_X2 FILLER_128_368 ();
 FILLCELL_X1 FILLER_128_394 ();
 FILLCELL_X1 FILLER_128_402 ();
 FILLCELL_X2 FILLER_128_410 ();
 FILLCELL_X4 FILLER_128_429 ();
 FILLCELL_X2 FILLER_128_450 ();
 FILLCELL_X4 FILLER_128_459 ();
 FILLCELL_X16 FILLER_128_487 ();
 FILLCELL_X8 FILLER_128_503 ();
 FILLCELL_X1 FILLER_128_511 ();
 FILLCELL_X8 FILLER_128_519 ();
 FILLCELL_X4 FILLER_128_527 ();
 FILLCELL_X8 FILLER_128_548 ();
 FILLCELL_X1 FILLER_128_556 ();
 FILLCELL_X1 FILLER_128_578 ();
 FILLCELL_X1 FILLER_128_584 ();
 FILLCELL_X16 FILLER_128_589 ();
 FILLCELL_X8 FILLER_128_605 ();
 FILLCELL_X8 FILLER_128_620 ();
 FILLCELL_X2 FILLER_128_628 ();
 FILLCELL_X1 FILLER_128_630 ();
 FILLCELL_X4 FILLER_128_632 ();
 FILLCELL_X2 FILLER_128_636 ();
 FILLCELL_X1 FILLER_128_638 ();
 FILLCELL_X1 FILLER_128_652 ();
 FILLCELL_X1 FILLER_128_667 ();
 FILLCELL_X8 FILLER_128_672 ();
 FILLCELL_X2 FILLER_128_680 ();
 FILLCELL_X1 FILLER_128_686 ();
 FILLCELL_X1 FILLER_128_712 ();
 FILLCELL_X2 FILLER_128_718 ();
 FILLCELL_X2 FILLER_128_723 ();
 FILLCELL_X1 FILLER_128_732 ();
 FILLCELL_X2 FILLER_128_754 ();
 FILLCELL_X1 FILLER_128_756 ();
 FILLCELL_X4 FILLER_128_764 ();
 FILLCELL_X2 FILLER_128_768 ();
 FILLCELL_X2 FILLER_128_780 ();
 FILLCELL_X8 FILLER_128_789 ();
 FILLCELL_X2 FILLER_128_797 ();
 FILLCELL_X16 FILLER_128_851 ();
 FILLCELL_X1 FILLER_128_887 ();
 FILLCELL_X8 FILLER_128_905 ();
 FILLCELL_X4 FILLER_128_913 ();
 FILLCELL_X1 FILLER_128_917 ();
 FILLCELL_X8 FILLER_128_934 ();
 FILLCELL_X1 FILLER_128_945 ();
 FILLCELL_X2 FILLER_128_952 ();
 FILLCELL_X2 FILLER_128_957 ();
 FILLCELL_X1 FILLER_128_959 ();
 FILLCELL_X2 FILLER_128_972 ();
 FILLCELL_X16 FILLER_128_978 ();
 FILLCELL_X4 FILLER_128_994 ();
 FILLCELL_X1 FILLER_128_998 ();
 FILLCELL_X1 FILLER_128_1005 ();
 FILLCELL_X16 FILLER_128_1016 ();
 FILLCELL_X1 FILLER_128_1032 ();
 FILLCELL_X2 FILLER_128_1039 ();
 FILLCELL_X2 FILLER_128_1044 ();
 FILLCELL_X4 FILLER_128_1049 ();
 FILLCELL_X1 FILLER_128_1056 ();
 FILLCELL_X8 FILLER_128_1060 ();
 FILLCELL_X4 FILLER_128_1074 ();
 FILLCELL_X16 FILLER_128_1081 ();
 FILLCELL_X2 FILLER_128_1115 ();
 FILLCELL_X4 FILLER_128_1130 ();
 FILLCELL_X2 FILLER_128_1134 ();
 FILLCELL_X1 FILLER_128_1152 ();
 FILLCELL_X16 FILLER_128_1202 ();
 FILLCELL_X4 FILLER_128_1221 ();
 FILLCELL_X8 FILLER_129_1 ();
 FILLCELL_X2 FILLER_129_9 ();
 FILLCELL_X1 FILLER_129_11 ();
 FILLCELL_X1 FILLER_129_43 ();
 FILLCELL_X4 FILLER_129_55 ();
 FILLCELL_X1 FILLER_129_59 ();
 FILLCELL_X16 FILLER_129_74 ();
 FILLCELL_X8 FILLER_129_90 ();
 FILLCELL_X1 FILLER_129_98 ();
 FILLCELL_X1 FILLER_129_116 ();
 FILLCELL_X4 FILLER_129_131 ();
 FILLCELL_X8 FILLER_129_142 ();
 FILLCELL_X1 FILLER_129_157 ();
 FILLCELL_X4 FILLER_129_172 ();
 FILLCELL_X1 FILLER_129_176 ();
 FILLCELL_X8 FILLER_129_200 ();
 FILLCELL_X4 FILLER_129_208 ();
 FILLCELL_X4 FILLER_129_219 ();
 FILLCELL_X1 FILLER_129_223 ();
 FILLCELL_X4 FILLER_129_228 ();
 FILLCELL_X1 FILLER_129_232 ();
 FILLCELL_X16 FILLER_129_257 ();
 FILLCELL_X8 FILLER_129_273 ();
 FILLCELL_X4 FILLER_129_281 ();
 FILLCELL_X2 FILLER_129_292 ();
 FILLCELL_X1 FILLER_129_301 ();
 FILLCELL_X4 FILLER_129_309 ();
 FILLCELL_X2 FILLER_129_313 ();
 FILLCELL_X2 FILLER_129_339 ();
 FILLCELL_X8 FILLER_129_348 ();
 FILLCELL_X8 FILLER_129_363 ();
 FILLCELL_X2 FILLER_129_371 ();
 FILLCELL_X4 FILLER_129_404 ();
 FILLCELL_X2 FILLER_129_408 ();
 FILLCELL_X4 FILLER_129_417 ();
 FILLCELL_X2 FILLER_129_421 ();
 FILLCELL_X1 FILLER_129_423 ();
 FILLCELL_X32 FILLER_129_455 ();
 FILLCELL_X32 FILLER_129_487 ();
 FILLCELL_X8 FILLER_129_519 ();
 FILLCELL_X2 FILLER_129_527 ();
 FILLCELL_X4 FILLER_129_546 ();
 FILLCELL_X1 FILLER_129_550 ();
 FILLCELL_X2 FILLER_129_565 ();
 FILLCELL_X1 FILLER_129_567 ();
 FILLCELL_X8 FILLER_129_584 ();
 FILLCELL_X4 FILLER_129_592 ();
 FILLCELL_X2 FILLER_129_599 ();
 FILLCELL_X32 FILLER_129_608 ();
 FILLCELL_X4 FILLER_129_666 ();
 FILLCELL_X4 FILLER_129_705 ();
 FILLCELL_X2 FILLER_129_709 ();
 FILLCELL_X1 FILLER_129_720 ();
 FILLCELL_X1 FILLER_129_738 ();
 FILLCELL_X1 FILLER_129_744 ();
 FILLCELL_X2 FILLER_129_754 ();
 FILLCELL_X1 FILLER_129_765 ();
 FILLCELL_X1 FILLER_129_769 ();
 FILLCELL_X8 FILLER_129_774 ();
 FILLCELL_X2 FILLER_129_786 ();
 FILLCELL_X1 FILLER_129_788 ();
 FILLCELL_X16 FILLER_129_791 ();
 FILLCELL_X4 FILLER_129_822 ();
 FILLCELL_X32 FILLER_129_830 ();
 FILLCELL_X1 FILLER_129_880 ();
 FILLCELL_X16 FILLER_129_902 ();
 FILLCELL_X1 FILLER_129_918 ();
 FILLCELL_X8 FILLER_129_943 ();
 FILLCELL_X2 FILLER_129_951 ();
 FILLCELL_X1 FILLER_129_956 ();
 FILLCELL_X16 FILLER_129_963 ();
 FILLCELL_X8 FILLER_129_979 ();
 FILLCELL_X4 FILLER_129_994 ();
 FILLCELL_X1 FILLER_129_998 ();
 FILLCELL_X8 FILLER_129_1006 ();
 FILLCELL_X8 FILLER_129_1039 ();
 FILLCELL_X4 FILLER_129_1047 ();
 FILLCELL_X2 FILLER_129_1051 ();
 FILLCELL_X8 FILLER_129_1060 ();
 FILLCELL_X4 FILLER_129_1068 ();
 FILLCELL_X2 FILLER_129_1072 ();
 FILLCELL_X1 FILLER_129_1074 ();
 FILLCELL_X8 FILLER_129_1082 ();
 FILLCELL_X1 FILLER_129_1090 ();
 FILLCELL_X8 FILLER_129_1117 ();
 FILLCELL_X4 FILLER_129_1125 ();
 FILLCELL_X2 FILLER_129_1129 ();
 FILLCELL_X1 FILLER_129_1131 ();
 FILLCELL_X4 FILLER_129_1137 ();
 FILLCELL_X8 FILLER_129_1146 ();
 FILLCELL_X4 FILLER_129_1154 ();
 FILLCELL_X2 FILLER_129_1158 ();
 FILLCELL_X1 FILLER_129_1160 ();
 FILLCELL_X8 FILLER_129_1164 ();
 FILLCELL_X2 FILLER_129_1172 ();
 FILLCELL_X1 FILLER_129_1191 ();
 FILLCELL_X4 FILLER_129_1209 ();
 FILLCELL_X1 FILLER_129_1213 ();
 FILLCELL_X4 FILLER_129_1235 ();
 FILLCELL_X1 FILLER_129_1239 ();
 FILLCELL_X8 FILLER_130_1 ();
 FILLCELL_X4 FILLER_130_9 ();
 FILLCELL_X1 FILLER_130_13 ();
 FILLCELL_X4 FILLER_130_31 ();
 FILLCELL_X2 FILLER_130_35 ();
 FILLCELL_X8 FILLER_130_42 ();
 FILLCELL_X4 FILLER_130_50 ();
 FILLCELL_X2 FILLER_130_54 ();
 FILLCELL_X16 FILLER_130_63 ();
 FILLCELL_X8 FILLER_130_79 ();
 FILLCELL_X4 FILLER_130_87 ();
 FILLCELL_X2 FILLER_130_91 ();
 FILLCELL_X4 FILLER_130_103 ();
 FILLCELL_X1 FILLER_130_107 ();
 FILLCELL_X2 FILLER_130_115 ();
 FILLCELL_X8 FILLER_130_141 ();
 FILLCELL_X2 FILLER_130_149 ();
 FILLCELL_X1 FILLER_130_151 ();
 FILLCELL_X32 FILLER_130_169 ();
 FILLCELL_X2 FILLER_130_201 ();
 FILLCELL_X8 FILLER_130_210 ();
 FILLCELL_X8 FILLER_130_225 ();
 FILLCELL_X1 FILLER_130_233 ();
 FILLCELL_X8 FILLER_130_241 ();
 FILLCELL_X4 FILLER_130_249 ();
 FILLCELL_X2 FILLER_130_253 ();
 FILLCELL_X1 FILLER_130_255 ();
 FILLCELL_X2 FILLER_130_270 ();
 FILLCELL_X4 FILLER_130_296 ();
 FILLCELL_X2 FILLER_130_300 ();
 FILLCELL_X1 FILLER_130_302 ();
 FILLCELL_X8 FILLER_130_307 ();
 FILLCELL_X4 FILLER_130_315 ();
 FILLCELL_X32 FILLER_130_324 ();
 FILLCELL_X16 FILLER_130_356 ();
 FILLCELL_X8 FILLER_130_372 ();
 FILLCELL_X4 FILLER_130_380 ();
 FILLCELL_X1 FILLER_130_384 ();
 FILLCELL_X32 FILLER_130_390 ();
 FILLCELL_X16 FILLER_130_422 ();
 FILLCELL_X8 FILLER_130_438 ();
 FILLCELL_X2 FILLER_130_446 ();
 FILLCELL_X32 FILLER_130_455 ();
 FILLCELL_X32 FILLER_130_487 ();
 FILLCELL_X8 FILLER_130_519 ();
 FILLCELL_X2 FILLER_130_546 ();
 FILLCELL_X1 FILLER_130_548 ();
 FILLCELL_X1 FILLER_130_569 ();
 FILLCELL_X1 FILLER_130_575 ();
 FILLCELL_X1 FILLER_130_582 ();
 FILLCELL_X1 FILLER_130_585 ();
 FILLCELL_X8 FILLER_130_612 ();
 FILLCELL_X1 FILLER_130_620 ();
 FILLCELL_X1 FILLER_130_630 ();
 FILLCELL_X4 FILLER_130_632 ();
 FILLCELL_X8 FILLER_130_660 ();
 FILLCELL_X4 FILLER_130_668 ();
 FILLCELL_X1 FILLER_130_672 ();
 FILLCELL_X8 FILLER_130_697 ();
 FILLCELL_X2 FILLER_130_705 ();
 FILLCELL_X4 FILLER_130_711 ();
 FILLCELL_X2 FILLER_130_715 ();
 FILLCELL_X1 FILLER_130_717 ();
 FILLCELL_X8 FILLER_130_723 ();
 FILLCELL_X4 FILLER_130_731 ();
 FILLCELL_X1 FILLER_130_759 ();
 FILLCELL_X2 FILLER_130_764 ();
 FILLCELL_X1 FILLER_130_770 ();
 FILLCELL_X2 FILLER_130_780 ();
 FILLCELL_X32 FILLER_130_800 ();
 FILLCELL_X4 FILLER_130_832 ();
 FILLCELL_X1 FILLER_130_836 ();
 FILLCELL_X16 FILLER_130_842 ();
 FILLCELL_X4 FILLER_130_858 ();
 FILLCELL_X2 FILLER_130_862 ();
 FILLCELL_X1 FILLER_130_864 ();
 FILLCELL_X2 FILLER_130_886 ();
 FILLCELL_X16 FILLER_130_900 ();
 FILLCELL_X4 FILLER_130_916 ();
 FILLCELL_X1 FILLER_130_920 ();
 FILLCELL_X8 FILLER_130_936 ();
 FILLCELL_X2 FILLER_130_944 ();
 FILLCELL_X4 FILLER_130_963 ();
 FILLCELL_X2 FILLER_130_967 ();
 FILLCELL_X1 FILLER_130_969 ();
 FILLCELL_X2 FILLER_130_981 ();
 FILLCELL_X4 FILLER_130_992 ();
 FILLCELL_X2 FILLER_130_996 ();
 FILLCELL_X4 FILLER_130_1011 ();
 FILLCELL_X1 FILLER_130_1015 ();
 FILLCELL_X2 FILLER_130_1020 ();
 FILLCELL_X1 FILLER_130_1038 ();
 FILLCELL_X16 FILLER_130_1042 ();
 FILLCELL_X4 FILLER_130_1058 ();
 FILLCELL_X1 FILLER_130_1062 ();
 FILLCELL_X1 FILLER_130_1067 ();
 FILLCELL_X2 FILLER_130_1070 ();
 FILLCELL_X8 FILLER_130_1086 ();
 FILLCELL_X1 FILLER_130_1094 ();
 FILLCELL_X1 FILLER_130_1114 ();
 FILLCELL_X2 FILLER_130_1122 ();
 FILLCELL_X4 FILLER_130_1144 ();
 FILLCELL_X2 FILLER_130_1148 ();
 FILLCELL_X1 FILLER_130_1150 ();
 FILLCELL_X16 FILLER_130_1158 ();
 FILLCELL_X4 FILLER_130_1174 ();
 FILLCELL_X2 FILLER_130_1203 ();
 FILLCELL_X1 FILLER_130_1239 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X8 FILLER_131_33 ();
 FILLCELL_X4 FILLER_131_41 ();
 FILLCELL_X16 FILLER_131_86 ();
 FILLCELL_X32 FILLER_131_119 ();
 FILLCELL_X32 FILLER_131_151 ();
 FILLCELL_X8 FILLER_131_183 ();
 FILLCELL_X2 FILLER_131_191 ();
 FILLCELL_X1 FILLER_131_215 ();
 FILLCELL_X2 FILLER_131_247 ();
 FILLCELL_X8 FILLER_131_273 ();
 FILLCELL_X16 FILLER_131_288 ();
 FILLCELL_X4 FILLER_131_304 ();
 FILLCELL_X1 FILLER_131_308 ();
 FILLCELL_X32 FILLER_131_313 ();
 FILLCELL_X32 FILLER_131_345 ();
 FILLCELL_X16 FILLER_131_377 ();
 FILLCELL_X4 FILLER_131_393 ();
 FILLCELL_X2 FILLER_131_397 ();
 FILLCELL_X1 FILLER_131_399 ();
 FILLCELL_X2 FILLER_131_407 ();
 FILLCELL_X1 FILLER_131_409 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X8 FILLER_131_513 ();
 FILLCELL_X4 FILLER_131_521 ();
 FILLCELL_X2 FILLER_131_525 ();
 FILLCELL_X1 FILLER_131_527 ();
 FILLCELL_X4 FILLER_131_545 ();
 FILLCELL_X2 FILLER_131_549 ();
 FILLCELL_X1 FILLER_131_551 ();
 FILLCELL_X4 FILLER_131_572 ();
 FILLCELL_X2 FILLER_131_576 ();
 FILLCELL_X1 FILLER_131_616 ();
 FILLCELL_X8 FILLER_131_656 ();
 FILLCELL_X4 FILLER_131_664 ();
 FILLCELL_X2 FILLER_131_668 ();
 FILLCELL_X1 FILLER_131_670 ();
 FILLCELL_X2 FILLER_131_717 ();
 FILLCELL_X8 FILLER_131_733 ();
 FILLCELL_X4 FILLER_131_741 ();
 FILLCELL_X16 FILLER_131_765 ();
 FILLCELL_X8 FILLER_131_781 ();
 FILLCELL_X1 FILLER_131_789 ();
 FILLCELL_X4 FILLER_131_807 ();
 FILLCELL_X2 FILLER_131_811 ();
 FILLCELL_X1 FILLER_131_813 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X1 FILLER_131_888 ();
 FILLCELL_X2 FILLER_131_902 ();
 FILLCELL_X1 FILLER_131_909 ();
 FILLCELL_X4 FILLER_131_917 ();
 FILLCELL_X2 FILLER_131_925 ();
 FILLCELL_X1 FILLER_131_927 ();
 FILLCELL_X1 FILLER_131_932 ();
 FILLCELL_X8 FILLER_131_937 ();
 FILLCELL_X2 FILLER_131_1021 ();
 FILLCELL_X8 FILLER_131_1048 ();
 FILLCELL_X2 FILLER_131_1109 ();
 FILLCELL_X4 FILLER_131_1128 ();
 FILLCELL_X2 FILLER_131_1132 ();
 FILLCELL_X1 FILLER_131_1134 ();
 FILLCELL_X8 FILLER_131_1159 ();
 FILLCELL_X4 FILLER_131_1167 ();
 FILLCELL_X2 FILLER_131_1171 ();
 FILLCELL_X1 FILLER_131_1173 ();
 FILLCELL_X1 FILLER_131_1226 ();
 FILLCELL_X1 FILLER_131_1239 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X4 FILLER_132_65 ();
 FILLCELL_X1 FILLER_132_69 ();
 FILLCELL_X16 FILLER_132_94 ();
 FILLCELL_X1 FILLER_132_124 ();
 FILLCELL_X16 FILLER_132_132 ();
 FILLCELL_X16 FILLER_132_165 ();
 FILLCELL_X4 FILLER_132_181 ();
 FILLCELL_X1 FILLER_132_185 ();
 FILLCELL_X32 FILLER_132_234 ();
 FILLCELL_X8 FILLER_132_266 ();
 FILLCELL_X4 FILLER_132_274 ();
 FILLCELL_X1 FILLER_132_278 ();
 FILLCELL_X8 FILLER_132_296 ();
 FILLCELL_X4 FILLER_132_304 ();
 FILLCELL_X2 FILLER_132_308 ();
 FILLCELL_X1 FILLER_132_310 ();
 FILLCELL_X2 FILLER_132_318 ();
 FILLCELL_X1 FILLER_132_327 ();
 FILLCELL_X2 FILLER_132_335 ();
 FILLCELL_X2 FILLER_132_344 ();
 FILLCELL_X2 FILLER_132_353 ();
 FILLCELL_X4 FILLER_132_362 ();
 FILLCELL_X8 FILLER_132_373 ();
 FILLCELL_X4 FILLER_132_381 ();
 FILLCELL_X1 FILLER_132_385 ();
 FILLCELL_X4 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_442 ();
 FILLCELL_X32 FILLER_132_474 ();
 FILLCELL_X32 FILLER_132_506 ();
 FILLCELL_X32 FILLER_132_538 ();
 FILLCELL_X8 FILLER_132_570 ();
 FILLCELL_X16 FILLER_132_608 ();
 FILLCELL_X4 FILLER_132_624 ();
 FILLCELL_X2 FILLER_132_628 ();
 FILLCELL_X1 FILLER_132_630 ();
 FILLCELL_X2 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_648 ();
 FILLCELL_X16 FILLER_132_680 ();
 FILLCELL_X4 FILLER_132_696 ();
 FILLCELL_X4 FILLER_132_717 ();
 FILLCELL_X1 FILLER_132_721 ();
 FILLCELL_X16 FILLER_132_770 ();
 FILLCELL_X2 FILLER_132_786 ();
 FILLCELL_X1 FILLER_132_788 ();
 FILLCELL_X1 FILLER_132_804 ();
 FILLCELL_X4 FILLER_132_812 ();
 FILLCELL_X8 FILLER_132_820 ();
 FILLCELL_X2 FILLER_132_828 ();
 FILLCELL_X8 FILLER_132_835 ();
 FILLCELL_X4 FILLER_132_843 ();
 FILLCELL_X1 FILLER_132_868 ();
 FILLCELL_X2 FILLER_132_875 ();
 FILLCELL_X1 FILLER_132_889 ();
 FILLCELL_X1 FILLER_132_897 ();
 FILLCELL_X4 FILLER_132_902 ();
 FILLCELL_X1 FILLER_132_906 ();
 FILLCELL_X1 FILLER_132_911 ();
 FILLCELL_X4 FILLER_132_922 ();
 FILLCELL_X2 FILLER_132_926 ();
 FILLCELL_X4 FILLER_132_936 ();
 FILLCELL_X2 FILLER_132_940 ();
 FILLCELL_X1 FILLER_132_942 ();
 FILLCELL_X1 FILLER_132_968 ();
 FILLCELL_X1 FILLER_132_982 ();
 FILLCELL_X4 FILLER_132_1017 ();
 FILLCELL_X2 FILLER_132_1021 ();
 FILLCELL_X4 FILLER_132_1050 ();
 FILLCELL_X2 FILLER_132_1095 ();
 FILLCELL_X1 FILLER_132_1103 ();
 FILLCELL_X2 FILLER_132_1107 ();
 FILLCELL_X2 FILLER_132_1113 ();
 FILLCELL_X16 FILLER_132_1120 ();
 FILLCELL_X2 FILLER_132_1160 ();
 FILLCELL_X4 FILLER_132_1169 ();
 FILLCELL_X2 FILLER_132_1173 ();
 FILLCELL_X1 FILLER_132_1209 ();
 FILLCELL_X1 FILLER_132_1235 ();
 FILLCELL_X1 FILLER_132_1239 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X8 FILLER_133_33 ();
 FILLCELL_X2 FILLER_133_65 ();
 FILLCELL_X1 FILLER_133_67 ();
 FILLCELL_X4 FILLER_133_75 ();
 FILLCELL_X2 FILLER_133_79 ();
 FILLCELL_X1 FILLER_133_81 ();
 FILLCELL_X8 FILLER_133_89 ();
 FILLCELL_X2 FILLER_133_131 ();
 FILLCELL_X4 FILLER_133_140 ();
 FILLCELL_X4 FILLER_133_151 ();
 FILLCELL_X2 FILLER_133_162 ();
 FILLCELL_X1 FILLER_133_164 ();
 FILLCELL_X16 FILLER_133_172 ();
 FILLCELL_X2 FILLER_133_188 ();
 FILLCELL_X1 FILLER_133_197 ();
 FILLCELL_X1 FILLER_133_205 ();
 FILLCELL_X8 FILLER_133_213 ();
 FILLCELL_X2 FILLER_133_221 ();
 FILLCELL_X1 FILLER_133_223 ();
 FILLCELL_X2 FILLER_133_248 ();
 FILLCELL_X8 FILLER_133_267 ();
 FILLCELL_X4 FILLER_133_275 ();
 FILLCELL_X2 FILLER_133_279 ();
 FILLCELL_X1 FILLER_133_281 ();
 FILLCELL_X2 FILLER_133_316 ();
 FILLCELL_X8 FILLER_133_383 ();
 FILLCELL_X2 FILLER_133_391 ();
 FILLCELL_X1 FILLER_133_393 ();
 FILLCELL_X2 FILLER_133_418 ();
 FILLCELL_X1 FILLER_133_420 ();
 FILLCELL_X2 FILLER_133_435 ();
 FILLCELL_X1 FILLER_133_437 ();
 FILLCELL_X32 FILLER_133_453 ();
 FILLCELL_X32 FILLER_133_485 ();
 FILLCELL_X4 FILLER_133_517 ();
 FILLCELL_X2 FILLER_133_521 ();
 FILLCELL_X32 FILLER_133_528 ();
 FILLCELL_X16 FILLER_133_560 ();
 FILLCELL_X8 FILLER_133_576 ();
 FILLCELL_X4 FILLER_133_584 ();
 FILLCELL_X2 FILLER_133_588 ();
 FILLCELL_X32 FILLER_133_593 ();
 FILLCELL_X4 FILLER_133_625 ();
 FILLCELL_X1 FILLER_133_629 ();
 FILLCELL_X16 FILLER_133_647 ();
 FILLCELL_X8 FILLER_133_663 ();
 FILLCELL_X1 FILLER_133_671 ();
 FILLCELL_X32 FILLER_133_679 ();
 FILLCELL_X2 FILLER_133_711 ();
 FILLCELL_X1 FILLER_133_713 ();
 FILLCELL_X4 FILLER_133_731 ();
 FILLCELL_X2 FILLER_133_735 ();
 FILLCELL_X1 FILLER_133_737 ();
 FILLCELL_X2 FILLER_133_755 ();
 FILLCELL_X1 FILLER_133_757 ();
 FILLCELL_X2 FILLER_133_762 ();
 FILLCELL_X1 FILLER_133_764 ();
 FILLCELL_X4 FILLER_133_772 ();
 FILLCELL_X2 FILLER_133_776 ();
 FILLCELL_X2 FILLER_133_785 ();
 FILLCELL_X1 FILLER_133_787 ();
 FILLCELL_X1 FILLER_133_821 ();
 FILLCELL_X8 FILLER_133_839 ();
 FILLCELL_X4 FILLER_133_847 ();
 FILLCELL_X1 FILLER_133_851 ();
 FILLCELL_X1 FILLER_133_881 ();
 FILLCELL_X4 FILLER_133_904 ();
 FILLCELL_X2 FILLER_133_908 ();
 FILLCELL_X1 FILLER_133_910 ();
 FILLCELL_X4 FILLER_133_916 ();
 FILLCELL_X1 FILLER_133_936 ();
 FILLCELL_X1 FILLER_133_939 ();
 FILLCELL_X2 FILLER_133_947 ();
 FILLCELL_X2 FILLER_133_953 ();
 FILLCELL_X2 FILLER_133_959 ();
 FILLCELL_X2 FILLER_133_966 ();
 FILLCELL_X2 FILLER_133_977 ();
 FILLCELL_X1 FILLER_133_979 ();
 FILLCELL_X2 FILLER_133_1024 ();
 FILLCELL_X16 FILLER_133_1049 ();
 FILLCELL_X4 FILLER_133_1093 ();
 FILLCELL_X2 FILLER_133_1097 ();
 FILLCELL_X1 FILLER_133_1124 ();
 FILLCELL_X8 FILLER_133_1132 ();
 FILLCELL_X4 FILLER_133_1140 ();
 FILLCELL_X1 FILLER_133_1144 ();
 FILLCELL_X8 FILLER_133_1152 ();
 FILLCELL_X4 FILLER_133_1160 ();
 FILLCELL_X1 FILLER_133_1181 ();
 FILLCELL_X2 FILLER_133_1185 ();
 FILLCELL_X4 FILLER_134_1 ();
 FILLCELL_X2 FILLER_134_5 ();
 FILLCELL_X8 FILLER_134_24 ();
 FILLCELL_X8 FILLER_134_87 ();
 FILLCELL_X1 FILLER_134_95 ();
 FILLCELL_X8 FILLER_134_103 ();
 FILLCELL_X4 FILLER_134_111 ();
 FILLCELL_X2 FILLER_134_115 ();
 FILLCELL_X2 FILLER_134_124 ();
 FILLCELL_X4 FILLER_134_140 ();
 FILLCELL_X2 FILLER_134_168 ();
 FILLCELL_X8 FILLER_134_184 ();
 FILLCELL_X2 FILLER_134_192 ();
 FILLCELL_X2 FILLER_134_211 ();
 FILLCELL_X16 FILLER_134_220 ();
 FILLCELL_X4 FILLER_134_243 ();
 FILLCELL_X1 FILLER_134_261 ();
 FILLCELL_X4 FILLER_134_269 ();
 FILLCELL_X2 FILLER_134_273 ();
 FILLCELL_X2 FILLER_134_287 ();
 FILLCELL_X1 FILLER_134_289 ();
 FILLCELL_X1 FILLER_134_304 ();
 FILLCELL_X8 FILLER_134_312 ();
 FILLCELL_X1 FILLER_134_320 ();
 FILLCELL_X2 FILLER_134_335 ();
 FILLCELL_X1 FILLER_134_337 ();
 FILLCELL_X16 FILLER_134_362 ();
 FILLCELL_X4 FILLER_134_378 ();
 FILLCELL_X32 FILLER_134_447 ();
 FILLCELL_X32 FILLER_134_479 ();
 FILLCELL_X32 FILLER_134_511 ();
 FILLCELL_X4 FILLER_134_543 ();
 FILLCELL_X2 FILLER_134_547 ();
 FILLCELL_X1 FILLER_134_549 ();
 FILLCELL_X16 FILLER_134_553 ();
 FILLCELL_X2 FILLER_134_569 ();
 FILLCELL_X32 FILLER_134_591 ();
 FILLCELL_X8 FILLER_134_623 ();
 FILLCELL_X4 FILLER_134_639 ();
 FILLCELL_X4 FILLER_134_650 ();
 FILLCELL_X2 FILLER_134_654 ();
 FILLCELL_X4 FILLER_134_663 ();
 FILLCELL_X8 FILLER_134_674 ();
 FILLCELL_X4 FILLER_134_682 ();
 FILLCELL_X1 FILLER_134_686 ();
 FILLCELL_X2 FILLER_134_711 ();
 FILLCELL_X16 FILLER_134_722 ();
 FILLCELL_X1 FILLER_134_738 ();
 FILLCELL_X8 FILLER_134_758 ();
 FILLCELL_X1 FILLER_134_766 ();
 FILLCELL_X8 FILLER_134_776 ();
 FILLCELL_X4 FILLER_134_784 ();
 FILLCELL_X2 FILLER_134_832 ();
 FILLCELL_X8 FILLER_134_905 ();
 FILLCELL_X2 FILLER_134_913 ();
 FILLCELL_X2 FILLER_134_945 ();
 FILLCELL_X1 FILLER_134_965 ();
 FILLCELL_X1 FILLER_134_979 ();
 FILLCELL_X1 FILLER_134_986 ();
 FILLCELL_X2 FILLER_134_1000 ();
 FILLCELL_X2 FILLER_134_1015 ();
 FILLCELL_X16 FILLER_134_1036 ();
 FILLCELL_X4 FILLER_134_1052 ();
 FILLCELL_X2 FILLER_134_1056 ();
 FILLCELL_X4 FILLER_134_1066 ();
 FILLCELL_X1 FILLER_134_1070 ();
 FILLCELL_X4 FILLER_134_1074 ();
 FILLCELL_X1 FILLER_134_1078 ();
 FILLCELL_X32 FILLER_134_1081 ();
 FILLCELL_X16 FILLER_134_1113 ();
 FILLCELL_X8 FILLER_134_1129 ();
 FILLCELL_X4 FILLER_134_1137 ();
 FILLCELL_X8 FILLER_134_1165 ();
 FILLCELL_X2 FILLER_134_1173 ();
 FILLCELL_X2 FILLER_134_1192 ();
 FILLCELL_X1 FILLER_134_1216 ();
 FILLCELL_X2 FILLER_134_1220 ();
 FILLCELL_X1 FILLER_134_1222 ();
 FILLCELL_X8 FILLER_135_1 ();
 FILLCELL_X4 FILLER_135_33 ();
 FILLCELL_X2 FILLER_135_37 ();
 FILLCELL_X2 FILLER_135_46 ();
 FILLCELL_X1 FILLER_135_48 ();
 FILLCELL_X32 FILLER_135_80 ();
 FILLCELL_X4 FILLER_135_112 ();
 FILLCELL_X1 FILLER_135_116 ();
 FILLCELL_X16 FILLER_135_139 ();
 FILLCELL_X4 FILLER_135_155 ();
 FILLCELL_X1 FILLER_135_159 ();
 FILLCELL_X8 FILLER_135_184 ();
 FILLCELL_X2 FILLER_135_192 ();
 FILLCELL_X8 FILLER_135_201 ();
 FILLCELL_X2 FILLER_135_209 ();
 FILLCELL_X32 FILLER_135_218 ();
 FILLCELL_X4 FILLER_135_250 ();
 FILLCELL_X1 FILLER_135_254 ();
 FILLCELL_X2 FILLER_135_272 ();
 FILLCELL_X1 FILLER_135_274 ();
 FILLCELL_X4 FILLER_135_292 ();
 FILLCELL_X2 FILLER_135_296 ();
 FILLCELL_X4 FILLER_135_322 ();
 FILLCELL_X8 FILLER_135_343 ();
 FILLCELL_X1 FILLER_135_351 ();
 FILLCELL_X32 FILLER_135_360 ();
 FILLCELL_X32 FILLER_135_392 ();
 FILLCELL_X32 FILLER_135_424 ();
 FILLCELL_X32 FILLER_135_456 ();
 FILLCELL_X32 FILLER_135_488 ();
 FILLCELL_X8 FILLER_135_520 ();
 FILLCELL_X4 FILLER_135_528 ();
 FILLCELL_X1 FILLER_135_532 ();
 FILLCELL_X2 FILLER_135_554 ();
 FILLCELL_X16 FILLER_135_560 ();
 FILLCELL_X2 FILLER_135_576 ();
 FILLCELL_X1 FILLER_135_578 ();
 FILLCELL_X16 FILLER_135_594 ();
 FILLCELL_X1 FILLER_135_610 ();
 FILLCELL_X8 FILLER_135_630 ();
 FILLCELL_X4 FILLER_135_638 ();
 FILLCELL_X2 FILLER_135_656 ();
 FILLCELL_X2 FILLER_135_706 ();
 FILLCELL_X16 FILLER_135_739 ();
 FILLCELL_X4 FILLER_135_755 ();
 FILLCELL_X2 FILLER_135_759 ();
 FILLCELL_X8 FILLER_135_780 ();
 FILLCELL_X4 FILLER_135_788 ();
 FILLCELL_X1 FILLER_135_792 ();
 FILLCELL_X1 FILLER_135_805 ();
 FILLCELL_X2 FILLER_135_824 ();
 FILLCELL_X8 FILLER_135_843 ();
 FILLCELL_X4 FILLER_135_851 ();
 FILLCELL_X1 FILLER_135_855 ();
 FILLCELL_X2 FILLER_135_859 ();
 FILLCELL_X1 FILLER_135_865 ();
 FILLCELL_X1 FILLER_135_871 ();
 FILLCELL_X1 FILLER_135_881 ();
 FILLCELL_X1 FILLER_135_885 ();
 FILLCELL_X8 FILLER_135_911 ();
 FILLCELL_X2 FILLER_135_919 ();
 FILLCELL_X1 FILLER_135_921 ();
 FILLCELL_X2 FILLER_135_932 ();
 FILLCELL_X1 FILLER_135_934 ();
 FILLCELL_X8 FILLER_135_965 ();
 FILLCELL_X4 FILLER_135_973 ();
 FILLCELL_X2 FILLER_135_977 ();
 FILLCELL_X1 FILLER_135_979 ();
 FILLCELL_X2 FILLER_135_1005 ();
 FILLCELL_X8 FILLER_135_1014 ();
 FILLCELL_X8 FILLER_135_1041 ();
 FILLCELL_X4 FILLER_135_1049 ();
 FILLCELL_X2 FILLER_135_1077 ();
 FILLCELL_X8 FILLER_135_1088 ();
 FILLCELL_X4 FILLER_135_1096 ();
 FILLCELL_X2 FILLER_135_1100 ();
 FILLCELL_X1 FILLER_135_1102 ();
 FILLCELL_X32 FILLER_135_1120 ();
 FILLCELL_X16 FILLER_135_1152 ();
 FILLCELL_X4 FILLER_135_1175 ();
 FILLCELL_X2 FILLER_135_1207 ();
 FILLCELL_X1 FILLER_135_1209 ();
 FILLCELL_X8 FILLER_136_1 ();
 FILLCELL_X4 FILLER_136_9 ();
 FILLCELL_X2 FILLER_136_13 ();
 FILLCELL_X1 FILLER_136_15 ();
 FILLCELL_X8 FILLER_136_30 ();
 FILLCELL_X1 FILLER_136_38 ();
 FILLCELL_X32 FILLER_136_48 ();
 FILLCELL_X4 FILLER_136_80 ();
 FILLCELL_X2 FILLER_136_84 ();
 FILLCELL_X1 FILLER_136_86 ();
 FILLCELL_X1 FILLER_136_104 ();
 FILLCELL_X8 FILLER_136_136 ();
 FILLCELL_X4 FILLER_136_144 ();
 FILLCELL_X2 FILLER_136_148 ();
 FILLCELL_X2 FILLER_136_164 ();
 FILLCELL_X8 FILLER_136_190 ();
 FILLCELL_X2 FILLER_136_215 ();
 FILLCELL_X32 FILLER_136_241 ();
 FILLCELL_X16 FILLER_136_273 ();
 FILLCELL_X4 FILLER_136_289 ();
 FILLCELL_X2 FILLER_136_293 ();
 FILLCELL_X1 FILLER_136_295 ();
 FILLCELL_X16 FILLER_136_299 ();
 FILLCELL_X1 FILLER_136_315 ();
 FILLCELL_X8 FILLER_136_333 ();
 FILLCELL_X2 FILLER_136_341 ();
 FILLCELL_X32 FILLER_136_347 ();
 FILLCELL_X32 FILLER_136_379 ();
 FILLCELL_X4 FILLER_136_411 ();
 FILLCELL_X2 FILLER_136_415 ();
 FILLCELL_X32 FILLER_136_420 ();
 FILLCELL_X32 FILLER_136_452 ();
 FILLCELL_X1 FILLER_136_484 ();
 FILLCELL_X8 FILLER_136_489 ();
 FILLCELL_X1 FILLER_136_497 ();
 FILLCELL_X2 FILLER_136_501 ();
 FILLCELL_X4 FILLER_136_513 ();
 FILLCELL_X4 FILLER_136_526 ();
 FILLCELL_X2 FILLER_136_576 ();
 FILLCELL_X2 FILLER_136_607 ();
 FILLCELL_X8 FILLER_136_620 ();
 FILLCELL_X2 FILLER_136_628 ();
 FILLCELL_X1 FILLER_136_630 ();
 FILLCELL_X2 FILLER_136_632 ();
 FILLCELL_X1 FILLER_136_634 ();
 FILLCELL_X8 FILLER_136_669 ();
 FILLCELL_X2 FILLER_136_677 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X16 FILLER_136_728 ();
 FILLCELL_X8 FILLER_136_746 ();
 FILLCELL_X4 FILLER_136_754 ();
 FILLCELL_X2 FILLER_136_758 ();
 FILLCELL_X1 FILLER_136_760 ();
 FILLCELL_X1 FILLER_136_773 ();
 FILLCELL_X4 FILLER_136_781 ();
 FILLCELL_X2 FILLER_136_785 ();
 FILLCELL_X1 FILLER_136_787 ();
 FILLCELL_X1 FILLER_136_799 ();
 FILLCELL_X1 FILLER_136_804 ();
 FILLCELL_X2 FILLER_136_814 ();
 FILLCELL_X2 FILLER_136_835 ();
 FILLCELL_X1 FILLER_136_837 ();
 FILLCELL_X16 FILLER_136_848 ();
 FILLCELL_X8 FILLER_136_864 ();
 FILLCELL_X4 FILLER_136_872 ();
 FILLCELL_X2 FILLER_136_894 ();
 FILLCELL_X4 FILLER_136_903 ();
 FILLCELL_X2 FILLER_136_907 ();
 FILLCELL_X1 FILLER_136_909 ();
 FILLCELL_X8 FILLER_136_937 ();
 FILLCELL_X4 FILLER_136_945 ();
 FILLCELL_X2 FILLER_136_949 ();
 FILLCELL_X4 FILLER_136_959 ();
 FILLCELL_X4 FILLER_136_971 ();
 FILLCELL_X4 FILLER_136_988 ();
 FILLCELL_X8 FILLER_136_1008 ();
 FILLCELL_X1 FILLER_136_1016 ();
 FILLCELL_X8 FILLER_136_1036 ();
 FILLCELL_X2 FILLER_136_1044 ();
 FILLCELL_X8 FILLER_136_1051 ();
 FILLCELL_X1 FILLER_136_1059 ();
 FILLCELL_X1 FILLER_136_1086 ();
 FILLCELL_X1 FILLER_136_1096 ();
 FILLCELL_X1 FILLER_136_1102 ();
 FILLCELL_X16 FILLER_136_1106 ();
 FILLCELL_X8 FILLER_136_1122 ();
 FILLCELL_X4 FILLER_136_1130 ();
 FILLCELL_X2 FILLER_136_1134 ();
 FILLCELL_X8 FILLER_136_1160 ();
 FILLCELL_X4 FILLER_136_1168 ();
 FILLCELL_X2 FILLER_136_1172 ();
 FILLCELL_X1 FILLER_136_1174 ();
 FILLCELL_X8 FILLER_136_1192 ();
 FILLCELL_X8 FILLER_137_1 ();
 FILLCELL_X2 FILLER_137_9 ();
 FILLCELL_X8 FILLER_137_49 ();
 FILLCELL_X4 FILLER_137_57 ();
 FILLCELL_X2 FILLER_137_61 ();
 FILLCELL_X2 FILLER_137_70 ();
 FILLCELL_X1 FILLER_137_72 ();
 FILLCELL_X2 FILLER_137_87 ();
 FILLCELL_X4 FILLER_137_96 ();
 FILLCELL_X1 FILLER_137_100 ();
 FILLCELL_X8 FILLER_137_108 ();
 FILLCELL_X1 FILLER_137_116 ();
 FILLCELL_X16 FILLER_137_124 ();
 FILLCELL_X4 FILLER_137_140 ();
 FILLCELL_X4 FILLER_137_168 ();
 FILLCELL_X2 FILLER_137_172 ();
 FILLCELL_X16 FILLER_137_181 ();
 FILLCELL_X8 FILLER_137_197 ();
 FILLCELL_X1 FILLER_137_205 ();
 FILLCELL_X2 FILLER_137_223 ();
 FILLCELL_X1 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_240 ();
 FILLCELL_X32 FILLER_137_272 ();
 FILLCELL_X32 FILLER_137_304 ();
 FILLCELL_X32 FILLER_137_336 ();
 FILLCELL_X32 FILLER_137_368 ();
 FILLCELL_X32 FILLER_137_400 ();
 FILLCELL_X32 FILLER_137_432 ();
 FILLCELL_X16 FILLER_137_464 ();
 FILLCELL_X8 FILLER_137_480 ();
 FILLCELL_X1 FILLER_137_488 ();
 FILLCELL_X4 FILLER_137_491 ();
 FILLCELL_X1 FILLER_137_495 ();
 FILLCELL_X4 FILLER_137_523 ();
 FILLCELL_X2 FILLER_137_527 ();
 FILLCELL_X2 FILLER_137_533 ();
 FILLCELL_X1 FILLER_137_535 ();
 FILLCELL_X1 FILLER_137_572 ();
 FILLCELL_X1 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_594 ();
 FILLCELL_X16 FILLER_137_626 ();
 FILLCELL_X4 FILLER_137_642 ();
 FILLCELL_X2 FILLER_137_646 ();
 FILLCELL_X1 FILLER_137_648 ();
 FILLCELL_X16 FILLER_137_654 ();
 FILLCELL_X4 FILLER_137_670 ();
 FILLCELL_X1 FILLER_137_674 ();
 FILLCELL_X2 FILLER_137_682 ();
 FILLCELL_X8 FILLER_137_701 ();
 FILLCELL_X4 FILLER_137_709 ();
 FILLCELL_X2 FILLER_137_713 ();
 FILLCELL_X4 FILLER_137_751 ();
 FILLCELL_X1 FILLER_137_755 ();
 FILLCELL_X2 FILLER_137_776 ();
 FILLCELL_X1 FILLER_137_778 ();
 FILLCELL_X1 FILLER_137_786 ();
 FILLCELL_X2 FILLER_137_790 ();
 FILLCELL_X1 FILLER_137_792 ();
 FILLCELL_X1 FILLER_137_827 ();
 FILLCELL_X4 FILLER_137_832 ();
 FILLCELL_X1 FILLER_137_836 ();
 FILLCELL_X1 FILLER_137_842 ();
 FILLCELL_X16 FILLER_137_856 ();
 FILLCELL_X2 FILLER_137_872 ();
 FILLCELL_X1 FILLER_137_879 ();
 FILLCELL_X4 FILLER_137_893 ();
 FILLCELL_X2 FILLER_137_897 ();
 FILLCELL_X1 FILLER_137_908 ();
 FILLCELL_X8 FILLER_137_913 ();
 FILLCELL_X2 FILLER_137_921 ();
 FILLCELL_X8 FILLER_137_928 ();
 FILLCELL_X2 FILLER_137_936 ();
 FILLCELL_X1 FILLER_137_938 ();
 FILLCELL_X8 FILLER_137_941 ();
 FILLCELL_X2 FILLER_137_949 ();
 FILLCELL_X1 FILLER_137_951 ();
 FILLCELL_X8 FILLER_137_968 ();
 FILLCELL_X1 FILLER_137_976 ();
 FILLCELL_X4 FILLER_137_986 ();
 FILLCELL_X8 FILLER_137_993 ();
 FILLCELL_X4 FILLER_137_1001 ();
 FILLCELL_X8 FILLER_137_1008 ();
 FILLCELL_X4 FILLER_137_1016 ();
 FILLCELL_X2 FILLER_137_1020 ();
 FILLCELL_X1 FILLER_137_1041 ();
 FILLCELL_X2 FILLER_137_1089 ();
 FILLCELL_X16 FILLER_137_1117 ();
 FILLCELL_X1 FILLER_137_1133 ();
 FILLCELL_X16 FILLER_137_1158 ();
 FILLCELL_X4 FILLER_137_1174 ();
 FILLCELL_X1 FILLER_137_1178 ();
 FILLCELL_X4 FILLER_137_1196 ();
 FILLCELL_X1 FILLER_137_1200 ();
 FILLCELL_X2 FILLER_137_1204 ();
 FILLCELL_X1 FILLER_137_1209 ();
 FILLCELL_X8 FILLER_138_1 ();
 FILLCELL_X16 FILLER_138_12 ();
 FILLCELL_X1 FILLER_138_28 ();
 FILLCELL_X4 FILLER_138_46 ();
 FILLCELL_X2 FILLER_138_50 ();
 FILLCELL_X8 FILLER_138_76 ();
 FILLCELL_X4 FILLER_138_84 ();
 FILLCELL_X1 FILLER_138_88 ();
 FILLCELL_X4 FILLER_138_127 ();
 FILLCELL_X8 FILLER_138_138 ();
 FILLCELL_X1 FILLER_138_146 ();
 FILLCELL_X2 FILLER_138_168 ();
 FILLCELL_X1 FILLER_138_177 ();
 FILLCELL_X2 FILLER_138_185 ();
 FILLCELL_X16 FILLER_138_194 ();
 FILLCELL_X1 FILLER_138_210 ();
 FILLCELL_X1 FILLER_138_218 ();
 FILLCELL_X2 FILLER_138_230 ();
 FILLCELL_X1 FILLER_138_232 ();
 FILLCELL_X4 FILLER_138_245 ();
 FILLCELL_X1 FILLER_138_249 ();
 FILLCELL_X4 FILLER_138_264 ();
 FILLCELL_X2 FILLER_138_275 ();
 FILLCELL_X1 FILLER_138_277 ();
 FILLCELL_X32 FILLER_138_295 ();
 FILLCELL_X32 FILLER_138_327 ();
 FILLCELL_X32 FILLER_138_359 ();
 FILLCELL_X32 FILLER_138_391 ();
 FILLCELL_X32 FILLER_138_423 ();
 FILLCELL_X32 FILLER_138_455 ();
 FILLCELL_X4 FILLER_138_487 ();
 FILLCELL_X1 FILLER_138_491 ();
 FILLCELL_X32 FILLER_138_511 ();
 FILLCELL_X8 FILLER_138_543 ();
 FILLCELL_X4 FILLER_138_551 ();
 FILLCELL_X1 FILLER_138_562 ();
 FILLCELL_X1 FILLER_138_567 ();
 FILLCELL_X32 FILLER_138_587 ();
 FILLCELL_X8 FILLER_138_619 ();
 FILLCELL_X4 FILLER_138_627 ();
 FILLCELL_X8 FILLER_138_632 ();
 FILLCELL_X4 FILLER_138_640 ();
 FILLCELL_X2 FILLER_138_644 ();
 FILLCELL_X16 FILLER_138_663 ();
 FILLCELL_X2 FILLER_138_679 ();
 FILLCELL_X8 FILLER_138_703 ();
 FILLCELL_X4 FILLER_138_711 ();
 FILLCELL_X2 FILLER_138_715 ();
 FILLCELL_X32 FILLER_138_754 ();
 FILLCELL_X4 FILLER_138_786 ();
 FILLCELL_X2 FILLER_138_790 ();
 FILLCELL_X1 FILLER_138_797 ();
 FILLCELL_X2 FILLER_138_812 ();
 FILLCELL_X2 FILLER_138_819 ();
 FILLCELL_X2 FILLER_138_825 ();
 FILLCELL_X8 FILLER_138_829 ();
 FILLCELL_X1 FILLER_138_837 ();
 FILLCELL_X2 FILLER_138_865 ();
 FILLCELL_X2 FILLER_138_906 ();
 FILLCELL_X4 FILLER_138_919 ();
 FILLCELL_X2 FILLER_138_923 ();
 FILLCELL_X1 FILLER_138_925 ();
 FILLCELL_X16 FILLER_138_976 ();
 FILLCELL_X8 FILLER_138_992 ();
 FILLCELL_X4 FILLER_138_1000 ();
 FILLCELL_X2 FILLER_138_1004 ();
 FILLCELL_X1 FILLER_138_1012 ();
 FILLCELL_X2 FILLER_138_1022 ();
 FILLCELL_X1 FILLER_138_1024 ();
 FILLCELL_X16 FILLER_138_1032 ();
 FILLCELL_X8 FILLER_138_1048 ();
 FILLCELL_X4 FILLER_138_1056 ();
 FILLCELL_X2 FILLER_138_1083 ();
 FILLCELL_X4 FILLER_138_1123 ();
 FILLCELL_X2 FILLER_138_1127 ();
 FILLCELL_X8 FILLER_138_1160 ();
 FILLCELL_X4 FILLER_138_1168 ();
 FILLCELL_X2 FILLER_138_1172 ();
 FILLCELL_X8 FILLER_138_1197 ();
 FILLCELL_X2 FILLER_138_1205 ();
 FILLCELL_X1 FILLER_138_1207 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X16 FILLER_139_33 ();
 FILLCELL_X8 FILLER_139_49 ();
 FILLCELL_X2 FILLER_139_57 ();
 FILLCELL_X1 FILLER_139_59 ();
 FILLCELL_X16 FILLER_139_77 ();
 FILLCELL_X4 FILLER_139_136 ();
 FILLCELL_X2 FILLER_139_140 ();
 FILLCELL_X2 FILLER_139_159 ();
 FILLCELL_X1 FILLER_139_171 ();
 FILLCELL_X8 FILLER_139_196 ();
 FILLCELL_X1 FILLER_139_204 ();
 FILLCELL_X8 FILLER_139_212 ();
 FILLCELL_X1 FILLER_139_237 ();
 FILLCELL_X1 FILLER_139_272 ();
 FILLCELL_X32 FILLER_139_280 ();
 FILLCELL_X32 FILLER_139_312 ();
 FILLCELL_X32 FILLER_139_344 ();
 FILLCELL_X32 FILLER_139_376 ();
 FILLCELL_X32 FILLER_139_408 ();
 FILLCELL_X32 FILLER_139_440 ();
 FILLCELL_X32 FILLER_139_472 ();
 FILLCELL_X32 FILLER_139_504 ();
 FILLCELL_X4 FILLER_139_536 ();
 FILLCELL_X2 FILLER_139_540 ();
 FILLCELL_X8 FILLER_139_549 ();
 FILLCELL_X2 FILLER_139_557 ();
 FILLCELL_X1 FILLER_139_559 ();
 FILLCELL_X16 FILLER_139_594 ();
 FILLCELL_X4 FILLER_139_610 ();
 FILLCELL_X1 FILLER_139_614 ();
 FILLCELL_X2 FILLER_139_632 ();
 FILLCELL_X2 FILLER_139_641 ();
 FILLCELL_X1 FILLER_139_643 ();
 FILLCELL_X2 FILLER_139_651 ();
 FILLCELL_X1 FILLER_139_653 ();
 FILLCELL_X2 FILLER_139_661 ();
 FILLCELL_X4 FILLER_139_709 ();
 FILLCELL_X2 FILLER_139_713 ();
 FILLCELL_X1 FILLER_139_715 ();
 FILLCELL_X8 FILLER_139_751 ();
 FILLCELL_X4 FILLER_139_759 ();
 FILLCELL_X2 FILLER_139_763 ();
 FILLCELL_X4 FILLER_139_781 ();
 FILLCELL_X2 FILLER_139_790 ();
 FILLCELL_X4 FILLER_139_801 ();
 FILLCELL_X2 FILLER_139_809 ();
 FILLCELL_X1 FILLER_139_811 ();
 FILLCELL_X8 FILLER_139_816 ();
 FILLCELL_X4 FILLER_139_824 ();
 FILLCELL_X2 FILLER_139_828 ();
 FILLCELL_X1 FILLER_139_830 ();
 FILLCELL_X1 FILLER_139_844 ();
 FILLCELL_X8 FILLER_139_901 ();
 FILLCELL_X1 FILLER_139_909 ();
 FILLCELL_X1 FILLER_139_914 ();
 FILLCELL_X2 FILLER_139_940 ();
 FILLCELL_X1 FILLER_139_955 ();
 FILLCELL_X1 FILLER_139_991 ();
 FILLCELL_X4 FILLER_139_995 ();
 FILLCELL_X2 FILLER_139_999 ();
 FILLCELL_X1 FILLER_139_1011 ();
 FILLCELL_X8 FILLER_139_1040 ();
 FILLCELL_X4 FILLER_139_1051 ();
 FILLCELL_X32 FILLER_139_1059 ();
 FILLCELL_X4 FILLER_139_1091 ();
 FILLCELL_X1 FILLER_139_1095 ();
 FILLCELL_X16 FILLER_139_1120 ();
 FILLCELL_X4 FILLER_139_1145 ();
 FILLCELL_X1 FILLER_139_1149 ();
 FILLCELL_X8 FILLER_139_1167 ();
 FILLCELL_X4 FILLER_139_1199 ();
 FILLCELL_X1 FILLER_139_1213 ();
 FILLCELL_X1 FILLER_139_1217 ();
 FILLCELL_X1 FILLER_139_1230 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X16 FILLER_140_65 ();
 FILLCELL_X4 FILLER_140_81 ();
 FILLCELL_X1 FILLER_140_85 ();
 FILLCELL_X4 FILLER_140_110 ();
 FILLCELL_X2 FILLER_140_114 ();
 FILLCELL_X16 FILLER_140_123 ();
 FILLCELL_X2 FILLER_140_139 ();
 FILLCELL_X4 FILLER_140_148 ();
 FILLCELL_X1 FILLER_140_152 ();
 FILLCELL_X1 FILLER_140_175 ();
 FILLCELL_X8 FILLER_140_193 ();
 FILLCELL_X2 FILLER_140_201 ();
 FILLCELL_X1 FILLER_140_203 ();
 FILLCELL_X4 FILLER_140_221 ();
 FILLCELL_X1 FILLER_140_225 ();
 FILLCELL_X4 FILLER_140_233 ();
 FILLCELL_X2 FILLER_140_237 ();
 FILLCELL_X1 FILLER_140_239 ();
 FILLCELL_X2 FILLER_140_242 ();
 FILLCELL_X32 FILLER_140_275 ();
 FILLCELL_X32 FILLER_140_307 ();
 FILLCELL_X32 FILLER_140_339 ();
 FILLCELL_X32 FILLER_140_371 ();
 FILLCELL_X2 FILLER_140_403 ();
 FILLCELL_X32 FILLER_140_418 ();
 FILLCELL_X32 FILLER_140_450 ();
 FILLCELL_X8 FILLER_140_482 ();
 FILLCELL_X4 FILLER_140_490 ();
 FILLCELL_X1 FILLER_140_494 ();
 FILLCELL_X32 FILLER_140_498 ();
 FILLCELL_X32 FILLER_140_530 ();
 FILLCELL_X32 FILLER_140_562 ();
 FILLCELL_X32 FILLER_140_594 ();
 FILLCELL_X4 FILLER_140_626 ();
 FILLCELL_X1 FILLER_140_630 ();
 FILLCELL_X4 FILLER_140_632 ();
 FILLCELL_X2 FILLER_140_636 ();
 FILLCELL_X1 FILLER_140_638 ();
 FILLCELL_X2 FILLER_140_646 ();
 FILLCELL_X1 FILLER_140_648 ();
 FILLCELL_X4 FILLER_140_673 ();
 FILLCELL_X16 FILLER_140_711 ();
 FILLCELL_X4 FILLER_140_727 ();
 FILLCELL_X2 FILLER_140_731 ();
 FILLCELL_X1 FILLER_140_733 ();
 FILLCELL_X16 FILLER_140_737 ();
 FILLCELL_X8 FILLER_140_753 ();
 FILLCELL_X4 FILLER_140_761 ();
 FILLCELL_X2 FILLER_140_765 ();
 FILLCELL_X2 FILLER_140_770 ();
 FILLCELL_X1 FILLER_140_772 ();
 FILLCELL_X8 FILLER_140_777 ();
 FILLCELL_X2 FILLER_140_785 ();
 FILLCELL_X1 FILLER_140_787 ();
 FILLCELL_X8 FILLER_140_814 ();
 FILLCELL_X2 FILLER_140_822 ();
 FILLCELL_X1 FILLER_140_855 ();
 FILLCELL_X1 FILLER_140_864 ();
 FILLCELL_X2 FILLER_140_903 ();
 FILLCELL_X4 FILLER_140_910 ();
 FILLCELL_X2 FILLER_140_917 ();
 FILLCELL_X2 FILLER_140_926 ();
 FILLCELL_X2 FILLER_140_933 ();
 FILLCELL_X1 FILLER_140_935 ();
 FILLCELL_X1 FILLER_140_942 ();
 FILLCELL_X1 FILLER_140_945 ();
 FILLCELL_X2 FILLER_140_975 ();
 FILLCELL_X8 FILLER_140_980 ();
 FILLCELL_X2 FILLER_140_988 ();
 FILLCELL_X8 FILLER_140_1014 ();
 FILLCELL_X1 FILLER_140_1022 ();
 FILLCELL_X8 FILLER_140_1027 ();
 FILLCELL_X4 FILLER_140_1035 ();
 FILLCELL_X2 FILLER_140_1039 ();
 FILLCELL_X8 FILLER_140_1062 ();
 FILLCELL_X1 FILLER_140_1070 ();
 FILLCELL_X4 FILLER_140_1074 ();
 FILLCELL_X2 FILLER_140_1102 ();
 FILLCELL_X32 FILLER_140_1121 ();
 FILLCELL_X2 FILLER_140_1153 ();
 FILLCELL_X1 FILLER_140_1155 ();
 FILLCELL_X8 FILLER_140_1173 ();
 FILLCELL_X2 FILLER_140_1227 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X16 FILLER_141_65 ();
 FILLCELL_X8 FILLER_141_81 ();
 FILLCELL_X16 FILLER_141_130 ();
 FILLCELL_X8 FILLER_141_146 ();
 FILLCELL_X4 FILLER_141_154 ();
 FILLCELL_X2 FILLER_141_158 ();
 FILLCELL_X1 FILLER_141_160 ();
 FILLCELL_X32 FILLER_141_168 ();
 FILLCELL_X8 FILLER_141_200 ();
 FILLCELL_X2 FILLER_141_208 ();
 FILLCELL_X1 FILLER_141_210 ();
 FILLCELL_X32 FILLER_141_235 ();
 FILLCELL_X32 FILLER_141_267 ();
 FILLCELL_X32 FILLER_141_299 ();
 FILLCELL_X32 FILLER_141_331 ();
 FILLCELL_X32 FILLER_141_363 ();
 FILLCELL_X32 FILLER_141_395 ();
 FILLCELL_X32 FILLER_141_427 ();
 FILLCELL_X32 FILLER_141_459 ();
 FILLCELL_X32 FILLER_141_491 ();
 FILLCELL_X32 FILLER_141_523 ();
 FILLCELL_X32 FILLER_141_555 ();
 FILLCELL_X32 FILLER_141_587 ();
 FILLCELL_X8 FILLER_141_619 ();
 FILLCELL_X4 FILLER_141_627 ();
 FILLCELL_X2 FILLER_141_631 ();
 FILLCELL_X1 FILLER_141_633 ();
 FILLCELL_X8 FILLER_141_658 ();
 FILLCELL_X4 FILLER_141_666 ();
 FILLCELL_X32 FILLER_141_711 ();
 FILLCELL_X4 FILLER_141_743 ();
 FILLCELL_X2 FILLER_141_747 ();
 FILLCELL_X8 FILLER_141_752 ();
 FILLCELL_X4 FILLER_141_760 ();
 FILLCELL_X4 FILLER_141_781 ();
 FILLCELL_X2 FILLER_141_804 ();
 FILLCELL_X1 FILLER_141_806 ();
 FILLCELL_X16 FILLER_141_814 ();
 FILLCELL_X1 FILLER_141_830 ();
 FILLCELL_X2 FILLER_141_833 ();
 FILLCELL_X1 FILLER_141_835 ();
 FILLCELL_X1 FILLER_141_848 ();
 FILLCELL_X1 FILLER_141_857 ();
 FILLCELL_X8 FILLER_141_922 ();
 FILLCELL_X8 FILLER_141_947 ();
 FILLCELL_X2 FILLER_141_955 ();
 FILLCELL_X1 FILLER_141_960 ();
 FILLCELL_X4 FILLER_141_964 ();
 FILLCELL_X2 FILLER_141_968 ();
 FILLCELL_X1 FILLER_141_970 ();
 FILLCELL_X1 FILLER_141_985 ();
 FILLCELL_X2 FILLER_141_993 ();
 FILLCELL_X1 FILLER_141_995 ();
 FILLCELL_X1 FILLER_141_1013 ();
 FILLCELL_X4 FILLER_141_1060 ();
 FILLCELL_X2 FILLER_141_1064 ();
 FILLCELL_X1 FILLER_141_1066 ();
 FILLCELL_X1 FILLER_141_1084 ();
 FILLCELL_X2 FILLER_141_1089 ();
 FILLCELL_X1 FILLER_141_1091 ();
 FILLCELL_X16 FILLER_141_1113 ();
 FILLCELL_X4 FILLER_141_1129 ();
 FILLCELL_X2 FILLER_141_1133 ();
 FILLCELL_X1 FILLER_141_1135 ();
 FILLCELL_X2 FILLER_141_1160 ();
 FILLCELL_X1 FILLER_141_1162 ();
 FILLCELL_X4 FILLER_141_1168 ();
 FILLCELL_X2 FILLER_141_1238 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X8 FILLER_142_97 ();
 FILLCELL_X4 FILLER_142_105 ();
 FILLCELL_X2 FILLER_142_109 ();
 FILLCELL_X8 FILLER_142_118 ();
 FILLCELL_X4 FILLER_142_126 ();
 FILLCELL_X16 FILLER_142_137 ();
 FILLCELL_X32 FILLER_142_192 ();
 FILLCELL_X16 FILLER_142_224 ();
 FILLCELL_X8 FILLER_142_240 ();
 FILLCELL_X1 FILLER_142_248 ();
 FILLCELL_X32 FILLER_142_252 ();
 FILLCELL_X32 FILLER_142_284 ();
 FILLCELL_X32 FILLER_142_316 ();
 FILLCELL_X32 FILLER_142_348 ();
 FILLCELL_X32 FILLER_142_380 ();
 FILLCELL_X8 FILLER_142_412 ();
 FILLCELL_X1 FILLER_142_420 ();
 FILLCELL_X32 FILLER_142_426 ();
 FILLCELL_X32 FILLER_142_458 ();
 FILLCELL_X32 FILLER_142_490 ();
 FILLCELL_X32 FILLER_142_522 ();
 FILLCELL_X32 FILLER_142_554 ();
 FILLCELL_X32 FILLER_142_586 ();
 FILLCELL_X8 FILLER_142_618 ();
 FILLCELL_X4 FILLER_142_626 ();
 FILLCELL_X1 FILLER_142_630 ();
 FILLCELL_X16 FILLER_142_639 ();
 FILLCELL_X8 FILLER_142_655 ();
 FILLCELL_X2 FILLER_142_663 ();
 FILLCELL_X2 FILLER_142_672 ();
 FILLCELL_X4 FILLER_142_681 ();
 FILLCELL_X4 FILLER_142_692 ();
 FILLCELL_X4 FILLER_142_703 ();
 FILLCELL_X16 FILLER_142_716 ();
 FILLCELL_X8 FILLER_142_732 ();
 FILLCELL_X4 FILLER_142_740 ();
 FILLCELL_X1 FILLER_142_744 ();
 FILLCELL_X2 FILLER_142_755 ();
 FILLCELL_X2 FILLER_142_762 ();
 FILLCELL_X1 FILLER_142_764 ();
 FILLCELL_X1 FILLER_142_772 ();
 FILLCELL_X8 FILLER_142_780 ();
 FILLCELL_X4 FILLER_142_788 ();
 FILLCELL_X2 FILLER_142_806 ();
 FILLCELL_X2 FILLER_142_817 ();
 FILLCELL_X8 FILLER_142_836 ();
 FILLCELL_X1 FILLER_142_870 ();
 FILLCELL_X1 FILLER_142_885 ();
 FILLCELL_X2 FILLER_142_893 ();
 FILLCELL_X1 FILLER_142_895 ();
 FILLCELL_X2 FILLER_142_918 ();
 FILLCELL_X1 FILLER_142_920 ();
 FILLCELL_X2 FILLER_142_926 ();
 FILLCELL_X1 FILLER_142_928 ();
 FILLCELL_X16 FILLER_142_932 ();
 FILLCELL_X8 FILLER_142_997 ();
 FILLCELL_X4 FILLER_142_1005 ();
 FILLCELL_X1 FILLER_142_1009 ();
 FILLCELL_X1 FILLER_142_1020 ();
 FILLCELL_X1 FILLER_142_1033 ();
 FILLCELL_X2 FILLER_142_1043 ();
 FILLCELL_X1 FILLER_142_1061 ();
 FILLCELL_X32 FILLER_142_1065 ();
 FILLCELL_X8 FILLER_142_1097 ();
 FILLCELL_X1 FILLER_142_1105 ();
 FILLCELL_X16 FILLER_142_1122 ();
 FILLCELL_X8 FILLER_142_1138 ();
 FILLCELL_X4 FILLER_142_1146 ();
 FILLCELL_X2 FILLER_142_1150 ();
 FILLCELL_X16 FILLER_142_1159 ();
 FILLCELL_X8 FILLER_142_1175 ();
 FILLCELL_X2 FILLER_142_1214 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X16 FILLER_143_33 ();
 FILLCELL_X8 FILLER_143_49 ();
 FILLCELL_X4 FILLER_143_57 ();
 FILLCELL_X32 FILLER_143_64 ();
 FILLCELL_X16 FILLER_143_96 ();
 FILLCELL_X2 FILLER_143_112 ();
 FILLCELL_X32 FILLER_143_138 ();
 FILLCELL_X4 FILLER_143_170 ();
 FILLCELL_X2 FILLER_143_174 ();
 FILLCELL_X32 FILLER_143_183 ();
 FILLCELL_X32 FILLER_143_215 ();
 FILLCELL_X32 FILLER_143_247 ();
 FILLCELL_X32 FILLER_143_279 ();
 FILLCELL_X32 FILLER_143_311 ();
 FILLCELL_X32 FILLER_143_343 ();
 FILLCELL_X32 FILLER_143_375 ();
 FILLCELL_X32 FILLER_143_407 ();
 FILLCELL_X16 FILLER_143_439 ();
 FILLCELL_X8 FILLER_143_455 ();
 FILLCELL_X2 FILLER_143_463 ();
 FILLCELL_X1 FILLER_143_465 ();
 FILLCELL_X32 FILLER_143_483 ();
 FILLCELL_X32 FILLER_143_515 ();
 FILLCELL_X32 FILLER_143_547 ();
 FILLCELL_X32 FILLER_143_579 ();
 FILLCELL_X8 FILLER_143_611 ();
 FILLCELL_X4 FILLER_143_619 ();
 FILLCELL_X1 FILLER_143_630 ();
 FILLCELL_X1 FILLER_143_648 ();
 FILLCELL_X1 FILLER_143_656 ();
 FILLCELL_X32 FILLER_143_666 ();
 FILLCELL_X16 FILLER_143_698 ();
 FILLCELL_X8 FILLER_143_714 ();
 FILLCELL_X4 FILLER_143_722 ();
 FILLCELL_X2 FILLER_143_726 ();
 FILLCELL_X8 FILLER_143_733 ();
 FILLCELL_X4 FILLER_143_741 ();
 FILLCELL_X1 FILLER_143_745 ();
 FILLCELL_X1 FILLER_143_752 ();
 FILLCELL_X2 FILLER_143_760 ();
 FILLCELL_X32 FILLER_143_774 ();
 FILLCELL_X8 FILLER_143_806 ();
 FILLCELL_X1 FILLER_143_814 ();
 FILLCELL_X8 FILLER_143_818 ();
 FILLCELL_X4 FILLER_143_826 ();
 FILLCELL_X2 FILLER_143_830 ();
 FILLCELL_X1 FILLER_143_832 ();
 FILLCELL_X1 FILLER_143_840 ();
 FILLCELL_X1 FILLER_143_846 ();
 FILLCELL_X8 FILLER_143_852 ();
 FILLCELL_X4 FILLER_143_860 ();
 FILLCELL_X4 FILLER_143_868 ();
 FILLCELL_X2 FILLER_143_872 ();
 FILLCELL_X2 FILLER_143_877 ();
 FILLCELL_X4 FILLER_143_890 ();
 FILLCELL_X2 FILLER_143_894 ();
 FILLCELL_X2 FILLER_143_916 ();
 FILLCELL_X1 FILLER_143_918 ();
 FILLCELL_X8 FILLER_143_940 ();
 FILLCELL_X2 FILLER_143_951 ();
 FILLCELL_X32 FILLER_143_964 ();
 FILLCELL_X8 FILLER_143_996 ();
 FILLCELL_X4 FILLER_143_1004 ();
 FILLCELL_X2 FILLER_143_1008 ();
 FILLCELL_X16 FILLER_143_1023 ();
 FILLCELL_X1 FILLER_143_1039 ();
 FILLCELL_X4 FILLER_143_1046 ();
 FILLCELL_X4 FILLER_143_1054 ();
 FILLCELL_X32 FILLER_143_1064 ();
 FILLCELL_X4 FILLER_143_1096 ();
 FILLCELL_X8 FILLER_143_1121 ();
 FILLCELL_X4 FILLER_143_1129 ();
 FILLCELL_X1 FILLER_143_1133 ();
 FILLCELL_X4 FILLER_143_1167 ();
 FILLCELL_X2 FILLER_143_1207 ();
 FILLCELL_X2 FILLER_143_1235 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X16 FILLER_144_97 ();
 FILLCELL_X4 FILLER_144_113 ();
 FILLCELL_X2 FILLER_144_117 ();
 FILLCELL_X1 FILLER_144_119 ();
 FILLCELL_X32 FILLER_144_123 ();
 FILLCELL_X16 FILLER_144_155 ();
 FILLCELL_X4 FILLER_144_171 ();
 FILLCELL_X2 FILLER_144_175 ();
 FILLCELL_X1 FILLER_144_177 ();
 FILLCELL_X32 FILLER_144_195 ();
 FILLCELL_X32 FILLER_144_227 ();
 FILLCELL_X32 FILLER_144_259 ();
 FILLCELL_X32 FILLER_144_291 ();
 FILLCELL_X32 FILLER_144_323 ();
 FILLCELL_X32 FILLER_144_355 ();
 FILLCELL_X32 FILLER_144_387 ();
 FILLCELL_X32 FILLER_144_419 ();
 FILLCELL_X32 FILLER_144_451 ();
 FILLCELL_X32 FILLER_144_483 ();
 FILLCELL_X32 FILLER_144_515 ();
 FILLCELL_X32 FILLER_144_547 ();
 FILLCELL_X32 FILLER_144_579 ();
 FILLCELL_X2 FILLER_144_611 ();
 FILLCELL_X1 FILLER_144_613 ();
 FILLCELL_X4 FILLER_144_632 ();
 FILLCELL_X1 FILLER_144_636 ();
 FILLCELL_X8 FILLER_144_654 ();
 FILLCELL_X4 FILLER_144_662 ();
 FILLCELL_X2 FILLER_144_666 ();
 FILLCELL_X1 FILLER_144_668 ();
 FILLCELL_X4 FILLER_144_674 ();
 FILLCELL_X1 FILLER_144_678 ();
 FILLCELL_X4 FILLER_144_696 ();
 FILLCELL_X2 FILLER_144_700 ();
 FILLCELL_X8 FILLER_144_719 ();
 FILLCELL_X4 FILLER_144_727 ();
 FILLCELL_X1 FILLER_144_777 ();
 FILLCELL_X16 FILLER_144_781 ();
 FILLCELL_X2 FILLER_144_797 ();
 FILLCELL_X1 FILLER_144_799 ();
 FILLCELL_X1 FILLER_144_809 ();
 FILLCELL_X1 FILLER_144_836 ();
 FILLCELL_X4 FILLER_144_840 ();
 FILLCELL_X2 FILLER_144_844 ();
 FILLCELL_X4 FILLER_144_849 ();
 FILLCELL_X1 FILLER_144_871 ();
 FILLCELL_X2 FILLER_144_886 ();
 FILLCELL_X2 FILLER_144_893 ();
 FILLCELL_X2 FILLER_144_899 ();
 FILLCELL_X1 FILLER_144_910 ();
 FILLCELL_X1 FILLER_144_940 ();
 FILLCELL_X2 FILLER_144_944 ();
 FILLCELL_X1 FILLER_144_946 ();
 FILLCELL_X2 FILLER_144_957 ();
 FILLCELL_X2 FILLER_144_974 ();
 FILLCELL_X8 FILLER_144_983 ();
 FILLCELL_X4 FILLER_144_991 ();
 FILLCELL_X1 FILLER_144_995 ();
 FILLCELL_X4 FILLER_144_1000 ();
 FILLCELL_X2 FILLER_144_1004 ();
 FILLCELL_X4 FILLER_144_1013 ();
 FILLCELL_X2 FILLER_144_1017 ();
 FILLCELL_X1 FILLER_144_1019 ();
 FILLCELL_X16 FILLER_144_1052 ();
 FILLCELL_X8 FILLER_144_1068 ();
 FILLCELL_X4 FILLER_144_1076 ();
 FILLCELL_X2 FILLER_144_1080 ();
 FILLCELL_X16 FILLER_144_1104 ();
 FILLCELL_X2 FILLER_144_1120 ();
 FILLCELL_X8 FILLER_144_1129 ();
 FILLCELL_X2 FILLER_144_1137 ();
 FILLCELL_X8 FILLER_144_1163 ();
 FILLCELL_X4 FILLER_144_1171 ();
 FILLCELL_X2 FILLER_144_1175 ();
 FILLCELL_X1 FILLER_144_1201 ();
 FILLCELL_X1 FILLER_144_1209 ();
 FILLCELL_X1 FILLER_144_1217 ();
 FILLCELL_X1 FILLER_144_1234 ();
 FILLCELL_X2 FILLER_144_1238 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X4 FILLER_145_609 ();
 FILLCELL_X1 FILLER_145_613 ();
 FILLCELL_X16 FILLER_145_652 ();
 FILLCELL_X1 FILLER_145_692 ();
 FILLCELL_X4 FILLER_145_722 ();
 FILLCELL_X2 FILLER_145_726 ();
 FILLCELL_X1 FILLER_145_728 ();
 FILLCELL_X2 FILLER_145_756 ();
 FILLCELL_X4 FILLER_145_764 ();
 FILLCELL_X2 FILLER_145_776 ();
 FILLCELL_X16 FILLER_145_805 ();
 FILLCELL_X8 FILLER_145_821 ();
 FILLCELL_X2 FILLER_145_829 ();
 FILLCELL_X4 FILLER_145_838 ();
 FILLCELL_X1 FILLER_145_842 ();
 FILLCELL_X2 FILLER_145_851 ();
 FILLCELL_X2 FILLER_145_871 ();
 FILLCELL_X4 FILLER_145_880 ();
 FILLCELL_X4 FILLER_145_891 ();
 FILLCELL_X2 FILLER_145_895 ();
 FILLCELL_X1 FILLER_145_904 ();
 FILLCELL_X8 FILLER_145_908 ();
 FILLCELL_X1 FILLER_145_925 ();
 FILLCELL_X2 FILLER_145_933 ();
 FILLCELL_X2 FILLER_145_972 ();
 FILLCELL_X8 FILLER_145_981 ();
 FILLCELL_X4 FILLER_145_989 ();
 FILLCELL_X2 FILLER_145_993 ();
 FILLCELL_X2 FILLER_145_1008 ();
 FILLCELL_X1 FILLER_145_1010 ();
 FILLCELL_X2 FILLER_145_1037 ();
 FILLCELL_X16 FILLER_145_1048 ();
 FILLCELL_X8 FILLER_145_1064 ();
 FILLCELL_X4 FILLER_145_1072 ();
 FILLCELL_X2 FILLER_145_1076 ();
 FILLCELL_X4 FILLER_145_1091 ();
 FILLCELL_X1 FILLER_145_1095 ();
 FILLCELL_X32 FILLER_145_1113 ();
 FILLCELL_X8 FILLER_145_1145 ();
 FILLCELL_X16 FILLER_145_1167 ();
 FILLCELL_X2 FILLER_145_1183 ();
 FILLCELL_X2 FILLER_145_1192 ();
 FILLCELL_X1 FILLER_145_1194 ();
 FILLCELL_X16 FILLER_145_1198 ();
 FILLCELL_X2 FILLER_145_1214 ();
 FILLCELL_X1 FILLER_145_1216 ();
 FILLCELL_X2 FILLER_145_1229 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X16 FILLER_146_225 ();
 FILLCELL_X8 FILLER_146_241 ();
 FILLCELL_X2 FILLER_146_249 ();
 FILLCELL_X1 FILLER_146_251 ();
 FILLCELL_X32 FILLER_146_256 ();
 FILLCELL_X32 FILLER_146_288 ();
 FILLCELL_X32 FILLER_146_320 ();
 FILLCELL_X32 FILLER_146_352 ();
 FILLCELL_X32 FILLER_146_384 ();
 FILLCELL_X32 FILLER_146_416 ();
 FILLCELL_X32 FILLER_146_448 ();
 FILLCELL_X32 FILLER_146_480 ();
 FILLCELL_X32 FILLER_146_512 ();
 FILLCELL_X32 FILLER_146_544 ();
 FILLCELL_X32 FILLER_146_576 ();
 FILLCELL_X16 FILLER_146_608 ();
 FILLCELL_X4 FILLER_146_624 ();
 FILLCELL_X2 FILLER_146_628 ();
 FILLCELL_X1 FILLER_146_630 ();
 FILLCELL_X2 FILLER_146_632 ();
 FILLCELL_X1 FILLER_146_634 ();
 FILLCELL_X2 FILLER_146_649 ();
 FILLCELL_X16 FILLER_146_658 ();
 FILLCELL_X1 FILLER_146_674 ();
 FILLCELL_X2 FILLER_146_682 ();
 FILLCELL_X1 FILLER_146_684 ();
 FILLCELL_X8 FILLER_146_692 ();
 FILLCELL_X1 FILLER_146_700 ();
 FILLCELL_X2 FILLER_146_724 ();
 FILLCELL_X1 FILLER_146_726 ();
 FILLCELL_X2 FILLER_146_747 ();
 FILLCELL_X16 FILLER_146_756 ();
 FILLCELL_X2 FILLER_146_781 ();
 FILLCELL_X1 FILLER_146_783 ();
 FILLCELL_X4 FILLER_146_801 ();
 FILLCELL_X1 FILLER_146_805 ();
 FILLCELL_X8 FILLER_146_820 ();
 FILLCELL_X16 FILLER_146_835 ();
 FILLCELL_X1 FILLER_146_851 ();
 FILLCELL_X8 FILLER_146_863 ();
 FILLCELL_X2 FILLER_146_881 ();
 FILLCELL_X8 FILLER_146_888 ();
 FILLCELL_X2 FILLER_146_896 ();
 FILLCELL_X1 FILLER_146_898 ();
 FILLCELL_X1 FILLER_146_931 ();
 FILLCELL_X2 FILLER_146_936 ();
 FILLCELL_X2 FILLER_146_947 ();
 FILLCELL_X2 FILLER_146_971 ();
 FILLCELL_X8 FILLER_146_980 ();
 FILLCELL_X4 FILLER_146_988 ();
 FILLCELL_X4 FILLER_146_1010 ();
 FILLCELL_X2 FILLER_146_1014 ();
 FILLCELL_X1 FILLER_146_1016 ();
 FILLCELL_X4 FILLER_146_1027 ();
 FILLCELL_X2 FILLER_146_1031 ();
 FILLCELL_X2 FILLER_146_1041 ();
 FILLCELL_X8 FILLER_146_1057 ();
 FILLCELL_X4 FILLER_146_1065 ();
 FILLCELL_X2 FILLER_146_1069 ();
 FILLCELL_X1 FILLER_146_1071 ();
 FILLCELL_X2 FILLER_146_1075 ();
 FILLCELL_X2 FILLER_146_1109 ();
 FILLCELL_X16 FILLER_146_1122 ();
 FILLCELL_X4 FILLER_146_1138 ();
 FILLCELL_X2 FILLER_146_1142 ();
 FILLCELL_X1 FILLER_146_1144 ();
 FILLCELL_X16 FILLER_146_1162 ();
 FILLCELL_X4 FILLER_146_1178 ();
 FILLCELL_X2 FILLER_146_1182 ();
 FILLCELL_X2 FILLER_146_1201 ();
 FILLCELL_X1 FILLER_146_1203 ();
 FILLCELL_X16 FILLER_146_1207 ();
 FILLCELL_X8 FILLER_146_1226 ();
 FILLCELL_X4 FILLER_146_1234 ();
 FILLCELL_X2 FILLER_146_1238 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X16 FILLER_147_673 ();
 FILLCELL_X4 FILLER_147_689 ();
 FILLCELL_X2 FILLER_147_693 ();
 FILLCELL_X32 FILLER_147_700 ();
 FILLCELL_X8 FILLER_147_732 ();
 FILLCELL_X2 FILLER_147_740 ();
 FILLCELL_X2 FILLER_147_746 ();
 FILLCELL_X4 FILLER_147_759 ();
 FILLCELL_X4 FILLER_147_795 ();
 FILLCELL_X2 FILLER_147_799 ();
 FILLCELL_X4 FILLER_147_808 ();
 FILLCELL_X2 FILLER_147_812 ();
 FILLCELL_X1 FILLER_147_814 ();
 FILLCELL_X2 FILLER_147_832 ();
 FILLCELL_X2 FILLER_147_838 ();
 FILLCELL_X1 FILLER_147_840 ();
 FILLCELL_X1 FILLER_147_845 ();
 FILLCELL_X2 FILLER_147_850 ();
 FILLCELL_X1 FILLER_147_852 ();
 FILLCELL_X1 FILLER_147_865 ();
 FILLCELL_X1 FILLER_147_869 ();
 FILLCELL_X4 FILLER_147_889 ();
 FILLCELL_X2 FILLER_147_893 ();
 FILLCELL_X1 FILLER_147_895 ();
 FILLCELL_X4 FILLER_147_901 ();
 FILLCELL_X4 FILLER_147_908 ();
 FILLCELL_X4 FILLER_147_916 ();
 FILLCELL_X1 FILLER_147_920 ();
 FILLCELL_X2 FILLER_147_923 ();
 FILLCELL_X1 FILLER_147_925 ();
 FILLCELL_X1 FILLER_147_930 ();
 FILLCELL_X1 FILLER_147_937 ();
 FILLCELL_X1 FILLER_147_941 ();
 FILLCELL_X1 FILLER_147_945 ();
 FILLCELL_X1 FILLER_147_948 ();
 FILLCELL_X1 FILLER_147_967 ();
 FILLCELL_X1 FILLER_147_973 ();
 FILLCELL_X2 FILLER_147_992 ();
 FILLCELL_X2 FILLER_147_1043 ();
 FILLCELL_X1 FILLER_147_1045 ();
 FILLCELL_X8 FILLER_147_1050 ();
 FILLCELL_X2 FILLER_147_1058 ();
 FILLCELL_X4 FILLER_147_1065 ();
 FILLCELL_X1 FILLER_147_1069 ();
 FILLCELL_X1 FILLER_147_1108 ();
 FILLCELL_X32 FILLER_147_1126 ();
 FILLCELL_X32 FILLER_147_1158 ();
 FILLCELL_X8 FILLER_147_1190 ();
 FILLCELL_X4 FILLER_147_1198 ();
 FILLCELL_X2 FILLER_147_1202 ();
 FILLCELL_X8 FILLER_147_1207 ();
 FILLCELL_X2 FILLER_147_1215 ();
 FILLCELL_X1 FILLER_147_1217 ();
 FILLCELL_X4 FILLER_147_1221 ();
 FILLCELL_X1 FILLER_147_1225 ();
 FILLCELL_X8 FILLER_147_1232 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X1 FILLER_148_646 ();
 FILLCELL_X4 FILLER_148_654 ();
 FILLCELL_X2 FILLER_148_658 ();
 FILLCELL_X1 FILLER_148_660 ();
 FILLCELL_X1 FILLER_148_705 ();
 FILLCELL_X8 FILLER_148_723 ();
 FILLCELL_X1 FILLER_148_731 ();
 FILLCELL_X4 FILLER_148_749 ();
 FILLCELL_X2 FILLER_148_753 ();
 FILLCELL_X1 FILLER_148_759 ();
 FILLCELL_X1 FILLER_148_764 ();
 FILLCELL_X1 FILLER_148_777 ();
 FILLCELL_X1 FILLER_148_783 ();
 FILLCELL_X4 FILLER_148_798 ();
 FILLCELL_X8 FILLER_148_805 ();
 FILLCELL_X2 FILLER_148_813 ();
 FILLCELL_X4 FILLER_148_820 ();
 FILLCELL_X1 FILLER_148_824 ();
 FILLCELL_X1 FILLER_148_846 ();
 FILLCELL_X2 FILLER_148_857 ();
 FILLCELL_X1 FILLER_148_878 ();
 FILLCELL_X1 FILLER_148_882 ();
 FILLCELL_X8 FILLER_148_894 ();
 FILLCELL_X4 FILLER_148_902 ();
 FILLCELL_X4 FILLER_148_920 ();
 FILLCELL_X1 FILLER_148_924 ();
 FILLCELL_X4 FILLER_148_941 ();
 FILLCELL_X2 FILLER_148_945 ();
 FILLCELL_X1 FILLER_148_953 ();
 FILLCELL_X2 FILLER_148_966 ();
 FILLCELL_X1 FILLER_148_968 ();
 FILLCELL_X4 FILLER_148_977 ();
 FILLCELL_X4 FILLER_148_999 ();
 FILLCELL_X2 FILLER_148_1003 ();
 FILLCELL_X1 FILLER_148_1005 ();
 FILLCELL_X4 FILLER_148_1020 ();
 FILLCELL_X2 FILLER_148_1024 ();
 FILLCELL_X1 FILLER_148_1029 ();
 FILLCELL_X2 FILLER_148_1034 ();
 FILLCELL_X1 FILLER_148_1036 ();
 FILLCELL_X2 FILLER_148_1043 ();
 FILLCELL_X16 FILLER_148_1065 ();
 FILLCELL_X4 FILLER_148_1081 ();
 FILLCELL_X2 FILLER_148_1085 ();
 FILLCELL_X1 FILLER_148_1087 ();
 FILLCELL_X32 FILLER_148_1091 ();
 FILLCELL_X16 FILLER_148_1123 ();
 FILLCELL_X4 FILLER_148_1139 ();
 FILLCELL_X2 FILLER_148_1143 ();
 FILLCELL_X1 FILLER_148_1145 ();
 FILLCELL_X32 FILLER_148_1153 ();
 FILLCELL_X16 FILLER_148_1185 ();
 FILLCELL_X8 FILLER_148_1201 ();
 FILLCELL_X4 FILLER_148_1209 ();
 FILLCELL_X4 FILLER_148_1216 ();
 FILLCELL_X2 FILLER_148_1220 ();
 FILLCELL_X8 FILLER_148_1225 ();
 FILLCELL_X4 FILLER_148_1233 ();
 FILLCELL_X2 FILLER_148_1237 ();
 FILLCELL_X1 FILLER_148_1239 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X16 FILLER_149_609 ();
 FILLCELL_X4 FILLER_149_625 ();
 FILLCELL_X1 FILLER_149_629 ();
 FILLCELL_X2 FILLER_149_647 ();
 FILLCELL_X1 FILLER_149_649 ();
 FILLCELL_X4 FILLER_149_676 ();
 FILLCELL_X2 FILLER_149_680 ();
 FILLCELL_X2 FILLER_149_706 ();
 FILLCELL_X2 FILLER_149_715 ();
 FILLCELL_X1 FILLER_149_717 ();
 FILLCELL_X8 FILLER_149_734 ();
 FILLCELL_X4 FILLER_149_742 ();
 FILLCELL_X2 FILLER_149_762 ();
 FILLCELL_X2 FILLER_149_771 ();
 FILLCELL_X1 FILLER_149_773 ();
 FILLCELL_X2 FILLER_149_781 ();
 FILLCELL_X1 FILLER_149_783 ();
 FILLCELL_X8 FILLER_149_793 ();
 FILLCELL_X4 FILLER_149_801 ();
 FILLCELL_X2 FILLER_149_805 ();
 FILLCELL_X8 FILLER_149_831 ();
 FILLCELL_X4 FILLER_149_839 ();
 FILLCELL_X1 FILLER_149_865 ();
 FILLCELL_X1 FILLER_149_878 ();
 FILLCELL_X1 FILLER_149_883 ();
 FILLCELL_X2 FILLER_149_893 ();
 FILLCELL_X16 FILLER_149_899 ();
 FILLCELL_X4 FILLER_149_915 ();
 FILLCELL_X1 FILLER_149_919 ();
 FILLCELL_X8 FILLER_149_939 ();
 FILLCELL_X4 FILLER_149_947 ();
 FILLCELL_X1 FILLER_149_956 ();
 FILLCELL_X8 FILLER_149_961 ();
 FILLCELL_X4 FILLER_149_969 ();
 FILLCELL_X32 FILLER_149_1030 ();
 FILLCELL_X16 FILLER_149_1062 ();
 FILLCELL_X8 FILLER_149_1078 ();
 FILLCELL_X4 FILLER_149_1086 ();
 FILLCELL_X1 FILLER_149_1090 ();
 FILLCELL_X32 FILLER_149_1101 ();
 FILLCELL_X32 FILLER_149_1133 ();
 FILLCELL_X32 FILLER_149_1165 ();
 FILLCELL_X8 FILLER_149_1197 ();
 FILLCELL_X4 FILLER_149_1205 ();
 FILLCELL_X2 FILLER_149_1209 ();
 FILLCELL_X1 FILLER_149_1211 ();
 FILLCELL_X8 FILLER_149_1219 ();
 FILLCELL_X2 FILLER_149_1227 ();
 FILLCELL_X4 FILLER_149_1233 ();
 FILLCELL_X2 FILLER_149_1237 ();
 FILLCELL_X1 FILLER_149_1239 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X4 FILLER_150_609 ();
 FILLCELL_X1 FILLER_150_613 ();
 FILLCELL_X1 FILLER_150_632 ();
 FILLCELL_X1 FILLER_150_640 ();
 FILLCELL_X8 FILLER_150_648 ();
 FILLCELL_X4 FILLER_150_656 ();
 FILLCELL_X1 FILLER_150_660 ();
 FILLCELL_X1 FILLER_150_675 ();
 FILLCELL_X1 FILLER_150_685 ();
 FILLCELL_X1 FILLER_150_693 ();
 FILLCELL_X1 FILLER_150_708 ();
 FILLCELL_X4 FILLER_150_733 ();
 FILLCELL_X1 FILLER_150_737 ();
 FILLCELL_X4 FILLER_150_755 ();
 FILLCELL_X2 FILLER_150_768 ();
 FILLCELL_X1 FILLER_150_770 ();
 FILLCELL_X8 FILLER_150_792 ();
 FILLCELL_X2 FILLER_150_817 ();
 FILLCELL_X4 FILLER_150_834 ();
 FILLCELL_X1 FILLER_150_838 ();
 FILLCELL_X1 FILLER_150_850 ();
 FILLCELL_X2 FILLER_150_899 ();
 FILLCELL_X1 FILLER_150_901 ();
 FILLCELL_X2 FILLER_150_911 ();
 FILLCELL_X2 FILLER_150_937 ();
 FILLCELL_X8 FILLER_150_943 ();
 FILLCELL_X1 FILLER_150_967 ();
 FILLCELL_X16 FILLER_150_975 ();
 FILLCELL_X1 FILLER_150_991 ();
 FILLCELL_X32 FILLER_150_1030 ();
 FILLCELL_X2 FILLER_150_1084 ();
 FILLCELL_X1 FILLER_150_1086 ();
 FILLCELL_X32 FILLER_150_1109 ();
 FILLCELL_X32 FILLER_150_1141 ();
 FILLCELL_X16 FILLER_150_1173 ();
 FILLCELL_X8 FILLER_150_1189 ();
 FILLCELL_X4 FILLER_150_1197 ();
 FILLCELL_X8 FILLER_150_1204 ();
 FILLCELL_X4 FILLER_150_1212 ();
 FILLCELL_X16 FILLER_150_1219 ();
 FILLCELL_X4 FILLER_150_1235 ();
 FILLCELL_X1 FILLER_150_1239 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X8 FILLER_151_609 ();
 FILLCELL_X4 FILLER_151_617 ();
 FILLCELL_X2 FILLER_151_621 ();
 FILLCELL_X1 FILLER_151_623 ();
 FILLCELL_X32 FILLER_151_658 ();
 FILLCELL_X16 FILLER_151_690 ();
 FILLCELL_X4 FILLER_151_706 ();
 FILLCELL_X2 FILLER_151_710 ();
 FILLCELL_X16 FILLER_151_729 ();
 FILLCELL_X4 FILLER_151_745 ();
 FILLCELL_X2 FILLER_151_749 ();
 FILLCELL_X1 FILLER_151_751 ();
 FILLCELL_X32 FILLER_151_772 ();
 FILLCELL_X16 FILLER_151_804 ();
 FILLCELL_X2 FILLER_151_820 ();
 FILLCELL_X8 FILLER_151_827 ();
 FILLCELL_X4 FILLER_151_835 ();
 FILLCELL_X2 FILLER_151_839 ();
 FILLCELL_X1 FILLER_151_841 ();
 FILLCELL_X1 FILLER_151_862 ();
 FILLCELL_X8 FILLER_151_878 ();
 FILLCELL_X1 FILLER_151_886 ();
 FILLCELL_X1 FILLER_151_895 ();
 FILLCELL_X2 FILLER_151_918 ();
 FILLCELL_X1 FILLER_151_920 ();
 FILLCELL_X4 FILLER_151_928 ();
 FILLCELL_X2 FILLER_151_932 ();
 FILLCELL_X1 FILLER_151_936 ();
 FILLCELL_X1 FILLER_151_944 ();
 FILLCELL_X32 FILLER_151_982 ();
 FILLCELL_X32 FILLER_151_1014 ();
 FILLCELL_X1 FILLER_151_1046 ();
 FILLCELL_X1 FILLER_151_1072 ();
 FILLCELL_X1 FILLER_151_1077 ();
 FILLCELL_X4 FILLER_151_1084 ();
 FILLCELL_X1 FILLER_151_1101 ();
 FILLCELL_X2 FILLER_151_1118 ();
 FILLCELL_X1 FILLER_151_1120 ();
 FILLCELL_X32 FILLER_151_1123 ();
 FILLCELL_X32 FILLER_151_1155 ();
 FILLCELL_X16 FILLER_151_1187 ();
 FILLCELL_X8 FILLER_151_1203 ();
 FILLCELL_X4 FILLER_151_1211 ();
 FILLCELL_X2 FILLER_151_1215 ();
 FILLCELL_X1 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1221 ();
 FILLCELL_X4 FILLER_151_1229 ();
 FILLCELL_X1 FILLER_151_1239 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X8 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_617 ();
 FILLCELL_X2 FILLER_152_621 ();
 FILLCELL_X1 FILLER_152_623 ();
 FILLCELL_X8 FILLER_152_639 ();
 FILLCELL_X4 FILLER_152_647 ();
 FILLCELL_X2 FILLER_152_651 ();
 FILLCELL_X1 FILLER_152_653 ();
 FILLCELL_X2 FILLER_152_666 ();
 FILLCELL_X1 FILLER_152_668 ();
 FILLCELL_X16 FILLER_152_676 ();
 FILLCELL_X8 FILLER_152_699 ();
 FILLCELL_X1 FILLER_152_707 ();
 FILLCELL_X4 FILLER_152_733 ();
 FILLCELL_X2 FILLER_152_737 ();
 FILLCELL_X1 FILLER_152_739 ();
 FILLCELL_X32 FILLER_152_750 ();
 FILLCELL_X32 FILLER_152_782 ();
 FILLCELL_X4 FILLER_152_814 ();
 FILLCELL_X4 FILLER_152_825 ();
 FILLCELL_X2 FILLER_152_829 ();
 FILLCELL_X1 FILLER_152_831 ();
 FILLCELL_X8 FILLER_152_884 ();
 FILLCELL_X4 FILLER_152_909 ();
 FILLCELL_X8 FILLER_152_923 ();
 FILLCELL_X1 FILLER_152_931 ();
 FILLCELL_X1 FILLER_152_945 ();
 FILLCELL_X1 FILLER_152_949 ();
 FILLCELL_X1 FILLER_152_954 ();
 FILLCELL_X1 FILLER_152_958 ();
 FILLCELL_X1 FILLER_152_964 ();
 FILLCELL_X32 FILLER_152_968 ();
 FILLCELL_X4 FILLER_152_1000 ();
 FILLCELL_X2 FILLER_152_1004 ();
 FILLCELL_X1 FILLER_152_1006 ();
 FILLCELL_X8 FILLER_152_1011 ();
 FILLCELL_X4 FILLER_152_1019 ();
 FILLCELL_X2 FILLER_152_1023 ();
 FILLCELL_X1 FILLER_152_1069 ();
 FILLCELL_X1 FILLER_152_1084 ();
 FILLCELL_X32 FILLER_152_1123 ();
 FILLCELL_X32 FILLER_152_1155 ();
 FILLCELL_X8 FILLER_152_1187 ();
 FILLCELL_X4 FILLER_152_1195 ();
 FILLCELL_X2 FILLER_152_1199 ();
 FILLCELL_X2 FILLER_152_1204 ();
 FILLCELL_X1 FILLER_152_1206 ();
 FILLCELL_X16 FILLER_152_1210 ();
 FILLCELL_X8 FILLER_152_1226 ();
 FILLCELL_X4 FILLER_152_1234 ();
 FILLCELL_X2 FILLER_152_1238 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X4 FILLER_153_641 ();
 FILLCELL_X2 FILLER_153_645 ();
 FILLCELL_X1 FILLER_153_647 ();
 FILLCELL_X4 FILLER_153_674 ();
 FILLCELL_X2 FILLER_153_678 ();
 FILLCELL_X1 FILLER_153_680 ();
 FILLCELL_X1 FILLER_153_698 ();
 FILLCELL_X1 FILLER_153_716 ();
 FILLCELL_X4 FILLER_153_727 ();
 FILLCELL_X2 FILLER_153_731 ();
 FILLCELL_X1 FILLER_153_733 ();
 FILLCELL_X4 FILLER_153_762 ();
 FILLCELL_X4 FILLER_153_769 ();
 FILLCELL_X2 FILLER_153_773 ();
 FILLCELL_X1 FILLER_153_775 ();
 FILLCELL_X4 FILLER_153_780 ();
 FILLCELL_X2 FILLER_153_784 ();
 FILLCELL_X2 FILLER_153_803 ();
 FILLCELL_X1 FILLER_153_805 ();
 FILLCELL_X4 FILLER_153_857 ();
 FILLCELL_X32 FILLER_153_878 ();
 FILLCELL_X16 FILLER_153_910 ();
 FILLCELL_X8 FILLER_153_926 ();
 FILLCELL_X4 FILLER_153_934 ();
 FILLCELL_X2 FILLER_153_938 ();
 FILLCELL_X1 FILLER_153_940 ();
 FILLCELL_X32 FILLER_153_966 ();
 FILLCELL_X16 FILLER_153_998 ();
 FILLCELL_X8 FILLER_153_1014 ();
 FILLCELL_X2 FILLER_153_1022 ();
 FILLCELL_X1 FILLER_153_1024 ();
 FILLCELL_X1 FILLER_153_1066 ();
 FILLCELL_X1 FILLER_153_1081 ();
 FILLCELL_X1 FILLER_153_1103 ();
 FILLCELL_X32 FILLER_153_1125 ();
 FILLCELL_X32 FILLER_153_1157 ();
 FILLCELL_X16 FILLER_153_1189 ();
 FILLCELL_X8 FILLER_153_1205 ();
 FILLCELL_X2 FILLER_153_1213 ();
 FILLCELL_X1 FILLER_153_1215 ();
 FILLCELL_X2 FILLER_153_1219 ();
 FILLCELL_X1 FILLER_153_1221 ();
 FILLCELL_X8 FILLER_153_1225 ();
 FILLCELL_X1 FILLER_153_1233 ();
 FILLCELL_X2 FILLER_153_1238 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X8 FILLER_154_609 ();
 FILLCELL_X2 FILLER_154_617 ();
 FILLCELL_X4 FILLER_154_624 ();
 FILLCELL_X2 FILLER_154_628 ();
 FILLCELL_X1 FILLER_154_630 ();
 FILLCELL_X16 FILLER_154_632 ();
 FILLCELL_X8 FILLER_154_648 ();
 FILLCELL_X8 FILLER_154_673 ();
 FILLCELL_X4 FILLER_154_681 ();
 FILLCELL_X1 FILLER_154_685 ();
 FILLCELL_X2 FILLER_154_693 ();
 FILLCELL_X1 FILLER_154_695 ();
 FILLCELL_X2 FILLER_154_703 ();
 FILLCELL_X4 FILLER_154_719 ();
 FILLCELL_X1 FILLER_154_723 ();
 FILLCELL_X1 FILLER_154_751 ();
 FILLCELL_X4 FILLER_154_758 ();
 FILLCELL_X1 FILLER_154_762 ();
 FILLCELL_X2 FILLER_154_780 ();
 FILLCELL_X8 FILLER_154_824 ();
 FILLCELL_X4 FILLER_154_832 ();
 FILLCELL_X2 FILLER_154_836 ();
 FILLCELL_X1 FILLER_154_838 ();
 FILLCELL_X32 FILLER_154_843 ();
 FILLCELL_X32 FILLER_154_875 ();
 FILLCELL_X8 FILLER_154_907 ();
 FILLCELL_X2 FILLER_154_915 ();
 FILLCELL_X8 FILLER_154_921 ();
 FILLCELL_X8 FILLER_154_936 ();
 FILLCELL_X4 FILLER_154_944 ();
 FILLCELL_X2 FILLER_154_948 ();
 FILLCELL_X4 FILLER_154_967 ();
 FILLCELL_X2 FILLER_154_975 ();
 FILLCELL_X4 FILLER_154_987 ();
 FILLCELL_X1 FILLER_154_1005 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X8 FILLER_154_1048 ();
 FILLCELL_X4 FILLER_154_1056 ();
 FILLCELL_X8 FILLER_154_1063 ();
 FILLCELL_X1 FILLER_154_1071 ();
 FILLCELL_X4 FILLER_154_1077 ();
 FILLCELL_X1 FILLER_154_1081 ();
 FILLCELL_X4 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1122 ();
 FILLCELL_X32 FILLER_154_1154 ();
 FILLCELL_X16 FILLER_154_1186 ();
 FILLCELL_X8 FILLER_154_1202 ();
 FILLCELL_X2 FILLER_154_1210 ();
 FILLCELL_X1 FILLER_154_1212 ();
 FILLCELL_X8 FILLER_154_1216 ();
 FILLCELL_X8 FILLER_154_1227 ();
 FILLCELL_X4 FILLER_154_1235 ();
 FILLCELL_X1 FILLER_154_1239 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X8 FILLER_155_673 ();
 FILLCELL_X4 FILLER_155_681 ();
 FILLCELL_X8 FILLER_155_702 ();
 FILLCELL_X8 FILLER_155_727 ();
 FILLCELL_X1 FILLER_155_735 ();
 FILLCELL_X4 FILLER_155_740 ();
 FILLCELL_X1 FILLER_155_744 ();
 FILLCELL_X1 FILLER_155_749 ();
 FILLCELL_X16 FILLER_155_773 ();
 FILLCELL_X4 FILLER_155_789 ();
 FILLCELL_X2 FILLER_155_793 ();
 FILLCELL_X1 FILLER_155_795 ();
 FILLCELL_X32 FILLER_155_821 ();
 FILLCELL_X32 FILLER_155_853 ();
 FILLCELL_X8 FILLER_155_885 ();
 FILLCELL_X4 FILLER_155_893 ();
 FILLCELL_X1 FILLER_155_897 ();
 FILLCELL_X4 FILLER_155_901 ();
 FILLCELL_X1 FILLER_155_905 ();
 FILLCELL_X16 FILLER_155_936 ();
 FILLCELL_X8 FILLER_155_952 ();
 FILLCELL_X4 FILLER_155_960 ();
 FILLCELL_X2 FILLER_155_964 ();
 FILLCELL_X1 FILLER_155_966 ();
 FILLCELL_X1 FILLER_155_970 ();
 FILLCELL_X2 FILLER_155_991 ();
 FILLCELL_X2 FILLER_155_996 ();
 FILLCELL_X4 FILLER_155_1012 ();
 FILLCELL_X2 FILLER_155_1016 ();
 FILLCELL_X1 FILLER_155_1023 ();
 FILLCELL_X32 FILLER_155_1037 ();
 FILLCELL_X16 FILLER_155_1069 ();
 FILLCELL_X4 FILLER_155_1085 ();
 FILLCELL_X1 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1111 ();
 FILLCELL_X32 FILLER_155_1143 ();
 FILLCELL_X32 FILLER_155_1175 ();
 FILLCELL_X8 FILLER_155_1207 ();
 FILLCELL_X4 FILLER_155_1215 ();
 FILLCELL_X2 FILLER_155_1219 ();
 FILLCELL_X1 FILLER_155_1221 ();
 FILLCELL_X8 FILLER_155_1225 ();
 FILLCELL_X1 FILLER_155_1233 ();
 FILLCELL_X2 FILLER_155_1237 ();
 FILLCELL_X1 FILLER_155_1239 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X16 FILLER_156_703 ();
 FILLCELL_X8 FILLER_156_719 ();
 FILLCELL_X4 FILLER_156_727 ();
 FILLCELL_X1 FILLER_156_731 ();
 FILLCELL_X32 FILLER_156_751 ();
 FILLCELL_X4 FILLER_156_783 ();
 FILLCELL_X1 FILLER_156_787 ();
 FILLCELL_X4 FILLER_156_791 ();
 FILLCELL_X2 FILLER_156_795 ();
 FILLCELL_X32 FILLER_156_810 ();
 FILLCELL_X8 FILLER_156_842 ();
 FILLCELL_X4 FILLER_156_850 ();
 FILLCELL_X2 FILLER_156_854 ();
 FILLCELL_X1 FILLER_156_856 ();
 FILLCELL_X2 FILLER_156_871 ();
 FILLCELL_X1 FILLER_156_876 ();
 FILLCELL_X16 FILLER_156_883 ();
 FILLCELL_X1 FILLER_156_899 ();
 FILLCELL_X16 FILLER_156_934 ();
 FILLCELL_X8 FILLER_156_950 ();
 FILLCELL_X2 FILLER_156_958 ();
 FILLCELL_X2 FILLER_156_992 ();
 FILLCELL_X1 FILLER_156_994 ();
 FILLCELL_X2 FILLER_156_1020 ();
 FILLCELL_X32 FILLER_156_1043 ();
 FILLCELL_X32 FILLER_156_1075 ();
 FILLCELL_X32 FILLER_156_1107 ();
 FILLCELL_X32 FILLER_156_1139 ();
 FILLCELL_X32 FILLER_156_1171 ();
 FILLCELL_X32 FILLER_156_1203 ();
 FILLCELL_X4 FILLER_156_1235 ();
 FILLCELL_X1 FILLER_156_1239 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X8 FILLER_157_737 ();
 FILLCELL_X2 FILLER_157_745 ();
 FILLCELL_X8 FILLER_157_755 ();
 FILLCELL_X16 FILLER_157_782 ();
 FILLCELL_X1 FILLER_157_798 ();
 FILLCELL_X1 FILLER_157_803 ();
 FILLCELL_X8 FILLER_157_818 ();
 FILLCELL_X2 FILLER_157_826 ();
 FILLCELL_X1 FILLER_157_828 ();
 FILLCELL_X2 FILLER_157_885 ();
 FILLCELL_X1 FILLER_157_887 ();
 FILLCELL_X16 FILLER_157_891 ();
 FILLCELL_X8 FILLER_157_907 ();
 FILLCELL_X4 FILLER_157_915 ();
 FILLCELL_X1 FILLER_157_932 ();
 FILLCELL_X16 FILLER_157_943 ();
 FILLCELL_X8 FILLER_157_959 ();
 FILLCELL_X1 FILLER_157_986 ();
 FILLCELL_X1 FILLER_157_990 ();
 FILLCELL_X1 FILLER_157_998 ();
 FILLCELL_X1 FILLER_157_1010 ();
 FILLCELL_X2 FILLER_157_1032 ();
 FILLCELL_X1 FILLER_157_1034 ();
 FILLCELL_X32 FILLER_157_1056 ();
 FILLCELL_X32 FILLER_157_1088 ();
 FILLCELL_X32 FILLER_157_1120 ();
 FILLCELL_X32 FILLER_157_1152 ();
 FILLCELL_X32 FILLER_157_1184 ();
 FILLCELL_X16 FILLER_157_1216 ();
 FILLCELL_X8 FILLER_157_1232 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X16 FILLER_158_760 ();
 FILLCELL_X8 FILLER_158_823 ();
 FILLCELL_X2 FILLER_158_831 ();
 FILLCELL_X8 FILLER_158_839 ();
 FILLCELL_X2 FILLER_158_847 ();
 FILLCELL_X2 FILLER_158_901 ();
 FILLCELL_X16 FILLER_158_958 ();
 FILLCELL_X8 FILLER_158_974 ();
 FILLCELL_X4 FILLER_158_982 ();
 FILLCELL_X2 FILLER_158_986 ();
 FILLCELL_X1 FILLER_158_1010 ();
 FILLCELL_X2 FILLER_158_1032 ();
 FILLCELL_X1 FILLER_158_1034 ();
 FILLCELL_X4 FILLER_158_1040 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X16 FILLER_159_737 ();
 FILLCELL_X8 FILLER_159_753 ();
 FILLCELL_X4 FILLER_159_761 ();
 FILLCELL_X2 FILLER_159_765 ();
 FILLCELL_X8 FILLER_159_770 ();
 FILLCELL_X4 FILLER_159_778 ();
 FILLCELL_X1 FILLER_159_782 ();
 FILLCELL_X1 FILLER_159_808 ();
 FILLCELL_X2 FILLER_159_826 ();
 FILLCELL_X1 FILLER_159_828 ();
 FILLCELL_X1 FILLER_159_879 ();
 FILLCELL_X4 FILLER_159_890 ();
 FILLCELL_X1 FILLER_159_894 ();
 FILLCELL_X8 FILLER_159_899 ();
 FILLCELL_X4 FILLER_159_907 ();
 FILLCELL_X1 FILLER_159_911 ();
 FILLCELL_X4 FILLER_159_920 ();
 FILLCELL_X2 FILLER_159_924 ();
 FILLCELL_X1 FILLER_159_926 ();
 FILLCELL_X1 FILLER_159_945 ();
 FILLCELL_X16 FILLER_159_967 ();
 FILLCELL_X2 FILLER_159_1002 ();
 FILLCELL_X32 FILLER_159_1039 ();
 FILLCELL_X32 FILLER_159_1071 ();
 FILLCELL_X32 FILLER_159_1103 ();
 FILLCELL_X32 FILLER_159_1135 ();
 FILLCELL_X32 FILLER_159_1167 ();
 FILLCELL_X32 FILLER_159_1199 ();
 FILLCELL_X8 FILLER_159_1231 ();
 FILLCELL_X1 FILLER_159_1239 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X16 FILLER_160_728 ();
 FILLCELL_X8 FILLER_160_744 ();
 FILLCELL_X4 FILLER_160_752 ();
 FILLCELL_X2 FILLER_160_756 ();
 FILLCELL_X1 FILLER_160_758 ();
 FILLCELL_X1 FILLER_160_818 ();
 FILLCELL_X16 FILLER_160_822 ();
 FILLCELL_X8 FILLER_160_838 ();
 FILLCELL_X4 FILLER_160_846 ();
 FILLCELL_X2 FILLER_160_850 ();
 FILLCELL_X1 FILLER_160_852 ();
 FILLCELL_X8 FILLER_160_899 ();
 FILLCELL_X4 FILLER_160_907 ();
 FILLCELL_X1 FILLER_160_914 ();
 FILLCELL_X4 FILLER_160_918 ();
 FILLCELL_X4 FILLER_160_929 ();
 FILLCELL_X1 FILLER_160_933 ();
 FILLCELL_X1 FILLER_160_938 ();
 FILLCELL_X4 FILLER_160_976 ();
 FILLCELL_X16 FILLER_160_984 ();
 FILLCELL_X8 FILLER_160_1000 ();
 FILLCELL_X4 FILLER_160_1008 ();
 FILLCELL_X8 FILLER_160_1022 ();
 FILLCELL_X1 FILLER_160_1030 ();
 FILLCELL_X32 FILLER_160_1050 ();
 FILLCELL_X32 FILLER_160_1082 ();
 FILLCELL_X32 FILLER_160_1114 ();
 FILLCELL_X32 FILLER_160_1146 ();
 FILLCELL_X32 FILLER_160_1178 ();
 FILLCELL_X16 FILLER_160_1210 ();
 FILLCELL_X8 FILLER_160_1226 ();
 FILLCELL_X4 FILLER_160_1234 ();
 FILLCELL_X2 FILLER_160_1238 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X4 FILLER_161_769 ();
 FILLCELL_X1 FILLER_161_773 ();
 FILLCELL_X1 FILLER_161_784 ();
 FILLCELL_X1 FILLER_161_805 ();
 FILLCELL_X2 FILLER_161_815 ();
 FILLCELL_X1 FILLER_161_817 ();
 FILLCELL_X16 FILLER_161_822 ();
 FILLCELL_X8 FILLER_161_838 ();
 FILLCELL_X1 FILLER_161_846 ();
 FILLCELL_X16 FILLER_161_862 ();
 FILLCELL_X16 FILLER_161_887 ();
 FILLCELL_X2 FILLER_161_903 ();
 FILLCELL_X1 FILLER_161_934 ();
 FILLCELL_X2 FILLER_161_962 ();
 FILLCELL_X16 FILLER_161_970 ();
 FILLCELL_X8 FILLER_161_986 ();
 FILLCELL_X1 FILLER_161_994 ();
 FILLCELL_X32 FILLER_161_999 ();
 FILLCELL_X32 FILLER_161_1031 ();
 FILLCELL_X32 FILLER_161_1063 ();
 FILLCELL_X32 FILLER_161_1095 ();
 FILLCELL_X32 FILLER_161_1127 ();
 FILLCELL_X32 FILLER_161_1159 ();
 FILLCELL_X32 FILLER_161_1191 ();
 FILLCELL_X16 FILLER_161_1223 ();
 FILLCELL_X1 FILLER_161_1239 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X16 FILLER_162_760 ();
 FILLCELL_X8 FILLER_162_776 ();
 FILLCELL_X4 FILLER_162_784 ();
 FILLCELL_X2 FILLER_162_788 ();
 FILLCELL_X4 FILLER_162_799 ();
 FILLCELL_X2 FILLER_162_803 ();
 FILLCELL_X16 FILLER_162_822 ();
 FILLCELL_X8 FILLER_162_868 ();
 FILLCELL_X16 FILLER_162_893 ();
 FILLCELL_X1 FILLER_162_928 ();
 FILLCELL_X2 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_960 ();
 FILLCELL_X4 FILLER_162_1011 ();
 FILLCELL_X2 FILLER_162_1015 ();
 FILLCELL_X1 FILLER_162_1017 ();
 FILLCELL_X8 FILLER_162_1022 ();
 FILLCELL_X2 FILLER_162_1030 ();
 FILLCELL_X1 FILLER_162_1032 ();
 FILLCELL_X32 FILLER_162_1037 ();
 FILLCELL_X32 FILLER_162_1069 ();
 FILLCELL_X32 FILLER_162_1101 ();
 FILLCELL_X32 FILLER_162_1133 ();
 FILLCELL_X32 FILLER_162_1165 ();
 FILLCELL_X32 FILLER_162_1197 ();
 FILLCELL_X8 FILLER_162_1229 ();
 FILLCELL_X2 FILLER_162_1237 ();
 FILLCELL_X1 FILLER_162_1239 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X1 FILLER_163_833 ();
 FILLCELL_X1 FILLER_163_838 ();
 FILLCELL_X2 FILLER_163_843 ();
 FILLCELL_X4 FILLER_163_877 ();
 FILLCELL_X1 FILLER_163_881 ();
 FILLCELL_X32 FILLER_163_886 ();
 FILLCELL_X8 FILLER_163_918 ();
 FILLCELL_X4 FILLER_163_926 ();
 FILLCELL_X1 FILLER_163_930 ();
 FILLCELL_X32 FILLER_163_951 ();
 FILLCELL_X8 FILLER_163_983 ();
 FILLCELL_X1 FILLER_163_991 ();
 FILLCELL_X4 FILLER_163_1019 ();
 FILLCELL_X32 FILLER_163_1027 ();
 FILLCELL_X32 FILLER_163_1059 ();
 FILLCELL_X32 FILLER_163_1091 ();
 FILLCELL_X32 FILLER_163_1123 ();
 FILLCELL_X32 FILLER_163_1155 ();
 FILLCELL_X32 FILLER_163_1187 ();
 FILLCELL_X16 FILLER_163_1219 ();
 FILLCELL_X4 FILLER_163_1235 ();
 FILLCELL_X1 FILLER_163_1239 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X8 FILLER_164_824 ();
 FILLCELL_X2 FILLER_164_832 ();
 FILLCELL_X1 FILLER_164_834 ();
 FILLCELL_X32 FILLER_164_852 ();
 FILLCELL_X32 FILLER_164_884 ();
 FILLCELL_X32 FILLER_164_916 ();
 FILLCELL_X32 FILLER_164_948 ();
 FILLCELL_X16 FILLER_164_980 ();
 FILLCELL_X4 FILLER_164_996 ();
 FILLCELL_X2 FILLER_164_1000 ();
 FILLCELL_X1 FILLER_164_1002 ();
 FILLCELL_X2 FILLER_164_1011 ();
 FILLCELL_X4 FILLER_164_1017 ();
 FILLCELL_X2 FILLER_164_1021 ();
 FILLCELL_X1 FILLER_164_1023 ();
 FILLCELL_X32 FILLER_164_1028 ();
 FILLCELL_X32 FILLER_164_1060 ();
 FILLCELL_X32 FILLER_164_1092 ();
 FILLCELL_X32 FILLER_164_1124 ();
 FILLCELL_X32 FILLER_164_1156 ();
 FILLCELL_X32 FILLER_164_1188 ();
 FILLCELL_X16 FILLER_164_1220 ();
 FILLCELL_X4 FILLER_164_1236 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X8 FILLER_165_577 ();
 FILLCELL_X4 FILLER_165_585 ();
 FILLCELL_X32 FILLER_165_593 ();
 FILLCELL_X32 FILLER_165_625 ();
 FILLCELL_X32 FILLER_165_657 ();
 FILLCELL_X32 FILLER_165_689 ();
 FILLCELL_X32 FILLER_165_721 ();
 FILLCELL_X32 FILLER_165_753 ();
 FILLCELL_X32 FILLER_165_785 ();
 FILLCELL_X32 FILLER_165_817 ();
 FILLCELL_X32 FILLER_165_849 ();
 FILLCELL_X32 FILLER_165_881 ();
 FILLCELL_X32 FILLER_165_913 ();
 FILLCELL_X32 FILLER_165_945 ();
 FILLCELL_X32 FILLER_165_977 ();
 FILLCELL_X32 FILLER_165_1009 ();
 FILLCELL_X32 FILLER_165_1041 ();
 FILLCELL_X32 FILLER_165_1073 ();
 FILLCELL_X32 FILLER_165_1105 ();
 FILLCELL_X32 FILLER_165_1137 ();
 FILLCELL_X32 FILLER_165_1169 ();
 FILLCELL_X32 FILLER_165_1201 ();
 FILLCELL_X4 FILLER_165_1233 ();
 FILLCELL_X2 FILLER_165_1237 ();
 FILLCELL_X1 FILLER_165_1239 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X16 FILLER_166_577 ();
 FILLCELL_X4 FILLER_166_597 ();
 FILLCELL_X2 FILLER_166_601 ();
 FILLCELL_X4 FILLER_166_607 ();
 FILLCELL_X2 FILLER_166_611 ();
 FILLCELL_X4 FILLER_166_617 ();
 FILLCELL_X1 FILLER_166_621 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X4 FILLER_166_632 ();
 FILLCELL_X8 FILLER_166_639 ();
 FILLCELL_X2 FILLER_166_647 ();
 FILLCELL_X1 FILLER_166_649 ();
 FILLCELL_X16 FILLER_166_656 ();
 FILLCELL_X8 FILLER_166_672 ();
 FILLCELL_X32 FILLER_166_683 ();
 FILLCELL_X1 FILLER_166_715 ();
 FILLCELL_X32 FILLER_166_719 ();
 FILLCELL_X16 FILLER_166_751 ();
 FILLCELL_X8 FILLER_166_767 ();
 FILLCELL_X16 FILLER_166_778 ();
 FILLCELL_X2 FILLER_166_794 ();
 FILLCELL_X1 FILLER_166_796 ();
 FILLCELL_X16 FILLER_166_800 ();
 FILLCELL_X8 FILLER_166_816 ();
 FILLCELL_X2 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_835 ();
 FILLCELL_X8 FILLER_166_867 ();
 FILLCELL_X4 FILLER_166_878 ();
 FILLCELL_X2 FILLER_166_882 ();
 FILLCELL_X1 FILLER_166_884 ();
 FILLCELL_X16 FILLER_166_888 ();
 FILLCELL_X4 FILLER_166_904 ();
 FILLCELL_X2 FILLER_166_908 ();
 FILLCELL_X8 FILLER_166_913 ();
 FILLCELL_X2 FILLER_166_921 ();
 FILLCELL_X16 FILLER_166_926 ();
 FILLCELL_X8 FILLER_166_942 ();
 FILLCELL_X4 FILLER_166_950 ();
 FILLCELL_X32 FILLER_166_957 ();
 FILLCELL_X4 FILLER_166_989 ();
 FILLCELL_X1 FILLER_166_993 ();
 FILLCELL_X8 FILLER_166_1000 ();
 FILLCELL_X4 FILLER_166_1008 ();
 FILLCELL_X8 FILLER_166_1015 ();
 FILLCELL_X2 FILLER_166_1023 ();
 FILLCELL_X1 FILLER_166_1025 ();
 FILLCELL_X32 FILLER_166_1029 ();
 FILLCELL_X32 FILLER_166_1061 ();
 FILLCELL_X32 FILLER_166_1093 ();
 FILLCELL_X32 FILLER_166_1125 ();
 FILLCELL_X32 FILLER_166_1157 ();
 FILLCELL_X32 FILLER_166_1189 ();
 FILLCELL_X16 FILLER_166_1221 ();
 FILLCELL_X2 FILLER_166_1237 ();
 FILLCELL_X1 FILLER_166_1239 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X16 FILLER_167_449 ();
 FILLCELL_X4 FILLER_167_465 ();
 FILLCELL_X1 FILLER_167_469 ();
 FILLCELL_X8 FILLER_167_473 ();
 FILLCELL_X1 FILLER_167_481 ();
 FILLCELL_X8 FILLER_167_485 ();
 FILLCELL_X1 FILLER_167_493 ();
 FILLCELL_X8 FILLER_167_498 ();
 FILLCELL_X1 FILLER_167_506 ();
 FILLCELL_X16 FILLER_167_510 ();
 FILLCELL_X4 FILLER_167_526 ();
 FILLCELL_X1 FILLER_167_530 ();
 FILLCELL_X2 FILLER_167_543 ();
 FILLCELL_X2 FILLER_167_549 ();
 FILLCELL_X4 FILLER_167_555 ();
 FILLCELL_X1 FILLER_167_559 ();
 FILLCELL_X8 FILLER_167_564 ();
 FILLCELL_X4 FILLER_167_572 ();
 FILLCELL_X1 FILLER_167_576 ();
 FILLCELL_X2 FILLER_167_592 ();
 FILLCELL_X1 FILLER_167_598 ();
 FILLCELL_X1 FILLER_167_607 ();
 FILLCELL_X4 FILLER_167_620 ();
 FILLCELL_X1 FILLER_167_624 ();
 FILLCELL_X2 FILLER_167_629 ();
 FILLCELL_X2 FILLER_167_636 ();
 FILLCELL_X1 FILLER_167_638 ();
 FILLCELL_X2 FILLER_167_649 ();
 FILLCELL_X1 FILLER_167_651 ();
 FILLCELL_X2 FILLER_167_656 ();
 FILLCELL_X1 FILLER_167_658 ();
 FILLCELL_X2 FILLER_167_662 ();
 FILLCELL_X1 FILLER_167_664 ();
 FILLCELL_X1 FILLER_167_668 ();
 FILLCELL_X1 FILLER_167_676 ();
 FILLCELL_X4 FILLER_167_686 ();
 FILLCELL_X1 FILLER_167_690 ();
 FILLCELL_X4 FILLER_167_697 ();
 FILLCELL_X2 FILLER_167_701 ();
 FILLCELL_X1 FILLER_167_703 ();
 FILLCELL_X16 FILLER_167_713 ();
 FILLCELL_X8 FILLER_167_729 ();
 FILLCELL_X4 FILLER_167_737 ();
 FILLCELL_X2 FILLER_167_741 ();
 FILLCELL_X4 FILLER_167_746 ();
 FILLCELL_X8 FILLER_167_753 ();
 FILLCELL_X4 FILLER_167_761 ();
 FILLCELL_X2 FILLER_167_765 ();
 FILLCELL_X1 FILLER_167_767 ();
 FILLCELL_X2 FILLER_167_771 ();
 FILLCELL_X1 FILLER_167_785 ();
 FILLCELL_X2 FILLER_167_795 ();
 FILLCELL_X2 FILLER_167_800 ();
 FILLCELL_X1 FILLER_167_802 ();
 FILLCELL_X1 FILLER_167_810 ();
 FILLCELL_X1 FILLER_167_814 ();
 FILLCELL_X1 FILLER_167_821 ();
 FILLCELL_X1 FILLER_167_825 ();
 FILLCELL_X4 FILLER_167_829 ();
 FILLCELL_X2 FILLER_167_833 ();
 FILLCELL_X1 FILLER_167_835 ();
 FILLCELL_X4 FILLER_167_839 ();
 FILLCELL_X2 FILLER_167_846 ();
 FILLCELL_X1 FILLER_167_848 ();
 FILLCELL_X4 FILLER_167_853 ();
 FILLCELL_X2 FILLER_167_863 ();
 FILLCELL_X1 FILLER_167_865 ();
 FILLCELL_X1 FILLER_167_869 ();
 FILLCELL_X8 FILLER_167_873 ();
 FILLCELL_X1 FILLER_167_881 ();
 FILLCELL_X16 FILLER_167_886 ();
 FILLCELL_X4 FILLER_167_902 ();
 FILLCELL_X1 FILLER_167_906 ();
 FILLCELL_X4 FILLER_167_910 ();
 FILLCELL_X1 FILLER_167_923 ();
 FILLCELL_X4 FILLER_167_930 ();
 FILLCELL_X1 FILLER_167_934 ();
 FILLCELL_X1 FILLER_167_945 ();
 FILLCELL_X8 FILLER_167_949 ();
 FILLCELL_X1 FILLER_167_957 ();
 FILLCELL_X4 FILLER_167_967 ();
 FILLCELL_X1 FILLER_167_971 ();
 FILLCELL_X16 FILLER_167_975 ();
 FILLCELL_X8 FILLER_167_991 ();
 FILLCELL_X4 FILLER_167_999 ();
 FILLCELL_X4 FILLER_167_1009 ();
 FILLCELL_X1 FILLER_167_1013 ();
 FILLCELL_X2 FILLER_167_1029 ();
 FILLCELL_X1 FILLER_167_1031 ();
 FILLCELL_X16 FILLER_167_1035 ();
 FILLCELL_X4 FILLER_167_1051 ();
 FILLCELL_X2 FILLER_167_1055 ();
 FILLCELL_X1 FILLER_167_1057 ();
 FILLCELL_X8 FILLER_167_1062 ();
 FILLCELL_X4 FILLER_167_1070 ();
 FILLCELL_X1 FILLER_167_1074 ();
 FILLCELL_X4 FILLER_167_1078 ();
 FILLCELL_X32 FILLER_167_1085 ();
 FILLCELL_X32 FILLER_167_1117 ();
 FILLCELL_X32 FILLER_167_1149 ();
 FILLCELL_X32 FILLER_167_1181 ();
 FILLCELL_X16 FILLER_167_1213 ();
 FILLCELL_X8 FILLER_167_1229 ();
 FILLCELL_X2 FILLER_167_1237 ();
 FILLCELL_X1 FILLER_167_1239 ();
endmodule
