module dma_controller (clk,
    debug_has_active_channels,
    rst_n,
    channel_busy,
    channel_done,
    channel_dst_addr,
    channel_enable,
    channel_error,
    channel_length,
    channel_mode,
    channel_src_addr,
    channel_start,
    debug_active_channels,
    debug_channel_state,
    debug_transfer_count,
    dst_addr,
    dst_wdata,
    dst_wready,
    dst_write,
    dst_wstrb,
    src_addr,
    src_rdata,
    src_read,
    src_rready,
    src_rvalid);
 input clk;
 output debug_has_active_channels;
 input rst_n;
 output [3:0] channel_busy;
 output [3:0] channel_done;
 input [127:0] channel_dst_addr;
 input [3:0] channel_enable;
 output [3:0] channel_error;
 input [127:0] channel_length;
 input [7:0] channel_mode;
 input [127:0] channel_src_addr;
 input [3:0] channel_start;
 output [3:0] debug_active_channels;
 output [11:0] debug_channel_state;
 output [127:0] debug_transfer_count;
 output [127:0] dst_addr;
 output [127:0] dst_wdata;
 input [3:0] dst_wready;
 output [3:0] dst_write;
 output [15:0] dst_wstrb;
 output [127:0] src_addr;
 input [127:0] src_rdata;
 output [3:0] src_read;
 output [3:0] src_rready;
 input [3:0] src_rvalid;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire clknet_0_clk;
 wire \active_channel_count[0] ;
 wire \active_channel_count[1] ;
 wire \active_channel_count[2] ;
 wire \active_channel_count[3] ;
 wire \channel_state[0][0] ;
 wire \channel_state[0][1] ;
 wire \channel_state[0][2] ;
 wire \channel_state[0][3] ;
 wire \channel_state[0][4] ;
 wire \channel_state[0][5] ;
 wire \channel_state[1][0] ;
 wire \channel_state[1][1] ;
 wire \channel_state[1][2] ;
 wire \channel_state[1][3] ;
 wire \channel_state[1][4] ;
 wire \channel_state[1][5] ;
 wire \channel_state[2][0] ;
 wire \channel_state[2][1] ;
 wire \channel_state[2][2] ;
 wire \channel_state[2][3] ;
 wire \channel_state[2][4] ;
 wire \channel_state[2][5] ;
 wire \channel_state[3][0] ;
 wire \channel_state[3][1] ;
 wire \channel_state[3][2] ;
 wire \channel_state[3][3] ;
 wire \channel_state[3][4] ;
 wire \channel_state[3][5] ;
 wire \transfer_count[0][0] ;
 wire \transfer_count[0][10] ;
 wire \transfer_count[0][11] ;
 wire \transfer_count[0][12] ;
 wire \transfer_count[0][13] ;
 wire \transfer_count[0][14] ;
 wire \transfer_count[0][15] ;
 wire \transfer_count[0][16] ;
 wire \transfer_count[0][17] ;
 wire \transfer_count[0][18] ;
 wire \transfer_count[0][19] ;
 wire \transfer_count[0][1] ;
 wire \transfer_count[0][20] ;
 wire \transfer_count[0][21] ;
 wire \transfer_count[0][22] ;
 wire \transfer_count[0][23] ;
 wire \transfer_count[0][24] ;
 wire \transfer_count[0][25] ;
 wire \transfer_count[0][26] ;
 wire \transfer_count[0][27] ;
 wire \transfer_count[0][28] ;
 wire \transfer_count[0][29] ;
 wire \transfer_count[0][2] ;
 wire \transfer_count[0][30] ;
 wire \transfer_count[0][31] ;
 wire \transfer_count[0][3] ;
 wire \transfer_count[0][4] ;
 wire \transfer_count[0][5] ;
 wire \transfer_count[0][6] ;
 wire \transfer_count[0][7] ;
 wire \transfer_count[0][8] ;
 wire \transfer_count[0][9] ;
 wire \transfer_count[1][0] ;
 wire \transfer_count[1][10] ;
 wire \transfer_count[1][11] ;
 wire \transfer_count[1][12] ;
 wire \transfer_count[1][13] ;
 wire \transfer_count[1][14] ;
 wire \transfer_count[1][15] ;
 wire \transfer_count[1][16] ;
 wire \transfer_count[1][17] ;
 wire \transfer_count[1][18] ;
 wire \transfer_count[1][19] ;
 wire \transfer_count[1][1] ;
 wire \transfer_count[1][20] ;
 wire \transfer_count[1][21] ;
 wire \transfer_count[1][22] ;
 wire \transfer_count[1][23] ;
 wire \transfer_count[1][24] ;
 wire \transfer_count[1][25] ;
 wire \transfer_count[1][26] ;
 wire \transfer_count[1][27] ;
 wire \transfer_count[1][28] ;
 wire \transfer_count[1][29] ;
 wire \transfer_count[1][2] ;
 wire \transfer_count[1][30] ;
 wire \transfer_count[1][31] ;
 wire \transfer_count[1][3] ;
 wire \transfer_count[1][4] ;
 wire \transfer_count[1][5] ;
 wire \transfer_count[1][6] ;
 wire \transfer_count[1][7] ;
 wire \transfer_count[1][8] ;
 wire \transfer_count[1][9] ;
 wire \transfer_count[2][0] ;
 wire \transfer_count[2][10] ;
 wire \transfer_count[2][11] ;
 wire \transfer_count[2][12] ;
 wire \transfer_count[2][13] ;
 wire \transfer_count[2][14] ;
 wire \transfer_count[2][15] ;
 wire \transfer_count[2][16] ;
 wire \transfer_count[2][17] ;
 wire \transfer_count[2][18] ;
 wire \transfer_count[2][19] ;
 wire \transfer_count[2][1] ;
 wire \transfer_count[2][20] ;
 wire \transfer_count[2][21] ;
 wire \transfer_count[2][22] ;
 wire \transfer_count[2][23] ;
 wire \transfer_count[2][24] ;
 wire \transfer_count[2][25] ;
 wire \transfer_count[2][26] ;
 wire \transfer_count[2][27] ;
 wire \transfer_count[2][28] ;
 wire \transfer_count[2][29] ;
 wire \transfer_count[2][2] ;
 wire \transfer_count[2][30] ;
 wire \transfer_count[2][31] ;
 wire \transfer_count[2][3] ;
 wire \transfer_count[2][4] ;
 wire \transfer_count[2][5] ;
 wire \transfer_count[2][6] ;
 wire \transfer_count[2][7] ;
 wire \transfer_count[2][8] ;
 wire \transfer_count[2][9] ;
 wire \transfer_count[3][0] ;
 wire \transfer_count[3][10] ;
 wire \transfer_count[3][11] ;
 wire \transfer_count[3][12] ;
 wire \transfer_count[3][13] ;
 wire \transfer_count[3][14] ;
 wire \transfer_count[3][15] ;
 wire \transfer_count[3][16] ;
 wire \transfer_count[3][17] ;
 wire \transfer_count[3][18] ;
 wire \transfer_count[3][19] ;
 wire \transfer_count[3][1] ;
 wire \transfer_count[3][20] ;
 wire \transfer_count[3][21] ;
 wire \transfer_count[3][22] ;
 wire \transfer_count[3][23] ;
 wire \transfer_count[3][24] ;
 wire \transfer_count[3][25] ;
 wire \transfer_count[3][26] ;
 wire \transfer_count[3][27] ;
 wire \transfer_count[3][28] ;
 wire \transfer_count[3][29] ;
 wire \transfer_count[3][2] ;
 wire \transfer_count[3][30] ;
 wire \transfer_count[3][31] ;
 wire \transfer_count[3][3] ;
 wire \transfer_count[3][4] ;
 wire \transfer_count[3][5] ;
 wire \transfer_count[3][6] ;
 wire \transfer_count[3][7] ;
 wire \transfer_count[3][8] ;
 wire \transfer_count[3][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X8 _1868_ (.A(rst_n),
    .Z(_1087_));
 BUF_X4 _1869_ (.A(_1087_),
    .Z(_1088_));
 BUF_X4 _1870_ (.A(_1088_),
    .Z(_1089_));
 BUF_X4 _1871_ (.A(_1089_),
    .Z(_1090_));
 CLKBUF_X3 _1872_ (.A(\channel_state[2][0] ),
    .Z(_1091_));
 NOR2_X1 _1873_ (.A1(\channel_state[2][4] ),
    .A2(_1091_),
    .ZN(_1092_));
 INV_X1 _1874_ (.A(net129),
    .ZN(_1093_));
 BUF_X2 _1875_ (.A(channel_enable[2]),
    .Z(_1094_));
 INV_X1 _1876_ (.A(_1094_),
    .ZN(_1095_));
 AOI21_X1 _1877_ (.A(_1093_),
    .B1(_1091_),
    .B2(_1095_),
    .ZN(_1096_));
 OAI21_X1 _1878_ (.A(_1090_),
    .B1(_1092_),
    .B2(_1096_),
    .ZN(_0014_));
 BUF_X2 _1879_ (.A(\transfer_count[2][5] ),
    .Z(_1097_));
 CLKBUF_X3 _1880_ (.A(\transfer_count[2][3] ),
    .Z(_1098_));
 BUF_X2 _1881_ (.A(\transfer_count[2][4] ),
    .Z(_1099_));
 CLKBUF_X3 _1882_ (.A(\transfer_count[2][2] ),
    .Z(_1100_));
 NAND3_X2 _1883_ (.A1(_1100_),
    .A2(\transfer_count[2][1] ),
    .A3(\transfer_count[2][0] ),
    .ZN(_1101_));
 INV_X1 _1884_ (.A(_1101_),
    .ZN(_1102_));
 NAND3_X1 _1885_ (.A1(_1098_),
    .A2(_1099_),
    .A3(_1102_),
    .ZN(_1103_));
 XOR2_X2 _1886_ (.A(_1097_),
    .B(_1103_),
    .Z(_1486_));
 INV_X1 _1887_ (.A(\transfer_count[2][13] ),
    .ZN(_1104_));
 BUF_X1 _1888_ (.A(\transfer_count[2][12] ),
    .Z(_1105_));
 INV_X1 _1889_ (.A(_1105_),
    .ZN(_1106_));
 INV_X1 _1890_ (.A(\transfer_count[2][11] ),
    .ZN(_1107_));
 BUF_X2 _1891_ (.A(\transfer_count[2][7] ),
    .Z(_1108_));
 NAND4_X4 _1892_ (.A1(_1100_),
    .A2(\transfer_count[2][1] ),
    .A3(\transfer_count[2][0] ),
    .A4(_1108_),
    .ZN(_1109_));
 INV_X1 _1893_ (.A(\transfer_count[2][10] ),
    .ZN(_1110_));
 INV_X1 _1894_ (.A(\transfer_count[2][9] ),
    .ZN(_1111_));
 CLKBUF_X2 _1895_ (.A(\transfer_count[2][8] ),
    .Z(_1112_));
 INV_X1 _1896_ (.A(_1112_),
    .ZN(_1113_));
 NAND4_X4 _1897_ (.A1(_1098_),
    .A2(\transfer_count[2][6] ),
    .A3(_1097_),
    .A4(_1099_),
    .ZN(_1114_));
 OR4_X1 _1898_ (.A1(_1110_),
    .A2(_1111_),
    .A3(_1113_),
    .A4(_1114_),
    .ZN(_1115_));
 OR4_X1 _1899_ (.A1(_1106_),
    .A2(_1107_),
    .A3(_1109_),
    .A4(_1115_),
    .ZN(_1116_));
 XNOR2_X1 _1900_ (.A(_1104_),
    .B(_1116_),
    .ZN(_1498_));
 NOR3_X2 _1901_ (.A1(_1113_),
    .A2(_1109_),
    .A3(_1114_),
    .ZN(_1117_));
 XNOR2_X2 _1902_ (.A(\transfer_count[2][9] ),
    .B(_1117_),
    .ZN(_1510_));
 BUF_X1 _1903_ (.A(\transfer_count[2][29] ),
    .Z(_1118_));
 NAND4_X1 _1904_ (.A1(\transfer_count[2][11] ),
    .A2(\transfer_count[2][10] ),
    .A3(\transfer_count[2][9] ),
    .A4(_1112_),
    .ZN(_1119_));
 OR3_X4 _1905_ (.A1(_1109_),
    .A2(_1114_),
    .A3(_1119_),
    .ZN(_1120_));
 CLKBUF_X2 _1906_ (.A(\transfer_count[2][28] ),
    .Z(_1121_));
 CLKBUF_X2 _1907_ (.A(\transfer_count[2][27] ),
    .Z(_1122_));
 BUF_X2 _1908_ (.A(\transfer_count[2][26] ),
    .Z(_1123_));
 NAND3_X1 _1909_ (.A1(_1121_),
    .A2(_1122_),
    .A3(_1123_),
    .ZN(_1124_));
 BUF_X2 _1910_ (.A(\transfer_count[2][24] ),
    .Z(_1125_));
 BUF_X2 _1911_ (.A(\transfer_count[2][21] ),
    .Z(_1126_));
 CLKBUF_X3 _1912_ (.A(\transfer_count[2][20] ),
    .Z(_1127_));
 AND4_X2 _1913_ (.A1(\transfer_count[2][23] ),
    .A2(\transfer_count[2][22] ),
    .A3(_1126_),
    .A4(_1127_),
    .ZN(_1128_));
 NAND3_X4 _1914_ (.A1(\transfer_count[2][25] ),
    .A2(_1125_),
    .A3(_1128_),
    .ZN(_1129_));
 BUF_X2 _1915_ (.A(\transfer_count[2][16] ),
    .Z(_1130_));
 BUF_X1 _1916_ (.A(\transfer_count[2][14] ),
    .Z(_1131_));
 AND4_X1 _1917_ (.A1(_1131_),
    .A2(\transfer_count[2][13] ),
    .A3(_1105_),
    .A4(\transfer_count[2][15] ),
    .ZN(_1132_));
 BUF_X1 _1918_ (.A(\transfer_count[2][18] ),
    .Z(_1133_));
 BUF_X1 _1919_ (.A(\transfer_count[2][17] ),
    .Z(_1134_));
 AND3_X1 _1920_ (.A1(\transfer_count[2][19] ),
    .A2(_1133_),
    .A3(_1134_),
    .ZN(_1135_));
 NAND3_X4 _1921_ (.A1(_1130_),
    .A2(_1132_),
    .A3(_1135_),
    .ZN(_1136_));
 NOR4_X2 _1922_ (.A1(_1120_),
    .A2(_1124_),
    .A3(_1129_),
    .A4(_1136_),
    .ZN(_1137_));
 XNOR2_X1 _1923_ (.A(_1118_),
    .B(_1137_),
    .ZN(_1522_));
 INV_X1 _1924_ (.A(\transfer_count[2][25] ),
    .ZN(_1138_));
 AND2_X1 _1925_ (.A1(_1125_),
    .A2(_1128_),
    .ZN(_1139_));
 NOR2_X4 _1926_ (.A1(_1120_),
    .A2(_1136_),
    .ZN(_1140_));
 NAND2_X1 _1927_ (.A1(_1139_),
    .A2(_1140_),
    .ZN(_1141_));
 XNOR2_X1 _1928_ (.A(_1138_),
    .B(_1141_),
    .ZN(_1534_));
 NAND2_X1 _1929_ (.A1(_1127_),
    .A2(_1140_),
    .ZN(_1142_));
 XOR2_X2 _1930_ (.A(_1126_),
    .B(_1142_),
    .Z(_1546_));
 NAND2_X1 _1931_ (.A1(_1130_),
    .A2(_1132_),
    .ZN(_1143_));
 NOR2_X2 _1932_ (.A1(_1120_),
    .A2(_1143_),
    .ZN(_1144_));
 XNOR2_X1 _1933_ (.A(_1134_),
    .B(_1144_),
    .ZN(_1558_));
 NAND4_X2 _1934_ (.A1(_1518_),
    .A2(_1524_),
    .A3(_1521_),
    .A4(_1527_),
    .ZN(_1145_));
 NAND4_X1 _1935_ (.A1(_1530_),
    .A2(_1536_),
    .A3(_1533_),
    .A4(_1539_),
    .ZN(_1146_));
 NAND4_X2 _1936_ (.A1(_1542_),
    .A2(_1548_),
    .A3(_1545_),
    .A4(_1551_),
    .ZN(_1147_));
 NOR3_X1 _1937_ (.A1(_1145_),
    .A2(_1146_),
    .A3(_1147_),
    .ZN(_1148_));
 AOI21_X1 _1938_ (.A(_1553_),
    .B1(_1556_),
    .B2(_1554_),
    .ZN(_1149_));
 AOI21_X1 _1939_ (.A(_1559_),
    .B1(_1562_),
    .B2(_1560_),
    .ZN(_1150_));
 NAND2_X1 _1940_ (.A1(_1554_),
    .A2(_1557_),
    .ZN(_1151_));
 OAI21_X1 _1941_ (.A(_1149_),
    .B1(_1150_),
    .B2(_1151_),
    .ZN(_1152_));
 NAND3_X1 _1942_ (.A1(_1524_),
    .A2(_1521_),
    .A3(_1526_),
    .ZN(_1153_));
 AOI21_X1 _1943_ (.A(_1520_),
    .B1(_1523_),
    .B2(_1521_),
    .ZN(_1154_));
 NAND2_X1 _1944_ (.A1(_1153_),
    .A2(_1154_),
    .ZN(_1155_));
 AOI221_X2 _1945_ (.A(_1517_),
    .B1(_1148_),
    .B2(_1152_),
    .C1(_1155_),
    .C2(_1518_),
    .ZN(_1156_));
 AND2_X1 _1946_ (.A1(_1542_),
    .A2(_1545_),
    .ZN(_1157_));
 AOI21_X1 _1947_ (.A(_1547_),
    .B1(_1550_),
    .B2(_1548_),
    .ZN(_1158_));
 INV_X1 _1948_ (.A(_1158_),
    .ZN(_1159_));
 AOI221_X2 _1949_ (.A(_1541_),
    .B1(_1157_),
    .B2(_1159_),
    .C1(_1544_),
    .C2(_1542_),
    .ZN(_1160_));
 OR2_X2 _1950_ (.A1(_1145_),
    .A2(_1146_),
    .ZN(_1161_));
 INV_X1 _1951_ (.A(_1532_),
    .ZN(_1162_));
 AOI21_X1 _1952_ (.A(_1535_),
    .B1(_1538_),
    .B2(_1536_),
    .ZN(_1163_));
 INV_X1 _1953_ (.A(_1533_),
    .ZN(_1164_));
 OAI21_X1 _1954_ (.A(_1162_),
    .B1(_1163_),
    .B2(_1164_),
    .ZN(_1165_));
 AOI21_X1 _1955_ (.A(_1529_),
    .B1(_1165_),
    .B2(_1530_),
    .ZN(_1166_));
 OAI221_X2 _1956_ (.A(_1156_),
    .B1(_1160_),
    .B2(_1161_),
    .C1(_1145_),
    .C2(_1166_),
    .ZN(_1167_));
 AND2_X1 _1957_ (.A1(_1476_),
    .A2(_1479_),
    .ZN(_1168_));
 NAND4_X4 _1958_ (.A1(_1506_),
    .A2(_1512_),
    .A3(_1509_),
    .A4(_1515_),
    .ZN(_1169_));
 NAND4_X4 _1959_ (.A1(_1494_),
    .A2(_1500_),
    .A3(_1497_),
    .A4(_1503_),
    .ZN(_1170_));
 NAND2_X2 _1960_ (.A1(_1482_),
    .A2(_1485_),
    .ZN(_1171_));
 NAND2_X2 _1961_ (.A1(_1488_),
    .A2(_1491_),
    .ZN(_1172_));
 NOR4_X4 _1962_ (.A1(_1169_),
    .A2(_1170_),
    .A3(_1171_),
    .A4(_1172_),
    .ZN(_1173_));
 NAND2_X1 _1963_ (.A1(_1560_),
    .A2(_1563_),
    .ZN(_1174_));
 NOR4_X4 _1964_ (.A1(_1161_),
    .A2(_1147_),
    .A3(_1151_),
    .A4(_1174_),
    .ZN(_1175_));
 AND2_X1 _1965_ (.A1(_1473_),
    .A2(_1468_),
    .ZN(_1176_));
 NAND4_X4 _1966_ (.A1(_1168_),
    .A2(_1173_),
    .A3(_1175_),
    .A4(_1176_),
    .ZN(_1177_));
 INV_X8 _1967_ (.A(_1087_),
    .ZN(_1178_));
 CLKBUF_X3 _1968_ (.A(\channel_state[2][1] ),
    .Z(_1179_));
 NAND2_X4 _1969_ (.A1(net132),
    .A2(_1179_),
    .ZN(_1180_));
 NOR2_X4 _1970_ (.A1(_1178_),
    .A2(_1180_),
    .ZN(_1181_));
 NAND3_X1 _1971_ (.A1(_1167_),
    .A2(_1177_),
    .A3(_1181_),
    .ZN(_1182_));
 NAND2_X1 _1972_ (.A1(_1177_),
    .A2(_1181_),
    .ZN(_1183_));
 NOR2_X1 _1973_ (.A1(_1169_),
    .A2(_1170_),
    .ZN(_1184_));
 AOI21_X1 _1974_ (.A(_1481_),
    .B1(_1484_),
    .B2(_1482_),
    .ZN(_1185_));
 AOI21_X1 _1975_ (.A(_1487_),
    .B1(_1490_),
    .B2(_1488_),
    .ZN(_1186_));
 OAI21_X1 _1976_ (.A(_1185_),
    .B1(_1171_),
    .B2(_1186_),
    .ZN(_1187_));
 NAND3_X1 _1977_ (.A1(_1500_),
    .A2(_1497_),
    .A3(_1502_),
    .ZN(_1188_));
 AOI21_X1 _1978_ (.A(_1496_),
    .B1(_1499_),
    .B2(_1497_),
    .ZN(_1189_));
 NAND2_X1 _1979_ (.A1(_1188_),
    .A2(_1189_),
    .ZN(_1190_));
 AOI221_X2 _1980_ (.A(_1493_),
    .B1(_1184_),
    .B2(_1187_),
    .C1(_1190_),
    .C2(_1494_),
    .ZN(_1191_));
 INV_X1 _1981_ (.A(_1170_),
    .ZN(_1192_));
 AOI21_X1 _1982_ (.A(_1505_),
    .B1(_1508_),
    .B2(_1506_),
    .ZN(_1193_));
 NAND2_X1 _1983_ (.A1(_1506_),
    .A2(_1509_),
    .ZN(_1194_));
 AOI21_X1 _1984_ (.A(_1511_),
    .B1(_1514_),
    .B2(_1512_),
    .ZN(_1195_));
 OAI21_X1 _1985_ (.A(_1193_),
    .B1(_1194_),
    .B2(_1195_),
    .ZN(_1196_));
 NAND2_X1 _1986_ (.A1(_1192_),
    .A2(_1196_),
    .ZN(_1197_));
 INV_X1 _1987_ (.A(_1472_),
    .ZN(_1198_));
 INV_X1 _1988_ (.A(_1473_),
    .ZN(_1199_));
 OAI21_X1 _1989_ (.A(_1198_),
    .B1(_1467_),
    .B2(_1199_),
    .ZN(_1200_));
 AOI221_X2 _1990_ (.A(_1475_),
    .B1(_1200_),
    .B2(_1168_),
    .C1(_1478_),
    .C2(_1476_),
    .ZN(_1201_));
 OR4_X2 _1991_ (.A1(_1169_),
    .A2(_1170_),
    .A3(_1171_),
    .A4(_1172_),
    .ZN(_1202_));
 OAI211_X4 _1992_ (.A(_1191_),
    .B(_1197_),
    .C1(_1201_),
    .C2(_1202_),
    .ZN(_1203_));
 NAND2_X1 _1993_ (.A1(_1203_),
    .A2(_1175_),
    .ZN(_1204_));
 BUF_X8 _1994_ (.A(_1178_),
    .Z(_1205_));
 BUF_X4 _1995_ (.A(_1205_),
    .Z(_1206_));
 NAND3_X4 _1996_ (.A1(net129),
    .A2(_1091_),
    .A3(_1094_),
    .ZN(_1207_));
 OAI221_X1 _1997_ (.A(_1182_),
    .B1(_1183_),
    .B2(_1204_),
    .C1(_1206_),
    .C2(_1207_),
    .ZN(_0017_));
 CLKBUF_X2 _1998_ (.A(\transfer_count[1][28] ),
    .Z(_1208_));
 BUF_X2 _1999_ (.A(\transfer_count[1][27] ),
    .Z(_1209_));
 BUF_X1 _2000_ (.A(\transfer_count[1][26] ),
    .Z(_1210_));
 CLKBUF_X2 _2001_ (.A(\transfer_count[1][25] ),
    .Z(_1211_));
 BUF_X2 _2002_ (.A(\transfer_count[1][24] ),
    .Z(_1212_));
 BUF_X2 _2003_ (.A(\transfer_count[1][23] ),
    .Z(_1213_));
 AND4_X2 _2004_ (.A1(_1210_),
    .A2(_1211_),
    .A3(_1212_),
    .A4(_1213_),
    .ZN(_1214_));
 NAND3_X1 _2005_ (.A1(_1208_),
    .A2(_1209_),
    .A3(_1214_),
    .ZN(_1215_));
 BUF_X2 _2006_ (.A(\transfer_count[1][22] ),
    .Z(_1216_));
 CLKBUF_X3 _2007_ (.A(\transfer_count[1][21] ),
    .Z(_1217_));
 NAND2_X4 _2008_ (.A1(_1216_),
    .A2(_1217_),
    .ZN(_1218_));
 BUF_X2 _2009_ (.A(\transfer_count[1][20] ),
    .Z(_1219_));
 BUF_X2 _2010_ (.A(\transfer_count[1][16] ),
    .Z(_1220_));
 BUF_X2 _2011_ (.A(\transfer_count[1][15] ),
    .Z(_1221_));
 BUF_X4 _2012_ (.A(\transfer_count[1][14] ),
    .Z(_1222_));
 AND4_X2 _2013_ (.A1(\transfer_count[1][17] ),
    .A2(_1220_),
    .A3(_1221_),
    .A4(_1222_),
    .ZN(_1223_));
 BUF_X2 _2014_ (.A(\transfer_count[1][18] ),
    .Z(_1224_));
 AND2_X2 _2015_ (.A1(\transfer_count[1][19] ),
    .A2(_1224_),
    .ZN(_1225_));
 NAND3_X4 _2016_ (.A1(_1219_),
    .A2(_1223_),
    .A3(_1225_),
    .ZN(_1226_));
 BUF_X2 _2017_ (.A(\transfer_count[1][6] ),
    .Z(_1227_));
 BUF_X2 _2018_ (.A(\transfer_count[1][5] ),
    .Z(_1228_));
 BUF_X2 _2019_ (.A(\transfer_count[1][4] ),
    .Z(_1229_));
 NAND3_X4 _2020_ (.A1(_1227_),
    .A2(_1228_),
    .A3(_1229_),
    .ZN(_1230_));
 CLKBUF_X3 _2021_ (.A(\transfer_count[1][3] ),
    .Z(_1231_));
 CLKBUF_X3 _2022_ (.A(\transfer_count[1][2] ),
    .Z(_1232_));
 NAND4_X4 _2023_ (.A1(_1231_),
    .A2(_1232_),
    .A3(\transfer_count[1][1] ),
    .A4(\transfer_count[1][0] ),
    .ZN(_1233_));
 OR2_X2 _2024_ (.A1(_1230_),
    .A2(_1233_),
    .ZN(_1234_));
 BUF_X4 _2025_ (.A(\transfer_count[1][8] ),
    .Z(_1235_));
 BUF_X4 _2026_ (.A(\transfer_count[1][7] ),
    .Z(_1236_));
 NAND4_X4 _2027_ (.A1(\transfer_count[1][10] ),
    .A2(\transfer_count[1][9] ),
    .A3(_1235_),
    .A4(_1236_),
    .ZN(_1237_));
 BUF_X2 _2028_ (.A(\transfer_count[1][12] ),
    .Z(_1238_));
 CLKBUF_X3 _2029_ (.A(\transfer_count[1][11] ),
    .Z(_1239_));
 NAND3_X4 _2030_ (.A1(\transfer_count[1][13] ),
    .A2(_1238_),
    .A3(_1239_),
    .ZN(_1240_));
 OR2_X2 _2031_ (.A1(_1237_),
    .A2(_1240_),
    .ZN(_1241_));
 OR3_X4 _2032_ (.A1(_1226_),
    .A2(_1234_),
    .A3(_1241_),
    .ZN(_1242_));
 NOR3_X2 _2033_ (.A1(_1215_),
    .A2(_1218_),
    .A3(_1242_),
    .ZN(_1243_));
 XNOR2_X2 _2034_ (.A(\transfer_count[1][29] ),
    .B(_1243_),
    .ZN(_1570_));
 NOR4_X4 _2035_ (.A1(_1218_),
    .A2(_1226_),
    .A3(_1234_),
    .A4(_1241_),
    .ZN(_1244_));
 NAND2_X1 _2036_ (.A1(_1214_),
    .A2(_1244_),
    .ZN(_1245_));
 XOR2_X2 _2037_ (.A(_1209_),
    .B(_1245_),
    .Z(_1576_));
 NAND2_X1 _2038_ (.A1(_1212_),
    .A2(_1213_),
    .ZN(_1246_));
 NOR3_X2 _2039_ (.A1(_1246_),
    .A2(_1218_),
    .A3(_1242_),
    .ZN(_1247_));
 XNOR2_X2 _2040_ (.A(_1211_),
    .B(_1247_),
    .ZN(_1582_));
 XNOR2_X1 _2041_ (.A(_1213_),
    .B(_1244_),
    .ZN(_1588_));
 XOR2_X2 _2042_ (.A(_1217_),
    .B(_1242_),
    .Z(_1594_));
 NAND3_X1 _2043_ (.A1(_1224_),
    .A2(\transfer_count[1][17] ),
    .A3(_1220_),
    .ZN(_1248_));
 NOR4_X4 _2044_ (.A1(_1230_),
    .A2(_1233_),
    .A3(_1237_),
    .A4(_1240_),
    .ZN(_1249_));
 NAND3_X1 _2045_ (.A1(_1221_),
    .A2(_1222_),
    .A3(_1249_),
    .ZN(_1250_));
 NOR2_X2 _2046_ (.A1(_1248_),
    .A2(_1250_),
    .ZN(_1251_));
 XNOR2_X2 _2047_ (.A(\transfer_count[1][19] ),
    .B(_1251_),
    .ZN(_1600_));
 NAND2_X1 _2048_ (.A1(_1222_),
    .A2(_1249_),
    .ZN(_1252_));
 XOR2_X2 _2049_ (.A(_1221_),
    .B(_1252_),
    .Z(_1612_));
 NOR2_X2 _2050_ (.A1(_1234_),
    .A2(_1237_),
    .ZN(_1253_));
 NAND3_X2 _2051_ (.A1(_1238_),
    .A2(_1239_),
    .A3(_1253_),
    .ZN(_1254_));
 XOR2_X2 _2052_ (.A(\transfer_count[1][13] ),
    .B(_1254_),
    .Z(_1618_));
 XNOR2_X1 _2053_ (.A(_1239_),
    .B(_1253_),
    .ZN(_1624_));
 NOR2_X2 _2054_ (.A1(_1230_),
    .A2(_1233_),
    .ZN(_1255_));
 NAND3_X1 _2055_ (.A1(_1235_),
    .A2(_1236_),
    .A3(_1255_),
    .ZN(_1256_));
 XOR2_X2 _2056_ (.A(\transfer_count[1][9] ),
    .B(_1256_),
    .Z(_1630_));
 XNOR2_X1 _2057_ (.A(_1236_),
    .B(_1255_),
    .ZN(_1636_));
 INV_X1 _2058_ (.A(_1229_),
    .ZN(_1257_));
 NOR2_X1 _2059_ (.A1(_1257_),
    .A2(_1233_),
    .ZN(_1258_));
 XNOR2_X2 _2060_ (.A(_1228_),
    .B(_1258_),
    .ZN(_1642_));
 NAND3_X2 _2061_ (.A1(_1232_),
    .A2(\transfer_count[1][1] ),
    .A3(\transfer_count[1][0] ),
    .ZN(_1259_));
 XOR2_X2 _2062_ (.A(_1231_),
    .B(_1259_),
    .Z(_1648_));
 BUF_X2 _2063_ (.A(channel_start[1]),
    .Z(_1260_));
 BUF_X2 _2064_ (.A(\channel_state[1][0] ),
    .Z(_1261_));
 BUF_X2 _2065_ (.A(channel_enable[1]),
    .Z(_1262_));
 NAND2_X1 _2066_ (.A1(_1261_),
    .A2(_1262_),
    .ZN(_1263_));
 NAND4_X1 _2067_ (.A1(_1088_),
    .A2(_1260_),
    .A3(\channel_state[1][4] ),
    .A4(_1263_),
    .ZN(_1264_));
 AND2_X1 _2068_ (.A1(net131),
    .A2(\channel_state[1][1] ),
    .ZN(_1265_));
 CLKBUF_X3 _2069_ (.A(_1265_),
    .Z(_1266_));
 NAND2_X2 _2070_ (.A1(_1087_),
    .A2(_1266_),
    .ZN(_1267_));
 CLKBUF_X3 _2071_ (.A(_1267_),
    .Z(_1268_));
 NAND4_X4 _2072_ (.A1(_1566_),
    .A2(_1569_),
    .A3(_1575_),
    .A4(_1572_),
    .ZN(_1269_));
 INV_X1 _2073_ (.A(_1269_),
    .ZN(_1270_));
 AOI21_X1 _2074_ (.A(_1577_),
    .B1(_1580_),
    .B2(_1578_),
    .ZN(_1271_));
 NAND2_X1 _2075_ (.A1(_1578_),
    .A2(_1581_),
    .ZN(_1272_));
 AOI21_X1 _2076_ (.A(_1583_),
    .B1(_1584_),
    .B2(_1586_),
    .ZN(_1273_));
 OAI21_X1 _2077_ (.A(_1271_),
    .B1(_1272_),
    .B2(_1273_),
    .ZN(_1274_));
 AOI21_X1 _2078_ (.A(_1589_),
    .B1(_1592_),
    .B2(_1590_),
    .ZN(_1275_));
 NAND2_X1 _2079_ (.A1(_1590_),
    .A2(_1593_),
    .ZN(_1276_));
 AOI21_X1 _2080_ (.A(_1595_),
    .B1(_1596_),
    .B2(_1598_),
    .ZN(_1277_));
 OAI21_X1 _2081_ (.A(_1275_),
    .B1(_1276_),
    .B2(_1277_),
    .ZN(_1278_));
 NAND4_X2 _2082_ (.A1(_1578_),
    .A2(_1581_),
    .A3(_1587_),
    .A4(_1584_),
    .ZN(_1279_));
 NOR2_X2 _2083_ (.A1(_1269_),
    .A2(_1279_),
    .ZN(_1280_));
 AOI22_X2 _2084_ (.A1(_1270_),
    .A2(_1274_),
    .B1(_1278_),
    .B2(_1280_),
    .ZN(_1281_));
 AOI21_X1 _2085_ (.A(_1565_),
    .B1(_1568_),
    .B2(_1566_),
    .ZN(_1282_));
 AOI21_X1 _2086_ (.A(_1571_),
    .B1(_1572_),
    .B2(_1574_),
    .ZN(_1283_));
 NAND2_X1 _2087_ (.A1(_1566_),
    .A2(_1569_),
    .ZN(_1284_));
 OAI21_X2 _2088_ (.A(_1282_),
    .B1(_1283_),
    .B2(_1284_),
    .ZN(_1285_));
 AOI21_X1 _2089_ (.A(_1601_),
    .B1(_1604_),
    .B2(_1602_),
    .ZN(_1286_));
 NAND2_X1 _2090_ (.A1(_1602_),
    .A2(_1605_),
    .ZN(_1287_));
 AOI21_X1 _2091_ (.A(_1607_),
    .B1(_1608_),
    .B2(_1610_),
    .ZN(_1288_));
 OAI21_X1 _2092_ (.A(_1286_),
    .B1(_1287_),
    .B2(_1288_),
    .ZN(_1289_));
 NAND4_X2 _2093_ (.A1(_1590_),
    .A2(_1593_),
    .A3(_1599_),
    .A4(_1596_),
    .ZN(_0181_));
 NOR3_X2 _2094_ (.A1(_1269_),
    .A2(_1279_),
    .A3(_0181_),
    .ZN(_0182_));
 AOI21_X1 _2095_ (.A(_1285_),
    .B1(_1289_),
    .B2(_0182_),
    .ZN(_0183_));
 NAND2_X1 _2096_ (.A1(_1281_),
    .A2(_0183_),
    .ZN(_0184_));
 NAND3_X1 _2097_ (.A1(_1622_),
    .A2(_1617_),
    .A3(_1620_),
    .ZN(_0185_));
 AOI21_X1 _2098_ (.A(_1616_),
    .B1(_1619_),
    .B2(_1617_),
    .ZN(_0186_));
 NAND2_X1 _2099_ (.A1(_0185_),
    .A2(_0186_),
    .ZN(_0187_));
 AOI21_X1 _2100_ (.A(_1613_),
    .B1(_0187_),
    .B2(_1614_),
    .ZN(_0188_));
 NAND4_X2 _2101_ (.A1(_1614_),
    .A2(_1617_),
    .A3(_1623_),
    .A4(_1620_),
    .ZN(_0189_));
 INV_X1 _2102_ (.A(_0189_),
    .ZN(_0190_));
 AOI21_X1 _2103_ (.A(_1625_),
    .B1(_1628_),
    .B2(_1626_),
    .ZN(_0191_));
 NAND2_X1 _2104_ (.A1(_1626_),
    .A2(_1629_),
    .ZN(_0192_));
 AOI21_X1 _2105_ (.A(_1631_),
    .B1(_1632_),
    .B2(_1634_),
    .ZN(_0193_));
 OAI21_X1 _2106_ (.A(_0191_),
    .B1(_0192_),
    .B2(_0193_),
    .ZN(_0194_));
 NAND4_X1 _2107_ (.A1(_1626_),
    .A2(_1629_),
    .A3(_1635_),
    .A4(_1632_),
    .ZN(_0195_));
 NOR2_X1 _2108_ (.A1(_0189_),
    .A2(_0195_),
    .ZN(_0196_));
 AOI21_X1 _2109_ (.A(_1637_),
    .B1(_1640_),
    .B2(_1638_),
    .ZN(_0197_));
 NAND2_X1 _2110_ (.A1(_1638_),
    .A2(_1641_),
    .ZN(_0198_));
 AOI21_X1 _2111_ (.A(_1643_),
    .B1(_1644_),
    .B2(_1646_),
    .ZN(_0199_));
 OAI21_X1 _2112_ (.A(_0197_),
    .B1(_0198_),
    .B2(_0199_),
    .ZN(_0200_));
 AOI22_X2 _2113_ (.A1(_0190_),
    .A2(_0194_),
    .B1(_0196_),
    .B2(_0200_),
    .ZN(_0201_));
 NAND2_X1 _2114_ (.A1(_1647_),
    .A2(_1644_),
    .ZN(_0202_));
 OR4_X1 _2115_ (.A1(_0189_),
    .A2(_0195_),
    .A3(_0198_),
    .A4(_0202_),
    .ZN(_0203_));
 INV_X1 _2116_ (.A(_1657_),
    .ZN(_0204_));
 INV_X1 _2117_ (.A(_1658_),
    .ZN(_0205_));
 OAI21_X1 _2118_ (.A(_0204_),
    .B1(_1661_),
    .B2(_0205_),
    .ZN(_0206_));
 AND2_X1 _2119_ (.A1(_1650_),
    .A2(_1653_),
    .ZN(_0207_));
 AOI221_X2 _2120_ (.A(_1649_),
    .B1(_0206_),
    .B2(_0207_),
    .C1(_1652_),
    .C2(_1650_),
    .ZN(_0208_));
 OAI211_X2 _2121_ (.A(_0188_),
    .B(_0201_),
    .C1(_0203_),
    .C2(_0208_),
    .ZN(_0209_));
 OR2_X1 _2122_ (.A1(_0184_),
    .A2(_0209_),
    .ZN(_0210_));
 NAND2_X1 _2123_ (.A1(_1608_),
    .A2(_1611_),
    .ZN(_0211_));
 NOR3_X2 _2124_ (.A1(_0181_),
    .A2(_1287_),
    .A3(_0211_),
    .ZN(_0212_));
 AOI221_X2 _2125_ (.A(_1285_),
    .B1(_0212_),
    .B2(_1280_),
    .C1(_0182_),
    .C2(_1289_),
    .ZN(_0213_));
 NAND2_X2 _2126_ (.A1(_1281_),
    .A2(_0213_),
    .ZN(_0214_));
 NAND2_X1 _2127_ (.A1(_1280_),
    .A2(_0212_),
    .ZN(_0215_));
 NAND3_X1 _2128_ (.A1(_1658_),
    .A2(_1662_),
    .A3(_0207_),
    .ZN(_0216_));
 OR3_X2 _2129_ (.A1(_0203_),
    .A2(_0215_),
    .A3(_0216_),
    .ZN(_0217_));
 AND3_X1 _2130_ (.A1(_1264_),
    .A2(_0214_),
    .A3(_0217_),
    .ZN(_0218_));
 AOI22_X1 _2131_ (.A1(_1264_),
    .A2(_1268_),
    .B1(_0210_),
    .B2(_0218_),
    .ZN(_0013_));
 BUF_X8 _2132_ (.A(_1205_),
    .Z(_0219_));
 NAND3_X4 _2133_ (.A1(_1261_),
    .A2(_1260_),
    .A3(_1262_),
    .ZN(_0220_));
 NAND2_X2 _2134_ (.A1(net131),
    .A2(\channel_state[1][1] ),
    .ZN(_0221_));
 NOR2_X2 _2135_ (.A1(_1178_),
    .A2(_0221_),
    .ZN(_0222_));
 CLKBUF_X3 _2136_ (.A(_0222_),
    .Z(_0223_));
 NAND3_X1 _2137_ (.A1(_0223_),
    .A2(_0214_),
    .A3(_0217_),
    .ZN(_0224_));
 NOR2_X1 _2138_ (.A1(_0184_),
    .A2(_0209_),
    .ZN(_0225_));
 OAI22_X1 _2139_ (.A1(_0219_),
    .A2(_0220_),
    .B1(_0224_),
    .B2(_0225_),
    .ZN(_0012_));
 CLKBUF_X2 _2140_ (.A(\transfer_count[0][29] ),
    .Z(_0226_));
 BUF_X2 _2141_ (.A(\transfer_count[0][20] ),
    .Z(_0227_));
 BUF_X2 _2142_ (.A(\transfer_count[0][19] ),
    .Z(_0228_));
 BUF_X2 _2143_ (.A(\transfer_count[0][18] ),
    .Z(_0229_));
 CLKBUF_X2 _2144_ (.A(\transfer_count[0][16] ),
    .Z(_0230_));
 CLKBUF_X2 _2145_ (.A(\transfer_count[0][14] ),
    .Z(_0231_));
 AND4_X2 _2146_ (.A1(\transfer_count[0][17] ),
    .A2(_0230_),
    .A3(\transfer_count[0][15] ),
    .A4(_0231_),
    .ZN(_0232_));
 NAND4_X4 _2147_ (.A1(_0227_),
    .A2(_0228_),
    .A3(_0229_),
    .A4(_0232_),
    .ZN(_0233_));
 BUF_X2 _2148_ (.A(\transfer_count[0][13] ),
    .Z(_0234_));
 BUF_X2 _2149_ (.A(\transfer_count[0][12] ),
    .Z(_0235_));
 CLKBUF_X3 _2150_ (.A(\transfer_count[0][11] ),
    .Z(_0236_));
 NAND3_X4 _2151_ (.A1(_0234_),
    .A2(_0235_),
    .A3(_0236_),
    .ZN(_0237_));
 BUF_X2 _2152_ (.A(\transfer_count[0][3] ),
    .Z(_0238_));
 CLKBUF_X3 _2153_ (.A(\transfer_count[0][2] ),
    .Z(_0239_));
 NAND4_X4 _2154_ (.A1(_0238_),
    .A2(_0239_),
    .A3(\transfer_count[0][1] ),
    .A4(\transfer_count[0][0] ),
    .ZN(_0240_));
 BUF_X2 _2155_ (.A(\transfer_count[0][6] ),
    .Z(_0241_));
 BUF_X2 _2156_ (.A(\transfer_count[0][5] ),
    .Z(_0242_));
 BUF_X2 _2157_ (.A(\transfer_count[0][4] ),
    .Z(_0243_));
 NAND3_X4 _2158_ (.A1(_0241_),
    .A2(_0242_),
    .A3(_0243_),
    .ZN(_0244_));
 BUF_X2 _2159_ (.A(\transfer_count[0][10] ),
    .Z(_0245_));
 BUF_X2 _2160_ (.A(\transfer_count[0][9] ),
    .Z(_0246_));
 BUF_X2 _2161_ (.A(\transfer_count[0][8] ),
    .Z(_0247_));
 CLKBUF_X3 _2162_ (.A(\transfer_count[0][7] ),
    .Z(_0248_));
 NAND4_X4 _2163_ (.A1(_0245_),
    .A2(_0246_),
    .A3(_0247_),
    .A4(_0248_),
    .ZN(_0249_));
 OR3_X4 _2164_ (.A1(_0240_),
    .A2(_0244_),
    .A3(_0249_),
    .ZN(_0250_));
 CLKBUF_X2 _2165_ (.A(\transfer_count[0][28] ),
    .Z(_0251_));
 BUF_X2 _2166_ (.A(\transfer_count[0][27] ),
    .Z(_0252_));
 CLKBUF_X2 _2167_ (.A(\transfer_count[0][25] ),
    .Z(_0253_));
 CLKBUF_X2 _2168_ (.A(\transfer_count[0][24] ),
    .Z(_0254_));
 BUF_X2 _2169_ (.A(\transfer_count[0][23] ),
    .Z(_0255_));
 AND4_X2 _2170_ (.A1(\transfer_count[0][26] ),
    .A2(_0253_),
    .A3(_0254_),
    .A4(_0255_),
    .ZN(_0256_));
 BUF_X2 _2171_ (.A(\transfer_count[0][22] ),
    .Z(_0257_));
 BUF_X2 _2172_ (.A(\transfer_count[0][21] ),
    .Z(_0258_));
 AND2_X1 _2173_ (.A1(_0257_),
    .A2(_0258_),
    .ZN(_0259_));
 NAND4_X2 _2174_ (.A1(_0251_),
    .A2(_0252_),
    .A3(_0256_),
    .A4(_0259_),
    .ZN(_0260_));
 NOR4_X4 _2175_ (.A1(_0233_),
    .A2(_0237_),
    .A3(_0250_),
    .A4(_0260_),
    .ZN(_0261_));
 XNOR2_X2 _2176_ (.A(_0226_),
    .B(_0261_),
    .ZN(_1669_));
 NAND2_X1 _2177_ (.A1(_0256_),
    .A2(_0259_),
    .ZN(_0262_));
 NOR4_X4 _2178_ (.A1(_0233_),
    .A2(_0237_),
    .A3(_0250_),
    .A4(_0262_),
    .ZN(_0263_));
 XNOR2_X2 _2179_ (.A(_0252_),
    .B(_0263_),
    .ZN(_1675_));
 NAND2_X1 _2180_ (.A1(_0254_),
    .A2(_0255_),
    .ZN(_0264_));
 NAND2_X1 _2181_ (.A1(_0257_),
    .A2(_0258_),
    .ZN(_0265_));
 OR3_X4 _2182_ (.A1(_0233_),
    .A2(_0237_),
    .A3(_0250_),
    .ZN(_0266_));
 NOR3_X2 _2183_ (.A1(_0264_),
    .A2(_0265_),
    .A3(_0266_),
    .ZN(_0267_));
 XNOR2_X2 _2184_ (.A(_0253_),
    .B(_0267_),
    .ZN(_1681_));
 NOR2_X1 _2185_ (.A1(_0265_),
    .A2(_0266_),
    .ZN(_0268_));
 XNOR2_X2 _2186_ (.A(_0255_),
    .B(_0268_),
    .ZN(_1687_));
 INV_X1 _2187_ (.A(_0258_),
    .ZN(_0269_));
 XNOR2_X2 _2188_ (.A(_0269_),
    .B(_0266_),
    .ZN(_1693_));
 NOR4_X4 _2189_ (.A1(_0237_),
    .A2(_0240_),
    .A3(_0244_),
    .A4(_0249_),
    .ZN(_0270_));
 AND3_X1 _2190_ (.A1(_0229_),
    .A2(_0232_),
    .A3(_0270_),
    .ZN(_0271_));
 XNOR2_X1 _2191_ (.A(_0228_),
    .B(_0271_),
    .ZN(_1699_));
 INV_X1 _2192_ (.A(\transfer_count[0][15] ),
    .ZN(_0272_));
 NAND2_X1 _2193_ (.A1(_0231_),
    .A2(_0270_),
    .ZN(_0273_));
 XNOR2_X2 _2194_ (.A(_0272_),
    .B(_0273_),
    .ZN(_1711_));
 NAND2_X1 _2195_ (.A1(_0235_),
    .A2(_0236_),
    .ZN(_0274_));
 NOR2_X2 _2196_ (.A1(_0274_),
    .A2(_0250_),
    .ZN(_0275_));
 XNOR2_X2 _2197_ (.A(_0234_),
    .B(_0275_),
    .ZN(_1717_));
 XOR2_X2 _2198_ (.A(_0236_),
    .B(_0250_),
    .Z(_1723_));
 NOR2_X1 _2199_ (.A1(_0240_),
    .A2(_0244_),
    .ZN(_0276_));
 AND3_X1 _2200_ (.A1(_0247_),
    .A2(_0248_),
    .A3(_0276_),
    .ZN(_0277_));
 XNOR2_X1 _2201_ (.A(_0246_),
    .B(_0277_),
    .ZN(_1729_));
 XNOR2_X2 _2202_ (.A(_0248_),
    .B(_0276_),
    .ZN(_1735_));
 INV_X1 _2203_ (.A(_0243_),
    .ZN(_0278_));
 NOR2_X1 _2204_ (.A1(_0278_),
    .A2(_0240_),
    .ZN(_0279_));
 XNOR2_X2 _2205_ (.A(_0242_),
    .B(_0279_),
    .ZN(_1741_));
 NAND3_X1 _2206_ (.A1(_0239_),
    .A2(\transfer_count[0][1] ),
    .A3(\transfer_count[0][0] ),
    .ZN(_0280_));
 XOR2_X2 _2207_ (.A(_0238_),
    .B(_0280_),
    .Z(_1747_));
 CLKBUF_X2 _2208_ (.A(\channel_state[0][0] ),
    .Z(_0281_));
 CLKBUF_X2 _2209_ (.A(channel_start[0]),
    .Z(_0282_));
 CLKBUF_X2 _2210_ (.A(channel_enable[0]),
    .Z(_0283_));
 NAND3_X2 _2211_ (.A1(_0281_),
    .A2(_0282_),
    .A3(_0283_),
    .ZN(_0284_));
 CLKBUF_X3 _2212_ (.A(_0284_),
    .Z(_0285_));
 NAND4_X2 _2213_ (.A1(_1665_),
    .A2(_1668_),
    .A3(_1674_),
    .A4(_1671_),
    .ZN(_0286_));
 INV_X1 _2214_ (.A(_0286_),
    .ZN(_0287_));
 AOI21_X1 _2215_ (.A(_1676_),
    .B1(_1679_),
    .B2(_1677_),
    .ZN(_0288_));
 NAND2_X1 _2216_ (.A1(_1677_),
    .A2(_1680_),
    .ZN(_0289_));
 AOI21_X1 _2217_ (.A(_1682_),
    .B1(_1683_),
    .B2(_1685_),
    .ZN(_0290_));
 OAI21_X1 _2218_ (.A(_0288_),
    .B1(_0289_),
    .B2(_0290_),
    .ZN(_0291_));
 AOI21_X1 _2219_ (.A(_1688_),
    .B1(_1691_),
    .B2(_1689_),
    .ZN(_0292_));
 NAND2_X1 _2220_ (.A1(_1689_),
    .A2(_1692_),
    .ZN(_0293_));
 AOI21_X1 _2221_ (.A(_1694_),
    .B1(_1695_),
    .B2(_1697_),
    .ZN(_0294_));
 OAI21_X1 _2222_ (.A(_0292_),
    .B1(_0293_),
    .B2(_0294_),
    .ZN(_0295_));
 NAND4_X2 _2223_ (.A1(_1677_),
    .A2(_1680_),
    .A3(_1686_),
    .A4(_1683_),
    .ZN(_0296_));
 NOR2_X2 _2224_ (.A1(_0286_),
    .A2(_0296_),
    .ZN(_0297_));
 AOI22_X2 _2225_ (.A1(_0287_),
    .A2(_0291_),
    .B1(_0295_),
    .B2(_0297_),
    .ZN(_0298_));
 AOI21_X1 _2226_ (.A(_1664_),
    .B1(_1667_),
    .B2(_1665_),
    .ZN(_0299_));
 AOI21_X1 _2227_ (.A(_1670_),
    .B1(_1671_),
    .B2(_1673_),
    .ZN(_0300_));
 NAND2_X1 _2228_ (.A1(_1665_),
    .A2(_1668_),
    .ZN(_0301_));
 OAI21_X1 _2229_ (.A(_0299_),
    .B1(_0300_),
    .B2(_0301_),
    .ZN(_0302_));
 AOI21_X1 _2230_ (.A(_1700_),
    .B1(_1703_),
    .B2(_1701_),
    .ZN(_0303_));
 NAND2_X1 _2231_ (.A1(_1701_),
    .A2(_1704_),
    .ZN(_0304_));
 AOI21_X1 _2232_ (.A(_1706_),
    .B1(_1707_),
    .B2(_1709_),
    .ZN(_0305_));
 OAI21_X1 _2233_ (.A(_0303_),
    .B1(_0304_),
    .B2(_0305_),
    .ZN(_0306_));
 NAND4_X2 _2234_ (.A1(_1689_),
    .A2(_1692_),
    .A3(_1698_),
    .A4(_1695_),
    .ZN(_0307_));
 NOR3_X2 _2235_ (.A1(_0286_),
    .A2(_0296_),
    .A3(_0307_),
    .ZN(_0308_));
 AOI21_X1 _2236_ (.A(_0302_),
    .B1(_0306_),
    .B2(_0308_),
    .ZN(_0309_));
 NAND2_X1 _2237_ (.A1(_0298_),
    .A2(_0309_),
    .ZN(_0310_));
 NAND3_X1 _2238_ (.A1(_1721_),
    .A2(_1716_),
    .A3(_1719_),
    .ZN(_0311_));
 AOI21_X1 _2239_ (.A(_1715_),
    .B1(_1718_),
    .B2(_1716_),
    .ZN(_0312_));
 NAND2_X1 _2240_ (.A1(_0311_),
    .A2(_0312_),
    .ZN(_0313_));
 AOI21_X2 _2241_ (.A(_1712_),
    .B1(_0313_),
    .B2(_1713_),
    .ZN(_0314_));
 NAND4_X2 _2242_ (.A1(_1713_),
    .A2(_1716_),
    .A3(_1722_),
    .A4(_1719_),
    .ZN(_0315_));
 INV_X1 _2243_ (.A(_0315_),
    .ZN(_0316_));
 AOI21_X1 _2244_ (.A(_1724_),
    .B1(_1727_),
    .B2(_1725_),
    .ZN(_0317_));
 NAND2_X1 _2245_ (.A1(_1725_),
    .A2(_1728_),
    .ZN(_0318_));
 AOI21_X1 _2246_ (.A(_1730_),
    .B1(_1731_),
    .B2(_1733_),
    .ZN(_0319_));
 OAI21_X2 _2247_ (.A(_0317_),
    .B1(_0318_),
    .B2(_0319_),
    .ZN(_0320_));
 NAND4_X2 _2248_ (.A1(_1725_),
    .A2(_1728_),
    .A3(_1734_),
    .A4(_1731_),
    .ZN(_0321_));
 NOR2_X1 _2249_ (.A1(_0315_),
    .A2(_0321_),
    .ZN(_0322_));
 AOI21_X1 _2250_ (.A(_1736_),
    .B1(_1739_),
    .B2(_1737_),
    .ZN(_0323_));
 NAND2_X1 _2251_ (.A1(_1737_),
    .A2(_1740_),
    .ZN(_0324_));
 AOI21_X1 _2252_ (.A(_1742_),
    .B1(_1743_),
    .B2(_1745_),
    .ZN(_0325_));
 OAI21_X2 _2253_ (.A(_0323_),
    .B1(_0324_),
    .B2(_0325_),
    .ZN(_0326_));
 AOI22_X4 _2254_ (.A1(_0316_),
    .A2(_0320_),
    .B1(_0322_),
    .B2(_0326_),
    .ZN(_0327_));
 NAND4_X2 _2255_ (.A1(_1737_),
    .A2(_1740_),
    .A3(_1746_),
    .A4(_1743_),
    .ZN(_0328_));
 OR3_X1 _2256_ (.A1(_0315_),
    .A2(_0321_),
    .A3(_0328_),
    .ZN(_0329_));
 INV_X1 _2257_ (.A(_1756_),
    .ZN(_0330_));
 INV_X1 _2258_ (.A(_1757_),
    .ZN(_0331_));
 OAI21_X1 _2259_ (.A(_0330_),
    .B1(_1760_),
    .B2(_0331_),
    .ZN(_0332_));
 AND2_X1 _2260_ (.A1(_1749_),
    .A2(_1752_),
    .ZN(_0333_));
 AOI221_X2 _2261_ (.A(_1748_),
    .B1(_0332_),
    .B2(_0333_),
    .C1(_1751_),
    .C2(_1749_),
    .ZN(_0334_));
 OAI211_X4 _2262_ (.A(_0314_),
    .B(_0327_),
    .C1(_0329_),
    .C2(_0334_),
    .ZN(_0335_));
 NOR2_X1 _2263_ (.A1(_0310_),
    .A2(_0335_),
    .ZN(_0336_));
 CLKBUF_X2 _2264_ (.A(\channel_state[0][1] ),
    .Z(_0337_));
 NAND2_X4 _2265_ (.A1(_0337_),
    .A2(net130),
    .ZN(_0338_));
 NOR2_X1 _2266_ (.A1(_1178_),
    .A2(_0338_),
    .ZN(_0339_));
 CLKBUF_X3 _2267_ (.A(_0339_),
    .Z(_0340_));
 NAND2_X1 _2268_ (.A1(_1707_),
    .A2(_1710_),
    .ZN(_0341_));
 NOR3_X2 _2269_ (.A1(_0307_),
    .A2(_0304_),
    .A3(_0341_),
    .ZN(_0342_));
 AOI221_X2 _2270_ (.A(_0302_),
    .B1(_0342_),
    .B2(_0297_),
    .C1(_0308_),
    .C2(_0306_),
    .ZN(_0343_));
 NAND2_X2 _2271_ (.A1(_0298_),
    .A2(_0343_),
    .ZN(_0344_));
 NOR3_X2 _2272_ (.A1(_0315_),
    .A2(_0321_),
    .A3(_0328_),
    .ZN(_0345_));
 AND3_X1 _2273_ (.A1(_1757_),
    .A2(_1761_),
    .A3(_0333_),
    .ZN(_0346_));
 NAND4_X2 _2274_ (.A1(_0297_),
    .A2(_0345_),
    .A3(_0342_),
    .A4(_0346_),
    .ZN(_0347_));
 NAND3_X1 _2275_ (.A1(_0340_),
    .A2(_0344_),
    .A3(_0347_),
    .ZN(_0348_));
 OAI22_X1 _2276_ (.A1(_0219_),
    .A2(_0285_),
    .B1(_0336_),
    .B2(_0348_),
    .ZN(_0007_));
 BUF_X4 _2277_ (.A(_1206_),
    .Z(_0349_));
 INV_X1 _2278_ (.A(\channel_state[0][2] ),
    .ZN(_0350_));
 NOR2_X1 _2279_ (.A1(_0350_),
    .A2(net134),
    .ZN(_0351_));
 AOI21_X1 _2280_ (.A(\channel_state[0][3] ),
    .B1(_0285_),
    .B2(_0351_),
    .ZN(_0352_));
 NOR2_X1 _2281_ (.A1(_0349_),
    .A2(_0352_),
    .ZN(_0006_));
 AND2_X1 _2282_ (.A1(_1089_),
    .A2(\channel_state[2][3] ),
    .ZN(_0047_));
 AND3_X4 _2283_ (.A1(net129),
    .A2(_1091_),
    .A3(_1094_),
    .ZN(_0353_));
 NOR2_X4 _2284_ (.A1(_1178_),
    .A2(_0353_),
    .ZN(_0354_));
 INV_X1 _2285_ (.A(\channel_state[2][2] ),
    .ZN(_0355_));
 NOR2_X1 _2286_ (.A1(net136),
    .A2(_0355_),
    .ZN(_0356_));
 AOI21_X1 _2287_ (.A(_0047_),
    .B1(_0354_),
    .B2(_0356_),
    .ZN(_0357_));
 INV_X1 _2288_ (.A(_0357_),
    .ZN(_0016_));
 AND2_X1 _2289_ (.A1(_1088_),
    .A2(\channel_state[1][3] ),
    .ZN(_0046_));
 AND3_X2 _2290_ (.A1(_1261_),
    .A2(_1260_),
    .A3(_1262_),
    .ZN(_0358_));
 NOR2_X4 _2291_ (.A1(_1178_),
    .A2(_0358_),
    .ZN(_0359_));
 INV_X1 _2292_ (.A(\channel_state[1][2] ),
    .ZN(_0360_));
 NOR2_X1 _2293_ (.A1(_0360_),
    .A2(net135),
    .ZN(_0361_));
 AOI21_X1 _2294_ (.A(_0046_),
    .B1(_0359_),
    .B2(_0361_),
    .ZN(_0362_));
 INV_X1 _2295_ (.A(_0362_),
    .ZN(_0011_));
 NAND2_X1 _2296_ (.A1(_0281_),
    .A2(_0283_),
    .ZN(_0363_));
 NAND4_X1 _2297_ (.A1(_1087_),
    .A2(\channel_state[0][4] ),
    .A3(_0282_),
    .A4(_0363_),
    .ZN(_0364_));
 AND2_X1 _2298_ (.A1(_0347_),
    .A2(_0364_),
    .ZN(_0365_));
 OAI211_X2 _2299_ (.A(_0344_),
    .B(_0365_),
    .C1(_0310_),
    .C2(_0335_),
    .ZN(_0366_));
 AND2_X1 _2300_ (.A1(_0337_),
    .A2(net130),
    .ZN(_0367_));
 BUF_X4 _2301_ (.A(_0367_),
    .Z(_0368_));
 NAND2_X1 _2302_ (.A1(_1087_),
    .A2(_0368_),
    .ZN(_0369_));
 CLKBUF_X3 _2303_ (.A(_0369_),
    .Z(_0370_));
 NAND2_X1 _2304_ (.A1(_0370_),
    .A2(_0364_),
    .ZN(_0371_));
 AND2_X1 _2305_ (.A1(_0366_),
    .A2(_0371_),
    .ZN(_0008_));
 BUF_X4 _2306_ (.A(_1089_),
    .Z(_0372_));
 INV_X1 _2307_ (.A(_0337_),
    .ZN(_0373_));
 AND3_X2 _2308_ (.A1(_0281_),
    .A2(_0282_),
    .A3(_0283_),
    .ZN(_0374_));
 NOR3_X1 _2309_ (.A1(_0373_),
    .A2(net130),
    .A3(_0374_),
    .ZN(_0375_));
 OAI21_X1 _2310_ (.A(_0372_),
    .B1(\channel_state[0][5] ),
    .B2(_0375_),
    .ZN(_0376_));
 INV_X1 _2311_ (.A(_0376_),
    .ZN(_0005_));
 INV_X1 _2312_ (.A(_1179_),
    .ZN(_0377_));
 NOR3_X1 _2313_ (.A1(net132),
    .A2(_0377_),
    .A3(_0353_),
    .ZN(_0378_));
 OAI21_X1 _2314_ (.A(_0372_),
    .B1(\channel_state[2][5] ),
    .B2(_0378_),
    .ZN(_0379_));
 INV_X1 _2315_ (.A(_0379_),
    .ZN(_0015_));
 BUF_X4 _2316_ (.A(_1089_),
    .Z(_0380_));
 INV_X1 _2317_ (.A(\channel_state[1][1] ),
    .ZN(_0381_));
 NOR3_X1 _2318_ (.A1(net131),
    .A2(_0381_),
    .A3(_0358_),
    .ZN(_0382_));
 OAI21_X1 _2319_ (.A(_0380_),
    .B1(\channel_state[1][5] ),
    .B2(_0382_),
    .ZN(_0383_));
 INV_X1 _2320_ (.A(_0383_),
    .ZN(_0010_));
 AND2_X1 _2321_ (.A1(_0282_),
    .A2(_0283_),
    .ZN(_0384_));
 INV_X1 _2322_ (.A(_0282_),
    .ZN(_0385_));
 AOI21_X1 _2323_ (.A(_0281_),
    .B1(\channel_state[0][4] ),
    .B2(_0385_),
    .ZN(_0386_));
 OAI21_X1 _2324_ (.A(_1090_),
    .B1(_0384_),
    .B2(_0386_),
    .ZN(_0004_));
 AND2_X1 _2325_ (.A1(_1260_),
    .A2(_1262_),
    .ZN(_0387_));
 INV_X1 _2326_ (.A(_1260_),
    .ZN(_0388_));
 AOI21_X1 _2327_ (.A(_1261_),
    .B1(_0388_),
    .B2(\channel_state[1][4] ),
    .ZN(_0389_));
 OAI21_X1 _2328_ (.A(_1090_),
    .B1(_0387_),
    .B2(_0389_),
    .ZN(_0009_));
 BUF_X2 _2329_ (.A(\transfer_count[3][5] ),
    .Z(_0390_));
 BUF_X2 _2330_ (.A(\transfer_count[3][3] ),
    .Z(_0391_));
 BUF_X2 _2331_ (.A(\transfer_count[3][4] ),
    .Z(_0392_));
 BUF_X2 _2332_ (.A(\transfer_count[3][2] ),
    .Z(_0393_));
 AND3_X1 _2333_ (.A1(_0393_),
    .A2(\transfer_count[3][1] ),
    .A3(\transfer_count[3][0] ),
    .ZN(_0394_));
 BUF_X2 _2334_ (.A(_0394_),
    .Z(_0395_));
 NAND3_X1 _2335_ (.A1(_0391_),
    .A2(_0392_),
    .A3(_0395_),
    .ZN(_0396_));
 XOR2_X2 _2336_ (.A(_0390_),
    .B(_0396_),
    .Z(_1783_));
 BUF_X2 _2337_ (.A(\transfer_count[3][13] ),
    .Z(_0397_));
 CLKBUF_X2 _2338_ (.A(\transfer_count[3][11] ),
    .Z(_0398_));
 BUF_X2 _2339_ (.A(\transfer_count[3][10] ),
    .Z(_0399_));
 BUF_X4 _2340_ (.A(\transfer_count[3][9] ),
    .Z(_0400_));
 AND4_X2 _2341_ (.A1(\transfer_count[3][12] ),
    .A2(_0398_),
    .A3(_0399_),
    .A4(_0400_),
    .ZN(_0401_));
 BUF_X4 _2342_ (.A(\transfer_count[3][7] ),
    .Z(_0402_));
 CLKBUF_X3 _2343_ (.A(\transfer_count[3][8] ),
    .Z(_0403_));
 AND4_X4 _2344_ (.A1(_0391_),
    .A2(\transfer_count[3][6] ),
    .A3(_0390_),
    .A4(_0392_),
    .ZN(_0404_));
 AND4_X1 _2345_ (.A1(_0402_),
    .A2(_0403_),
    .A3(_0395_),
    .A4(_0404_),
    .ZN(_0405_));
 CLKBUF_X3 _2346_ (.A(_0405_),
    .Z(_0406_));
 NAND2_X1 _2347_ (.A1(_0401_),
    .A2(_0406_),
    .ZN(_0407_));
 XOR2_X2 _2348_ (.A(_0397_),
    .B(_0407_),
    .Z(_1795_));
 XNOR2_X1 _2349_ (.A(_0400_),
    .B(_0406_),
    .ZN(_1807_));
 BUF_X2 _2350_ (.A(\transfer_count[3][23] ),
    .Z(_0408_));
 AND2_X1 _2351_ (.A1(\transfer_count[3][24] ),
    .A2(_0408_),
    .ZN(_0409_));
 AND2_X1 _2352_ (.A1(\transfer_count[3][26] ),
    .A2(\transfer_count[3][25] ),
    .ZN(_0410_));
 AND3_X1 _2353_ (.A1(\transfer_count[3][27] ),
    .A2(_0409_),
    .A3(_0410_),
    .ZN(_0411_));
 INV_X1 _2354_ (.A(_0395_),
    .ZN(_0412_));
 NAND3_X2 _2355_ (.A1(_0402_),
    .A2(_0403_),
    .A3(_0404_),
    .ZN(_0413_));
 BUF_X2 _2356_ (.A(\transfer_count[3][22] ),
    .Z(_0414_));
 BUF_X2 _2357_ (.A(\transfer_count[3][21] ),
    .Z(_0415_));
 CLKBUF_X2 _2358_ (.A(\transfer_count[3][20] ),
    .Z(_0416_));
 BUF_X2 _2359_ (.A(\transfer_count[3][19] ),
    .Z(_0417_));
 BUF_X4 _2360_ (.A(\transfer_count[3][17] ),
    .Z(_0418_));
 AND4_X1 _2361_ (.A1(_0416_),
    .A2(_0417_),
    .A3(\transfer_count[3][18] ),
    .A4(_0418_),
    .ZN(_0419_));
 NAND3_X4 _2362_ (.A1(_0414_),
    .A2(_0415_),
    .A3(_0419_),
    .ZN(_0420_));
 BUF_X2 _2363_ (.A(\transfer_count[3][16] ),
    .Z(_0421_));
 AND3_X1 _2364_ (.A1(\transfer_count[3][14] ),
    .A2(_0397_),
    .A3(\transfer_count[3][15] ),
    .ZN(_0422_));
 NAND3_X4 _2365_ (.A1(_0421_),
    .A2(_0401_),
    .A3(_0422_),
    .ZN(_0423_));
 NOR4_X4 _2366_ (.A1(_0412_),
    .A2(_0413_),
    .A3(_0420_),
    .A4(_0423_),
    .ZN(_0424_));
 AND3_X1 _2367_ (.A1(\transfer_count[3][28] ),
    .A2(_0411_),
    .A3(_0424_),
    .ZN(_0425_));
 XNOR2_X1 _2368_ (.A(\transfer_count[3][29] ),
    .B(_0425_),
    .ZN(_1819_));
 INV_X1 _2369_ (.A(\transfer_count[3][25] ),
    .ZN(_0426_));
 NAND2_X1 _2370_ (.A1(_0409_),
    .A2(_0424_),
    .ZN(_0427_));
 XNOR2_X1 _2371_ (.A(_0426_),
    .B(_0427_),
    .ZN(_1831_));
 AND3_X1 _2372_ (.A1(_0421_),
    .A2(_0401_),
    .A3(_0422_),
    .ZN(_0428_));
 AND3_X1 _2373_ (.A1(_0406_),
    .A2(_0419_),
    .A3(_0428_),
    .ZN(_0429_));
 XNOR2_X1 _2374_ (.A(_0415_),
    .B(_0429_),
    .ZN(_1843_));
 NAND4_X4 _2375_ (.A1(_0402_),
    .A2(_0403_),
    .A3(_0395_),
    .A4(_0404_),
    .ZN(_0430_));
 NOR2_X2 _2376_ (.A1(_0430_),
    .A2(_0423_),
    .ZN(_0431_));
 XNOR2_X2 _2377_ (.A(_0418_),
    .B(_0431_),
    .ZN(_1855_));
 BUF_X2 _2378_ (.A(channel_start[3]),
    .Z(_0432_));
 NAND3_X1 _2379_ (.A1(_1088_),
    .A2(\channel_state[3][4] ),
    .A3(_0432_),
    .ZN(_0433_));
 BUF_X2 _2380_ (.A(channel_enable[3]),
    .Z(_0434_));
 BUF_X2 _2381_ (.A(\channel_state[3][0] ),
    .Z(_0435_));
 AOI21_X1 _2382_ (.A(_0433_),
    .B1(_0434_),
    .B2(_0435_),
    .ZN(_0436_));
 BUF_X2 _2383_ (.A(\channel_state[3][1] ),
    .Z(_0437_));
 NAND2_X4 _2384_ (.A1(_0437_),
    .A2(net133),
    .ZN(_0438_));
 NOR2_X4 _2385_ (.A1(_1178_),
    .A2(_0438_),
    .ZN(_0439_));
 AOI21_X1 _2386_ (.A(_1850_),
    .B1(_1853_),
    .B2(_1851_),
    .ZN(_0440_));
 NAND2_X1 _2387_ (.A1(_1851_),
    .A2(_1854_),
    .ZN(_0441_));
 AOI21_X1 _2388_ (.A(_1856_),
    .B1(_1859_),
    .B2(_1857_),
    .ZN(_0442_));
 OAI21_X1 _2389_ (.A(_0440_),
    .B1(_0441_),
    .B2(_0442_),
    .ZN(_0443_));
 NAND4_X4 _2390_ (.A1(_1815_),
    .A2(_1821_),
    .A3(_1818_),
    .A4(_1824_),
    .ZN(_0444_));
 NAND4_X4 _2391_ (.A1(_1827_),
    .A2(_1833_),
    .A3(_1830_),
    .A4(_1836_),
    .ZN(_0445_));
 NAND4_X2 _2392_ (.A1(_1839_),
    .A2(_1845_),
    .A3(_1842_),
    .A4(_1848_),
    .ZN(_0446_));
 NOR3_X1 _2393_ (.A1(_0444_),
    .A2(_0445_),
    .A3(_0446_),
    .ZN(_0447_));
 NAND3_X1 _2394_ (.A1(_1821_),
    .A2(_1818_),
    .A3(_1823_),
    .ZN(_0448_));
 AOI21_X1 _2395_ (.A(_1817_),
    .B1(_1820_),
    .B2(_1818_),
    .ZN(_0449_));
 NAND2_X1 _2396_ (.A1(_0448_),
    .A2(_0449_),
    .ZN(_0450_));
 AOI221_X2 _2397_ (.A(_1814_),
    .B1(_0443_),
    .B2(_0447_),
    .C1(_0450_),
    .C2(_1815_),
    .ZN(_0451_));
 INV_X1 _2398_ (.A(_0444_),
    .ZN(_0452_));
 AOI21_X1 _2399_ (.A(_1826_),
    .B1(_1829_),
    .B2(_1827_),
    .ZN(_0453_));
 NAND2_X1 _2400_ (.A1(_1827_),
    .A2(_1830_),
    .ZN(_0454_));
 AOI21_X1 _2401_ (.A(_1832_),
    .B1(_1835_),
    .B2(_1833_),
    .ZN(_0455_));
 OAI21_X1 _2402_ (.A(_0453_),
    .B1(_0454_),
    .B2(_0455_),
    .ZN(_0456_));
 NOR2_X1 _2403_ (.A1(_0444_),
    .A2(_0445_),
    .ZN(_0457_));
 AOI21_X1 _2404_ (.A(_1838_),
    .B1(_1841_),
    .B2(_1839_),
    .ZN(_0458_));
 NAND2_X1 _2405_ (.A1(_1839_),
    .A2(_1842_),
    .ZN(_0459_));
 AOI21_X1 _2406_ (.A(_1844_),
    .B1(_1847_),
    .B2(_1845_),
    .ZN(_0460_));
 OAI21_X1 _2407_ (.A(_0458_),
    .B1(_0459_),
    .B2(_0460_),
    .ZN(_0461_));
 AOI22_X2 _2408_ (.A1(_0452_),
    .A2(_0456_),
    .B1(_0457_),
    .B2(_0461_),
    .ZN(_0462_));
 NAND3_X1 _2409_ (.A1(_0439_),
    .A2(_0451_),
    .A3(_0462_),
    .ZN(_0463_));
 NAND4_X2 _2410_ (.A1(_1851_),
    .A2(_1857_),
    .A3(_1854_),
    .A4(_1860_),
    .ZN(_0464_));
 NOR4_X4 _2411_ (.A1(_0444_),
    .A2(_0445_),
    .A3(_0446_),
    .A4(_0464_),
    .ZN(_0465_));
 NAND4_X2 _2412_ (.A1(_1803_),
    .A2(_1809_),
    .A3(_1806_),
    .A4(_1812_),
    .ZN(_0466_));
 NAND4_X2 _2413_ (.A1(_1791_),
    .A2(_1797_),
    .A3(_1794_),
    .A4(_1800_),
    .ZN(_0467_));
 NOR2_X1 _2414_ (.A1(_0466_),
    .A2(_0467_),
    .ZN(_0468_));
 AOI21_X1 _2415_ (.A(_1778_),
    .B1(_1781_),
    .B2(_1779_),
    .ZN(_0469_));
 NAND2_X1 _2416_ (.A1(_1779_),
    .A2(_1782_),
    .ZN(_0470_));
 AOI21_X1 _2417_ (.A(_1784_),
    .B1(_1787_),
    .B2(_1785_),
    .ZN(_0471_));
 OAI21_X1 _2418_ (.A(_0469_),
    .B1(_0470_),
    .B2(_0471_),
    .ZN(_0472_));
 NAND3_X1 _2419_ (.A1(_1797_),
    .A2(_1794_),
    .A3(_1799_),
    .ZN(_0473_));
 AOI21_X1 _2420_ (.A(_1793_),
    .B1(_1796_),
    .B2(_1794_),
    .ZN(_0474_));
 NAND2_X1 _2421_ (.A1(_0473_),
    .A2(_0474_),
    .ZN(_0475_));
 AOI221_X2 _2422_ (.A(_1790_),
    .B1(_0468_),
    .B2(_0472_),
    .C1(_0475_),
    .C2(_1791_),
    .ZN(_0476_));
 INV_X1 _2423_ (.A(_0467_),
    .ZN(_0477_));
 AOI21_X1 _2424_ (.A(_1802_),
    .B1(_1805_),
    .B2(_1803_),
    .ZN(_0478_));
 NAND2_X1 _2425_ (.A1(_1803_),
    .A2(_1806_),
    .ZN(_0479_));
 AOI21_X1 _2426_ (.A(_1808_),
    .B1(_1811_),
    .B2(_1809_),
    .ZN(_0480_));
 OAI21_X1 _2427_ (.A(_0478_),
    .B1(_0479_),
    .B2(_0480_),
    .ZN(_0481_));
 NAND2_X1 _2428_ (.A1(_0477_),
    .A2(_0481_),
    .ZN(_0482_));
 INV_X1 _2429_ (.A(_1769_),
    .ZN(_0483_));
 INV_X1 _2430_ (.A(_1770_),
    .ZN(_0484_));
 OAI21_X1 _2431_ (.A(_0483_),
    .B1(_1764_),
    .B2(_0484_),
    .ZN(_0485_));
 AND2_X1 _2432_ (.A1(_1773_),
    .A2(_1776_),
    .ZN(_0486_));
 AOI221_X2 _2433_ (.A(_1772_),
    .B1(_0485_),
    .B2(_0486_),
    .C1(_1775_),
    .C2(_1773_),
    .ZN(_0487_));
 NAND2_X1 _2434_ (.A1(_1785_),
    .A2(_1788_),
    .ZN(_0488_));
 OR4_X1 _2435_ (.A1(_0466_),
    .A2(_0467_),
    .A3(_0470_),
    .A4(_0488_),
    .ZN(_0489_));
 OAI211_X2 _2436_ (.A(_0476_),
    .B(_0482_),
    .C1(_0487_),
    .C2(_0489_),
    .ZN(_0490_));
 AOI21_X1 _2437_ (.A(_0463_),
    .B1(_0465_),
    .B2(_0490_),
    .ZN(_0491_));
 AND2_X1 _2438_ (.A1(_0437_),
    .A2(net133),
    .ZN(_0492_));
 NAND2_X1 _2439_ (.A1(_1087_),
    .A2(_0492_),
    .ZN(_0493_));
 NOR4_X2 _2440_ (.A1(_0466_),
    .A2(_0467_),
    .A3(_0470_),
    .A4(_0488_),
    .ZN(_0494_));
 AND2_X1 _2441_ (.A1(_1770_),
    .A2(_1765_),
    .ZN(_0495_));
 NAND4_X2 _2442_ (.A1(_0486_),
    .A2(_0494_),
    .A3(_0495_),
    .A4(_0465_),
    .ZN(_0496_));
 NOR2_X1 _2443_ (.A1(_0493_),
    .A2(_0496_),
    .ZN(_0497_));
 OR3_X1 _2444_ (.A1(_0436_),
    .A2(_0491_),
    .A3(_0497_),
    .ZN(_0023_));
 CLKBUF_X3 _2445_ (.A(_0439_),
    .Z(_0498_));
 NAND2_X1 _2446_ (.A1(_0451_),
    .A2(_0462_),
    .ZN(_0499_));
 NAND3_X1 _2447_ (.A1(_0498_),
    .A2(_0499_),
    .A3(_0496_),
    .ZN(_0500_));
 NAND2_X1 _2448_ (.A1(_0439_),
    .A2(_0496_),
    .ZN(_0501_));
 NAND2_X1 _2449_ (.A1(_0490_),
    .A2(_0465_),
    .ZN(_0502_));
 NAND3_X4 _2450_ (.A1(_0435_),
    .A2(_0432_),
    .A3(_0434_),
    .ZN(_0503_));
 OAI221_X1 _2451_ (.A(_0500_),
    .B1(_0501_),
    .B2(_0502_),
    .C1(_1206_),
    .C2(_0503_),
    .ZN(_0022_));
 INV_X1 _2452_ (.A(\channel_state[3][2] ),
    .ZN(_0504_));
 NOR2_X1 _2453_ (.A1(_0504_),
    .A2(net137),
    .ZN(_0505_));
 AOI21_X1 _2454_ (.A(\channel_state[3][3] ),
    .B1(_0503_),
    .B2(_0505_),
    .ZN(_0506_));
 NOR2_X1 _2455_ (.A1(_0349_),
    .A2(_0506_),
    .ZN(_0021_));
 INV_X1 _2456_ (.A(_0437_),
    .ZN(_0507_));
 AND3_X2 _2457_ (.A1(_0435_),
    .A2(_0432_),
    .A3(_0434_),
    .ZN(_0508_));
 NOR3_X1 _2458_ (.A1(_0507_),
    .A2(net133),
    .A3(_0508_),
    .ZN(_0509_));
 OAI21_X1 _2459_ (.A(_0380_),
    .B1(\channel_state[3][5] ),
    .B2(_0509_),
    .ZN(_0510_));
 INV_X1 _2460_ (.A(_0510_),
    .ZN(_0020_));
 AND2_X1 _2461_ (.A1(_0432_),
    .A2(_0434_),
    .ZN(_0511_));
 INV_X1 _2462_ (.A(_0432_),
    .ZN(_0512_));
 AOI21_X1 _2463_ (.A(_0435_),
    .B1(\channel_state[3][4] ),
    .B2(_0512_),
    .ZN(_0513_));
 OAI21_X1 _2464_ (.A(_1090_),
    .B1(_0511_),
    .B2(_0513_),
    .ZN(_0019_));
 AND3_X1 _2465_ (.A1(net129),
    .A2(\channel_state[2][4] ),
    .A3(_0354_),
    .ZN(_0514_));
 AND2_X2 _2466_ (.A1(net132),
    .A2(_1179_),
    .ZN(_0515_));
 NAND2_X2 _2467_ (.A1(_1087_),
    .A2(_0515_),
    .ZN(_0516_));
 AOI211_X2 _2468_ (.A(_1167_),
    .B(_0516_),
    .C1(_1175_),
    .C2(_1203_),
    .ZN(_0517_));
 CLKBUF_X3 _2469_ (.A(_0516_),
    .Z(_0518_));
 NOR2_X2 _2470_ (.A1(_1177_),
    .A2(_0518_),
    .ZN(_0519_));
 OR3_X1 _2471_ (.A1(_0514_),
    .A2(_0517_),
    .A3(_0519_),
    .ZN(_0018_));
 AND3_X1 _2472_ (.A1(_0380_),
    .A2(\channel_state[1][2] ),
    .A3(net135),
    .ZN(_0001_));
 AND3_X1 _2473_ (.A1(_0380_),
    .A2(\channel_state[0][2] ),
    .A3(net134),
    .ZN(_0000_));
 AND3_X1 _2474_ (.A1(_0380_),
    .A2(\channel_state[3][2] ),
    .A3(net137),
    .ZN(_0003_));
 AND3_X1 _2475_ (.A1(_0380_),
    .A2(net136),
    .A3(\channel_state[2][2] ),
    .ZN(_0002_));
 INV_X1 _2476_ (.A(net89),
    .ZN(_1465_));
 NAND3_X2 _2477_ (.A1(_1100_),
    .A2(_1469_),
    .A3(_1108_),
    .ZN(_0520_));
 OR3_X1 _2478_ (.A1(_1114_),
    .A2(_1119_),
    .A3(_0520_),
    .ZN(_0521_));
 BUF_X4 _2479_ (.A(_0521_),
    .Z(_0522_));
 NOR3_X2 _2480_ (.A1(_1104_),
    .A2(_1106_),
    .A3(_0522_),
    .ZN(_0523_));
 XNOR2_X1 _2481_ (.A(_1131_),
    .B(_0523_),
    .ZN(_1495_));
 XNOR2_X1 _2482_ (.A(_1106_),
    .B(_0522_),
    .ZN(_1501_));
 INV_X1 _2483_ (.A(\transfer_count[2][30] ),
    .ZN(_0524_));
 NAND4_X2 _2484_ (.A1(_1118_),
    .A2(_1121_),
    .A3(_1122_),
    .A4(_1123_),
    .ZN(_0525_));
 OR2_X1 _2485_ (.A1(_0524_),
    .A2(_0525_),
    .ZN(_0526_));
 NOR4_X4 _2486_ (.A1(_1120_),
    .A2(_1129_),
    .A3(_1136_),
    .A4(_0526_),
    .ZN(_0527_));
 XNOR2_X2 _2487_ (.A(\transfer_count[2][31] ),
    .B(_0527_),
    .ZN(_1516_));
 INV_X1 _2488_ (.A(net54),
    .ZN(_1659_));
 INV_X1 _2489_ (.A(net1),
    .ZN(_1758_));
 INV_X2 _2490_ (.A(net124),
    .ZN(_1762_));
 XOR2_X2 _2491_ (.A(_1098_),
    .B(_1101_),
    .Z(_1474_));
 XNOR2_X2 _2492_ (.A(_1100_),
    .B(_1469_),
    .ZN(_1477_));
 NOR2_X1 _2493_ (.A1(_1101_),
    .A2(_1114_),
    .ZN(_0528_));
 XNOR2_X2 _2494_ (.A(_1108_),
    .B(_0528_),
    .ZN(_1480_));
 AND2_X1 _2495_ (.A1(_1100_),
    .A2(_1469_),
    .ZN(_0529_));
 NAND4_X2 _2496_ (.A1(_1098_),
    .A2(_1097_),
    .A3(_1099_),
    .A4(_0529_),
    .ZN(_0530_));
 XOR2_X2 _2497_ (.A(\transfer_count[2][6] ),
    .B(_0530_),
    .Z(_1483_));
 NAND2_X1 _2498_ (.A1(_1098_),
    .A2(_0529_),
    .ZN(_0531_));
 XOR2_X2 _2499_ (.A(_1099_),
    .B(_0531_),
    .Z(_1489_));
 NAND3_X1 _2500_ (.A1(_1131_),
    .A2(\transfer_count[2][13] ),
    .A3(_1105_),
    .ZN(_0532_));
 NOR2_X1 _2501_ (.A1(_1120_),
    .A2(_0532_),
    .ZN(_0533_));
 XNOR2_X1 _2502_ (.A(\transfer_count[2][15] ),
    .B(_0533_),
    .ZN(_1492_));
 NOR2_X1 _2503_ (.A1(_1109_),
    .A2(_1115_),
    .ZN(_0534_));
 XNOR2_X2 _2504_ (.A(\transfer_count[2][11] ),
    .B(_0534_),
    .ZN(_1504_));
 NOR4_X2 _2505_ (.A1(_1111_),
    .A2(_1113_),
    .A3(_1114_),
    .A4(_0520_),
    .ZN(_0535_));
 XNOR2_X2 _2506_ (.A(\transfer_count[2][10] ),
    .B(_0535_),
    .ZN(_1507_));
 NOR2_X2 _2507_ (.A1(_1114_),
    .A2(_0520_),
    .ZN(_0536_));
 XNOR2_X2 _2508_ (.A(_1112_),
    .B(_0536_),
    .ZN(_1513_));
 NOR4_X2 _2509_ (.A1(_1129_),
    .A2(_1136_),
    .A3(_0522_),
    .A4(_0525_),
    .ZN(_0537_));
 XNOR2_X1 _2510_ (.A(\transfer_count[2][30] ),
    .B(_0537_),
    .ZN(_1519_));
 NAND2_X1 _2511_ (.A1(_1122_),
    .A2(_1123_),
    .ZN(_0538_));
 NOR4_X2 _2512_ (.A1(_0538_),
    .A2(_1129_),
    .A3(_1136_),
    .A4(_0522_),
    .ZN(_0539_));
 XNOR2_X1 _2513_ (.A(_1121_),
    .B(_0539_),
    .ZN(_1525_));
 INV_X1 _2514_ (.A(_1122_),
    .ZN(_0540_));
 NAND4_X2 _2515_ (.A1(_1123_),
    .A2(\transfer_count[2][25] ),
    .A3(_1139_),
    .A4(_1140_),
    .ZN(_0541_));
 XNOR2_X2 _2516_ (.A(_0540_),
    .B(_0541_),
    .ZN(_1528_));
 OR2_X2 _2517_ (.A1(_1136_),
    .A2(_0521_),
    .ZN(_0542_));
 NOR2_X1 _2518_ (.A1(_1129_),
    .A2(_0542_),
    .ZN(_0543_));
 XNOR2_X1 _2519_ (.A(_1123_),
    .B(_0543_),
    .ZN(_1531_));
 INV_X1 _2520_ (.A(_1128_),
    .ZN(_0544_));
 NOR3_X2 _2521_ (.A1(_0544_),
    .A2(_1136_),
    .A3(_0522_),
    .ZN(_0545_));
 XNOR2_X1 _2522_ (.A(_1125_),
    .B(_0545_),
    .ZN(_1537_));
 AND3_X1 _2523_ (.A1(\transfer_count[2][22] ),
    .A2(_1126_),
    .A3(_1127_),
    .ZN(_0546_));
 NAND2_X1 _2524_ (.A1(_0546_),
    .A2(_1140_),
    .ZN(_0547_));
 XOR2_X2 _2525_ (.A(\transfer_count[2][23] ),
    .B(_0547_),
    .Z(_1540_));
 NAND2_X1 _2526_ (.A1(_1126_),
    .A2(_1127_),
    .ZN(_0548_));
 NOR2_X1 _2527_ (.A1(_0548_),
    .A2(_0542_),
    .ZN(_0549_));
 XNOR2_X2 _2528_ (.A(\transfer_count[2][22] ),
    .B(_0549_),
    .ZN(_1543_));
 XOR2_X2 _2529_ (.A(_1127_),
    .B(_0542_),
    .Z(_1549_));
 AND3_X1 _2530_ (.A1(_1133_),
    .A2(_1134_),
    .A3(_1144_),
    .ZN(_0550_));
 XNOR2_X1 _2531_ (.A(\transfer_count[2][19] ),
    .B(_0550_),
    .ZN(_1552_));
 INV_X1 _2532_ (.A(_1134_),
    .ZN(_0551_));
 NOR3_X2 _2533_ (.A1(_0551_),
    .A2(_1143_),
    .A3(_0522_),
    .ZN(_0552_));
 XNOR2_X1 _2534_ (.A(_1133_),
    .B(_0552_),
    .ZN(_1555_));
 INV_X1 _2535_ (.A(\transfer_count[2][15] ),
    .ZN(_0553_));
 NOR3_X2 _2536_ (.A1(_0553_),
    .A2(_0532_),
    .A3(_0522_),
    .ZN(_0554_));
 XNOR2_X1 _2537_ (.A(_1130_),
    .B(_0554_),
    .ZN(_1561_));
 INV_X1 _2538_ (.A(\transfer_count[1][31] ),
    .ZN(_0555_));
 INV_X1 _2539_ (.A(\transfer_count[1][30] ),
    .ZN(_0556_));
 AND3_X1 _2540_ (.A1(_1219_),
    .A2(_1223_),
    .A3(_1225_),
    .ZN(_0557_));
 NAND4_X2 _2541_ (.A1(_1216_),
    .A2(_1217_),
    .A3(_0557_),
    .A4(_1249_),
    .ZN(_0558_));
 NAND4_X2 _2542_ (.A1(\transfer_count[1][29] ),
    .A2(_1208_),
    .A3(_1209_),
    .A4(_1214_),
    .ZN(_0559_));
 OR3_X2 _2543_ (.A1(_0556_),
    .A2(_0558_),
    .A3(_0559_),
    .ZN(_0560_));
 XNOR2_X2 _2544_ (.A(_0555_),
    .B(_0560_),
    .ZN(_1564_));
 BUF_X2 _2545_ (.A(_1654_),
    .Z(_0561_));
 NAND3_X4 _2546_ (.A1(_1231_),
    .A2(_1232_),
    .A3(_0561_),
    .ZN(_0562_));
 OR4_X4 _2547_ (.A1(_1230_),
    .A2(_1237_),
    .A3(_1240_),
    .A4(_0562_),
    .ZN(_0563_));
 NOR4_X4 _2548_ (.A1(_1218_),
    .A2(_1226_),
    .A3(_0559_),
    .A4(_0563_),
    .ZN(_0564_));
 XNOR2_X1 _2549_ (.A(\transfer_count[1][30] ),
    .B(_0564_),
    .ZN(_1567_));
 NAND2_X1 _2550_ (.A1(_1209_),
    .A2(_1214_),
    .ZN(_0565_));
 NOR4_X2 _2551_ (.A1(_0565_),
    .A2(_1218_),
    .A3(_1226_),
    .A4(_0563_),
    .ZN(_0566_));
 XNOR2_X1 _2552_ (.A(_1208_),
    .B(_0566_),
    .ZN(_1573_));
 NAND3_X2 _2553_ (.A1(_1211_),
    .A2(_1212_),
    .A3(_1213_),
    .ZN(_0567_));
 NOR4_X4 _2554_ (.A1(_0567_),
    .A2(_1218_),
    .A3(_1226_),
    .A4(_0563_),
    .ZN(_0568_));
 XNOR2_X1 _2555_ (.A(_1210_),
    .B(_0568_),
    .ZN(_1579_));
 INV_X1 _2556_ (.A(_1213_),
    .ZN(_0569_));
 NOR4_X4 _2557_ (.A1(_0569_),
    .A2(_1218_),
    .A3(_1226_),
    .A4(_0563_),
    .ZN(_0570_));
 XNOR2_X1 _2558_ (.A(_1212_),
    .B(_0570_),
    .ZN(_1585_));
 NOR4_X4 _2559_ (.A1(_1230_),
    .A2(_1237_),
    .A3(_1240_),
    .A4(_0562_),
    .ZN(_0571_));
 AND3_X1 _2560_ (.A1(_1217_),
    .A2(_0557_),
    .A3(_0571_),
    .ZN(_0572_));
 XNOR2_X1 _2561_ (.A(_1216_),
    .B(_0572_),
    .ZN(_1591_));
 NAND3_X2 _2562_ (.A1(_1223_),
    .A2(_1225_),
    .A3(_0571_),
    .ZN(_0573_));
 XOR2_X2 _2563_ (.A(_1219_),
    .B(_0573_),
    .Z(_1597_));
 AND2_X1 _2564_ (.A1(_1223_),
    .A2(_0571_),
    .ZN(_0574_));
 XNOR2_X2 _2565_ (.A(_1224_),
    .B(_0574_),
    .ZN(_1603_));
 INV_X1 _2566_ (.A(\transfer_count[1][17] ),
    .ZN(_0575_));
 AND3_X1 _2567_ (.A1(_1220_),
    .A2(_1221_),
    .A3(_1222_),
    .ZN(_0576_));
 NAND2_X1 _2568_ (.A1(_0576_),
    .A2(_1249_),
    .ZN(_0577_));
 XNOR2_X2 _2569_ (.A(_0575_),
    .B(_0577_),
    .ZN(_1606_));
 AND3_X1 _2570_ (.A1(_1221_),
    .A2(_1222_),
    .A3(_0571_),
    .ZN(_0578_));
 XNOR2_X2 _2571_ (.A(_1220_),
    .B(_0578_),
    .ZN(_1609_));
 XNOR2_X2 _2572_ (.A(_1222_),
    .B(_0571_),
    .ZN(_1615_));
 INV_X1 _2573_ (.A(_1239_),
    .ZN(_0579_));
 NOR4_X2 _2574_ (.A1(_0579_),
    .A2(_1230_),
    .A3(_1237_),
    .A4(_0562_),
    .ZN(_0580_));
 XNOR2_X2 _2575_ (.A(_1238_),
    .B(_0580_),
    .ZN(_1621_));
 NOR2_X1 _2576_ (.A1(_1230_),
    .A2(_0562_),
    .ZN(_0581_));
 AND4_X1 _2577_ (.A1(\transfer_count[1][9] ),
    .A2(_1235_),
    .A3(_1236_),
    .A4(_0581_),
    .ZN(_0582_));
 XNOR2_X2 _2578_ (.A(\transfer_count[1][10] ),
    .B(_0582_),
    .ZN(_1627_));
 NAND2_X1 _2579_ (.A1(_1236_),
    .A2(_0581_),
    .ZN(_0583_));
 XOR2_X2 _2580_ (.A(_1235_),
    .B(_0583_),
    .Z(_1633_));
 AND3_X1 _2581_ (.A1(_1231_),
    .A2(_1232_),
    .A3(_0561_),
    .ZN(_0584_));
 AND3_X1 _2582_ (.A1(_1228_),
    .A2(_1229_),
    .A3(_0584_),
    .ZN(_0585_));
 XNOR2_X2 _2583_ (.A(_1227_),
    .B(_0585_),
    .ZN(_1639_));
 XNOR2_X2 _2584_ (.A(_1229_),
    .B(_0584_),
    .ZN(_1645_));
 XNOR2_X1 _2585_ (.A(_1232_),
    .B(_0561_),
    .ZN(_1651_));
 INV_X1 _2586_ (.A(\transfer_count[0][31] ),
    .ZN(_0586_));
 NAND3_X1 _2587_ (.A1(\transfer_count[0][30] ),
    .A2(_0226_),
    .A3(_0261_),
    .ZN(_0587_));
 XNOR2_X2 _2588_ (.A(_0586_),
    .B(_0587_),
    .ZN(_1663_));
 NAND4_X1 _2589_ (.A1(_0226_),
    .A2(_0251_),
    .A3(_0252_),
    .A4(_0256_),
    .ZN(_0588_));
 AND4_X2 _2590_ (.A1(_0227_),
    .A2(_0228_),
    .A3(_0229_),
    .A4(_0232_),
    .ZN(_0589_));
 NAND3_X4 _2591_ (.A1(_0238_),
    .A2(_0239_),
    .A3(_1753_),
    .ZN(_0590_));
 NOR4_X4 _2592_ (.A1(_0237_),
    .A2(_0244_),
    .A3(_0249_),
    .A4(_0590_),
    .ZN(_0591_));
 NAND4_X4 _2593_ (.A1(_0257_),
    .A2(_0258_),
    .A3(_0589_),
    .A4(_0591_),
    .ZN(_0592_));
 NOR2_X1 _2594_ (.A1(_0588_),
    .A2(_0592_),
    .ZN(_0593_));
 XNOR2_X2 _2595_ (.A(\transfer_count[0][30] ),
    .B(_0593_),
    .ZN(_1666_));
 NAND2_X1 _2596_ (.A1(_0252_),
    .A2(_0256_),
    .ZN(_0594_));
 NOR2_X1 _2597_ (.A1(_0594_),
    .A2(_0592_),
    .ZN(_0595_));
 XNOR2_X2 _2598_ (.A(_0251_),
    .B(_0595_),
    .ZN(_1672_));
 NAND3_X1 _2599_ (.A1(_0253_),
    .A2(_0254_),
    .A3(_0255_),
    .ZN(_0596_));
 NOR2_X1 _2600_ (.A1(_0596_),
    .A2(_0592_),
    .ZN(_0597_));
 XNOR2_X2 _2601_ (.A(\transfer_count[0][26] ),
    .B(_0597_),
    .ZN(_1678_));
 INV_X1 _2602_ (.A(_0255_),
    .ZN(_0598_));
 NOR2_X1 _2603_ (.A1(_0598_),
    .A2(_0592_),
    .ZN(_0599_));
 XNOR2_X2 _2604_ (.A(_0254_),
    .B(_0599_),
    .ZN(_1684_));
 NAND3_X2 _2605_ (.A1(_0246_),
    .A2(_0247_),
    .A3(_0248_),
    .ZN(_0600_));
 NOR3_X4 _2606_ (.A1(_0244_),
    .A2(_0600_),
    .A3(_0590_),
    .ZN(_0601_));
 INV_X1 _2607_ (.A(_0245_),
    .ZN(_0602_));
 NOR2_X1 _2608_ (.A1(_0602_),
    .A2(_0237_),
    .ZN(_0603_));
 NAND4_X2 _2609_ (.A1(_0258_),
    .A2(_0589_),
    .A3(_0601_),
    .A4(_0603_),
    .ZN(_0604_));
 XOR2_X2 _2610_ (.A(_0257_),
    .B(_0604_),
    .Z(_1690_));
 NAND3_X1 _2611_ (.A1(_0228_),
    .A2(_0229_),
    .A3(_0232_),
    .ZN(_0605_));
 OR4_X4 _2612_ (.A1(_0237_),
    .A2(_0244_),
    .A3(_0249_),
    .A4(_0590_),
    .ZN(_0606_));
 NOR2_X2 _2613_ (.A1(_0605_),
    .A2(_0606_),
    .ZN(_0607_));
 XNOR2_X2 _2614_ (.A(_0227_),
    .B(_0607_),
    .ZN(_1696_));
 INV_X1 _2615_ (.A(_0232_),
    .ZN(_0608_));
 NOR2_X1 _2616_ (.A1(_0608_),
    .A2(_0606_),
    .ZN(_0609_));
 XNOR2_X1 _2617_ (.A(_0229_),
    .B(_0609_),
    .ZN(_1702_));
 INV_X1 _2618_ (.A(\transfer_count[0][17] ),
    .ZN(_0610_));
 NAND4_X2 _2619_ (.A1(_0230_),
    .A2(\transfer_count[0][15] ),
    .A3(_0231_),
    .A4(_0270_),
    .ZN(_0611_));
 XNOR2_X2 _2620_ (.A(_0610_),
    .B(_0611_),
    .ZN(_1705_));
 INV_X1 _2621_ (.A(_0231_),
    .ZN(_0612_));
 NOR3_X2 _2622_ (.A1(_0272_),
    .A2(_0612_),
    .A3(_0606_),
    .ZN(_0613_));
 XNOR2_X1 _2623_ (.A(_0230_),
    .B(_0613_),
    .ZN(_1708_));
 XNOR2_X1 _2624_ (.A(_0612_),
    .B(_0606_),
    .ZN(_1714_));
 NAND3_X2 _2625_ (.A1(_0236_),
    .A2(_0245_),
    .A3(_0601_),
    .ZN(_0614_));
 XOR2_X2 _2626_ (.A(_0235_),
    .B(_0614_),
    .Z(_1720_));
 XNOR2_X1 _2627_ (.A(_0245_),
    .B(_0601_),
    .ZN(_1726_));
 INV_X1 _2628_ (.A(_0248_),
    .ZN(_0615_));
 NOR3_X2 _2629_ (.A1(_0615_),
    .A2(_0244_),
    .A3(_0590_),
    .ZN(_0616_));
 XNOR2_X2 _2630_ (.A(_0247_),
    .B(_0616_),
    .ZN(_1732_));
 INV_X1 _2631_ (.A(_0242_),
    .ZN(_0617_));
 NOR3_X2 _2632_ (.A1(_0617_),
    .A2(_0278_),
    .A3(_0590_),
    .ZN(_0618_));
 XNOR2_X1 _2633_ (.A(_0241_),
    .B(_0618_),
    .ZN(_1738_));
 XNOR2_X1 _2634_ (.A(_0278_),
    .B(_0590_),
    .ZN(_1744_));
 XNOR2_X2 _2635_ (.A(_0239_),
    .B(_1753_),
    .ZN(_1750_));
 XNOR2_X1 _2636_ (.A(_0391_),
    .B(_0395_),
    .ZN(_1771_));
 BUF_X1 _2637_ (.A(_1766_),
    .Z(_0619_));
 XNOR2_X1 _2638_ (.A(_0393_),
    .B(_0619_),
    .ZN(_1774_));
 NAND2_X1 _2639_ (.A1(_0395_),
    .A2(_0404_),
    .ZN(_0620_));
 XOR2_X2 _2640_ (.A(_0402_),
    .B(_0620_),
    .Z(_1777_));
 AND2_X2 _2641_ (.A1(_0393_),
    .A2(_0619_),
    .ZN(_0621_));
 NAND4_X2 _2642_ (.A1(_0391_),
    .A2(_0390_),
    .A3(_0392_),
    .A4(_0621_),
    .ZN(_0622_));
 XOR2_X2 _2643_ (.A(\transfer_count[3][6] ),
    .B(_0622_),
    .Z(_1780_));
 NAND2_X1 _2644_ (.A1(_0391_),
    .A2(_0621_),
    .ZN(_0623_));
 XOR2_X2 _2645_ (.A(_0392_),
    .B(_0623_),
    .Z(_1786_));
 AND4_X1 _2646_ (.A1(\transfer_count[3][14] ),
    .A2(_0397_),
    .A3(_0401_),
    .A4(_0406_),
    .ZN(_0624_));
 XNOR2_X1 _2647_ (.A(\transfer_count[3][15] ),
    .B(_0624_),
    .ZN(_1789_));
 INV_X1 _2648_ (.A(\transfer_count[3][14] ),
    .ZN(_0625_));
 AND4_X2 _2649_ (.A1(_0402_),
    .A2(_0403_),
    .A3(_0404_),
    .A4(_0621_),
    .ZN(_0626_));
 NAND3_X1 _2650_ (.A1(_0397_),
    .A2(_0401_),
    .A3(_0626_),
    .ZN(_0627_));
 XNOR2_X1 _2651_ (.A(_0625_),
    .B(_0627_),
    .ZN(_1792_));
 NAND4_X2 _2652_ (.A1(_0398_),
    .A2(_0399_),
    .A3(_0400_),
    .A4(_0626_),
    .ZN(_0628_));
 XOR2_X2 _2653_ (.A(\transfer_count[3][12] ),
    .B(_0628_),
    .Z(_1798_));
 NAND3_X2 _2654_ (.A1(_0399_),
    .A2(_0400_),
    .A3(_0406_),
    .ZN(_0629_));
 XOR2_X2 _2655_ (.A(_0398_),
    .B(_0629_),
    .Z(_1801_));
 NAND2_X1 _2656_ (.A1(_0400_),
    .A2(_0626_),
    .ZN(_0630_));
 XOR2_X2 _2657_ (.A(_0399_),
    .B(_0630_),
    .Z(_1804_));
 INV_X1 _2658_ (.A(_0403_),
    .ZN(_0631_));
 NAND3_X2 _2659_ (.A1(_0402_),
    .A2(_0404_),
    .A3(_0621_),
    .ZN(_0632_));
 XNOR2_X1 _2660_ (.A(_0631_),
    .B(_0632_),
    .ZN(_1810_));
 INV_X1 _2661_ (.A(\transfer_count[3][31] ),
    .ZN(_0633_));
 NOR3_X4 _2662_ (.A1(_0430_),
    .A2(_0420_),
    .A3(_0423_),
    .ZN(_0634_));
 AND3_X1 _2663_ (.A1(\transfer_count[3][29] ),
    .A2(\transfer_count[3][28] ),
    .A3(_0411_),
    .ZN(_0635_));
 NAND3_X1 _2664_ (.A1(\transfer_count[3][30] ),
    .A2(_0634_),
    .A3(_0635_),
    .ZN(_0636_));
 XNOR2_X1 _2665_ (.A(_0633_),
    .B(_0636_),
    .ZN(_1813_));
 INV_X1 _2666_ (.A(\transfer_count[3][30] ),
    .ZN(_0637_));
 NAND4_X4 _2667_ (.A1(_0402_),
    .A2(_0403_),
    .A3(_0404_),
    .A4(_0621_),
    .ZN(_0638_));
 NOR3_X4 _2668_ (.A1(_0420_),
    .A2(_0423_),
    .A3(_0638_),
    .ZN(_0639_));
 NAND2_X1 _2669_ (.A1(_0635_),
    .A2(_0639_),
    .ZN(_0640_));
 XNOR2_X1 _2670_ (.A(_0637_),
    .B(_0640_),
    .ZN(_1816_));
 INV_X1 _2671_ (.A(\transfer_count[3][28] ),
    .ZN(_0641_));
 NAND2_X1 _2672_ (.A1(_0411_),
    .A2(_0639_),
    .ZN(_0642_));
 XNOR2_X1 _2673_ (.A(_0641_),
    .B(_0642_),
    .ZN(_1822_));
 NAND3_X1 _2674_ (.A1(_0409_),
    .A2(_0410_),
    .A3(_0424_),
    .ZN(_0643_));
 XOR2_X2 _2675_ (.A(\transfer_count[3][27] ),
    .B(_0643_),
    .Z(_1825_));
 INV_X1 _2676_ (.A(\transfer_count[3][26] ),
    .ZN(_0644_));
 NAND3_X1 _2677_ (.A1(\transfer_count[3][25] ),
    .A2(_0409_),
    .A3(_0639_),
    .ZN(_0645_));
 XNOR2_X1 _2678_ (.A(_0644_),
    .B(_0645_),
    .ZN(_1828_));
 INV_X1 _2679_ (.A(\transfer_count[3][24] ),
    .ZN(_0646_));
 NAND2_X1 _2680_ (.A1(_0408_),
    .A2(_0639_),
    .ZN(_0647_));
 XNOR2_X1 _2681_ (.A(_0646_),
    .B(_0647_),
    .ZN(_1834_));
 XNOR2_X2 _2682_ (.A(_0408_),
    .B(_0634_),
    .ZN(_1837_));
 NAND3_X2 _2683_ (.A1(_0417_),
    .A2(\transfer_count[3][18] ),
    .A3(_0418_),
    .ZN(_0648_));
 NAND2_X1 _2684_ (.A1(_0415_),
    .A2(_0416_),
    .ZN(_0649_));
 NOR4_X4 _2685_ (.A1(_0648_),
    .A2(_0649_),
    .A3(_0423_),
    .A4(_0638_),
    .ZN(_0650_));
 XNOR2_X1 _2686_ (.A(_0414_),
    .B(_0650_),
    .ZN(_1840_));
 OR3_X2 _2687_ (.A1(_0648_),
    .A2(_0423_),
    .A3(_0638_),
    .ZN(_0651_));
 XOR2_X2 _2688_ (.A(_0416_),
    .B(_0651_),
    .Z(_1846_));
 AND4_X1 _2689_ (.A1(\transfer_count[3][18] ),
    .A2(_0418_),
    .A3(_0406_),
    .A4(_0428_),
    .ZN(_0652_));
 XNOR2_X1 _2690_ (.A(_0417_),
    .B(_0652_),
    .ZN(_1849_));
 INV_X1 _2691_ (.A(\transfer_count[3][18] ),
    .ZN(_0653_));
 NOR2_X1 _2692_ (.A1(_0423_),
    .A2(_0638_),
    .ZN(_0654_));
 NAND2_X1 _2693_ (.A1(_0418_),
    .A2(_0654_),
    .ZN(_0655_));
 XNOR2_X1 _2694_ (.A(_0653_),
    .B(_0655_),
    .ZN(_1852_));
 AND3_X1 _2695_ (.A1(_0401_),
    .A2(_0422_),
    .A3(_0626_),
    .ZN(_0656_));
 XNOR2_X2 _2696_ (.A(_0421_),
    .B(_0656_),
    .ZN(_1858_));
 INV_X1 _2697_ (.A(_1470_),
    .ZN(_1471_));
 INV_X1 _2698_ (.A(_1655_),
    .ZN(_1656_));
 INV_X1 _2699_ (.A(_1754_),
    .ZN(_1755_));
 INV_X1 _2700_ (.A(_1767_),
    .ZN(_1768_));
 NOR3_X1 _2701_ (.A1(_0281_),
    .A2(\channel_state[0][2] ),
    .A3(\channel_state[0][3] ),
    .ZN(_0657_));
 NOR2_X1 _2702_ (.A1(_0337_),
    .A2(\channel_state[0][5] ),
    .ZN(_0658_));
 NAND2_X1 _2703_ (.A1(_0657_),
    .A2(_0658_),
    .ZN(_0659_));
 NAND3_X1 _2704_ (.A1(_0283_),
    .A2(net138),
    .A3(_0659_),
    .ZN(_0660_));
 NOR2_X1 _2705_ (.A1(\active_channel_count[0] ),
    .A2(_0660_),
    .ZN(_0661_));
 NAND2_X1 _2706_ (.A1(_1094_),
    .A2(net140),
    .ZN(_0662_));
 NOR2_X2 _2707_ (.A1(_1179_),
    .A2(\channel_state[2][5] ),
    .ZN(_0663_));
 NOR3_X2 _2708_ (.A1(_1091_),
    .A2(\channel_state[2][2] ),
    .A3(\channel_state[2][3] ),
    .ZN(_0664_));
 AOI21_X4 _2709_ (.A(_0662_),
    .B1(_0663_),
    .B2(_0664_),
    .ZN(_0665_));
 NAND2_X1 _2710_ (.A1(_0434_),
    .A2(net141),
    .ZN(_0666_));
 NOR2_X2 _2711_ (.A1(\channel_state[3][5] ),
    .A2(_0437_),
    .ZN(_0667_));
 NOR3_X1 _2712_ (.A1(_0435_),
    .A2(\channel_state[3][2] ),
    .A3(\channel_state[3][3] ),
    .ZN(_0668_));
 AOI21_X2 _2713_ (.A(_0666_),
    .B1(_0667_),
    .B2(_0668_),
    .ZN(_0669_));
 NAND2_X1 _2714_ (.A1(_1262_),
    .A2(net139),
    .ZN(_0670_));
 NOR2_X2 _2715_ (.A1(\channel_state[1][1] ),
    .A2(\channel_state[1][5] ),
    .ZN(_0671_));
 NOR3_X2 _2716_ (.A1(_1261_),
    .A2(\channel_state[1][3] ),
    .A3(\channel_state[1][2] ),
    .ZN(_0672_));
 AOI21_X4 _2717_ (.A(_0670_),
    .B1(_0671_),
    .B2(_0672_),
    .ZN(_0673_));
 NOR3_X4 _2718_ (.A1(_0665_),
    .A2(_0669_),
    .A3(_0673_),
    .ZN(_0674_));
 MUX2_X1 _2719_ (.A(_1861_),
    .B(_0661_),
    .S(_0674_),
    .Z(_0675_));
 AND2_X1 _2720_ (.A1(_1090_),
    .A2(_0675_),
    .ZN(_0024_));
 NAND2_X1 _2721_ (.A1(_0674_),
    .A2(_0660_),
    .ZN(_0676_));
 AND3_X1 _2722_ (.A1(_0380_),
    .A2(_1864_),
    .A3(_0676_),
    .ZN(_0025_));
 BUF_X8 _2723_ (.A(_1088_),
    .Z(_0677_));
 NAND2_X1 _2724_ (.A1(_0677_),
    .A2(_0676_),
    .ZN(_0678_));
 XNOR2_X1 _2725_ (.A(_1865_),
    .B(\active_channel_count[2] ),
    .ZN(_0679_));
 NOR2_X1 _2726_ (.A1(_0678_),
    .A2(_0679_),
    .ZN(_0026_));
 NAND3_X1 _2727_ (.A1(\active_channel_count[0] ),
    .A2(\active_channel_count[2] ),
    .A3(\active_channel_count[1] ),
    .ZN(_0680_));
 XOR2_X1 _2728_ (.A(\active_channel_count[3] ),
    .B(_0680_),
    .Z(_0681_));
 NOR2_X1 _2729_ (.A1(_0678_),
    .A2(_0681_),
    .ZN(_0027_));
 OAI21_X1 _2730_ (.A(_0677_),
    .B1(net138),
    .B2(_0374_),
    .ZN(_0682_));
 INV_X1 _2731_ (.A(net138),
    .ZN(_0683_));
 AOI21_X1 _2732_ (.A(_1205_),
    .B1(_0683_),
    .B2(_0284_),
    .ZN(_0684_));
 NAND3_X1 _2733_ (.A1(_0344_),
    .A2(_0347_),
    .A3(_0684_),
    .ZN(_0685_));
 OAI22_X1 _2734_ (.A1(_0368_),
    .A2(_0682_),
    .B1(_0685_),
    .B2(_0336_),
    .ZN(_0028_));
 CLKBUF_X3 _2735_ (.A(_1266_),
    .Z(_0686_));
 OAI21_X1 _2736_ (.A(_0677_),
    .B1(net139),
    .B2(_0358_),
    .ZN(_0687_));
 INV_X1 _2737_ (.A(net139),
    .ZN(_0688_));
 AOI21_X1 _2738_ (.A(_1205_),
    .B1(_0688_),
    .B2(_0220_),
    .ZN(_0689_));
 NAND3_X1 _2739_ (.A1(_0214_),
    .A2(_0217_),
    .A3(_0689_),
    .ZN(_0690_));
 OAI22_X1 _2740_ (.A1(_0686_),
    .A2(_0687_),
    .B1(_0690_),
    .B2(_0225_),
    .ZN(_0029_));
 CLKBUF_X3 _2741_ (.A(_1180_),
    .Z(_0691_));
 OAI221_X1 _2742_ (.A(_0677_),
    .B1(net140),
    .B2(_0353_),
    .C1(_0691_),
    .C2(_1177_),
    .ZN(_0692_));
 CLKBUF_X3 _2743_ (.A(_1180_),
    .Z(_0693_));
 NOR2_X1 _2744_ (.A1(_0693_),
    .A2(_1167_),
    .ZN(_0694_));
 AOI21_X1 _2745_ (.A(_0692_),
    .B1(_0694_),
    .B2(_1204_),
    .ZN(_0030_));
 CLKBUF_X3 _2746_ (.A(_0438_),
    .Z(_0695_));
 OAI221_X1 _2747_ (.A(_0677_),
    .B1(_0695_),
    .B2(_0496_),
    .C1(_0508_),
    .C2(net141),
    .ZN(_0696_));
 CLKBUF_X3 _2748_ (.A(_0438_),
    .Z(_0697_));
 NOR2_X1 _2749_ (.A1(_0697_),
    .A2(_0499_),
    .ZN(_0698_));
 AOI21_X1 _2750_ (.A(_0696_),
    .B1(_0698_),
    .B2(_0502_),
    .ZN(_0031_));
 NAND3_X1 _2751_ (.A1(_0373_),
    .A2(\channel_state[0][4] ),
    .A3(_0385_),
    .ZN(_0699_));
 NAND4_X1 _2752_ (.A1(_1087_),
    .A2(net142),
    .A3(_0284_),
    .A4(_0699_),
    .ZN(_0700_));
 AND2_X1 _2753_ (.A1(_0347_),
    .A2(_0700_),
    .ZN(_0701_));
 OAI211_X2 _2754_ (.A(_0344_),
    .B(_0701_),
    .C1(_0310_),
    .C2(_0335_),
    .ZN(_0702_));
 NAND2_X1 _2755_ (.A1(_0370_),
    .A2(_0700_),
    .ZN(_0703_));
 AND2_X1 _2756_ (.A1(_0702_),
    .A2(_0703_),
    .ZN(_0032_));
 NAND3_X1 _2757_ (.A1(_0388_),
    .A2(\channel_state[1][4] ),
    .A3(_0381_),
    .ZN(_0704_));
 NAND3_X1 _2758_ (.A1(net143),
    .A2(_0359_),
    .A3(_0704_),
    .ZN(_0705_));
 AND3_X1 _2759_ (.A1(_0214_),
    .A2(_0217_),
    .A3(_0705_),
    .ZN(_0706_));
 AOI22_X1 _2760_ (.A1(_1268_),
    .A2(_0705_),
    .B1(_0706_),
    .B2(_0210_),
    .ZN(_0033_));
 NAND3_X1 _2761_ (.A1(_1093_),
    .A2(\channel_state[2][4] ),
    .A3(_0377_),
    .ZN(_0707_));
 AND3_X1 _2762_ (.A1(net144),
    .A2(_0354_),
    .A3(_0707_),
    .ZN(_0708_));
 OR3_X1 _2763_ (.A1(_0517_),
    .A2(_0519_),
    .A3(_0708_),
    .ZN(_0034_));
 NAND3_X1 _2764_ (.A1(_0507_),
    .A2(\channel_state[3][4] ),
    .A3(_0512_),
    .ZN(_0709_));
 AND4_X1 _2765_ (.A1(_1088_),
    .A2(net145),
    .A3(_0503_),
    .A4(_0709_),
    .ZN(_0710_));
 OR3_X1 _2766_ (.A1(_0491_),
    .A2(_0497_),
    .A3(_0710_),
    .ZN(_0035_));
 AND2_X1 _2767_ (.A1(_1090_),
    .A2(\active_channel_count[0] ),
    .ZN(_0036_));
 AND2_X1 _2768_ (.A1(_1090_),
    .A2(\active_channel_count[1] ),
    .ZN(_0037_));
 AND2_X1 _2769_ (.A1(_1090_),
    .A2(\active_channel_count[2] ),
    .ZN(_0038_));
 AND2_X1 _2770_ (.A1(_1090_),
    .A2(\active_channel_count[3] ),
    .ZN(_0039_));
 NOR2_X1 _2771_ (.A1(\active_channel_count[2] ),
    .A2(\active_channel_count[3] ),
    .ZN(_0711_));
 AOI21_X1 _2772_ (.A(_0219_),
    .B1(_1863_),
    .B2(_0711_),
    .ZN(_0040_));
 BUF_X4 _2773_ (.A(_1205_),
    .Z(_0712_));
 INV_X1 _2774_ (.A(\channel_state[0][4] ),
    .ZN(_0713_));
 AND2_X1 _2775_ (.A1(_0713_),
    .A2(_0657_),
    .ZN(_0714_));
 NAND2_X1 _2776_ (.A1(net151),
    .A2(_0714_),
    .ZN(_0715_));
 AOI21_X1 _2777_ (.A(_0712_),
    .B1(_0658_),
    .B2(_0715_),
    .ZN(_0041_));
 INV_X1 _2778_ (.A(\channel_state[1][4] ),
    .ZN(_0716_));
 AND2_X1 _2779_ (.A1(_0716_),
    .A2(_0672_),
    .ZN(_0717_));
 NAND2_X1 _2780_ (.A1(net152),
    .A2(_0717_),
    .ZN(_0718_));
 AOI21_X1 _2781_ (.A(_0712_),
    .B1(_0671_),
    .B2(_0718_),
    .ZN(_0042_));
 NOR4_X2 _2782_ (.A1(\channel_state[2][4] ),
    .A2(_1091_),
    .A3(\channel_state[2][2] ),
    .A4(\channel_state[2][3] ),
    .ZN(_0719_));
 NAND2_X1 _2783_ (.A1(net153),
    .A2(_0719_),
    .ZN(_0720_));
 AOI21_X1 _2784_ (.A(_0712_),
    .B1(_0663_),
    .B2(_0720_),
    .ZN(_0043_));
 INV_X1 _2785_ (.A(\channel_state[3][4] ),
    .ZN(_0721_));
 AND2_X1 _2786_ (.A1(_0721_),
    .A2(_0668_),
    .ZN(_0722_));
 NAND2_X1 _2787_ (.A1(net154),
    .A2(_0722_),
    .ZN(_0723_));
 AOI21_X1 _2788_ (.A(_0712_),
    .B1(_0667_),
    .B2(_0723_),
    .ZN(_0044_));
 AND2_X1 _2789_ (.A1(_1090_),
    .A2(\channel_state[0][3] ),
    .ZN(_0045_));
 BUF_X4 _2790_ (.A(_1089_),
    .Z(_0724_));
 AND2_X1 _2791_ (.A1(_0724_),
    .A2(\channel_state[3][3] ),
    .ZN(_0048_));
 NAND3_X1 _2792_ (.A1(net159),
    .A2(_0658_),
    .A3(_0714_),
    .ZN(_0725_));
 NOR2_X1 _2793_ (.A1(\channel_state[0][3] ),
    .A2(_0351_),
    .ZN(_0726_));
 AOI21_X1 _2794_ (.A(_0712_),
    .B1(_0725_),
    .B2(_0726_),
    .ZN(_0049_));
 NAND3_X1 _2795_ (.A1(net160),
    .A2(_0671_),
    .A3(_0717_),
    .ZN(_0727_));
 NOR2_X1 _2796_ (.A1(\channel_state[1][3] ),
    .A2(_0361_),
    .ZN(_0728_));
 AOI21_X1 _2797_ (.A(_0712_),
    .B1(_0727_),
    .B2(_0728_),
    .ZN(_0050_));
 NAND3_X1 _2798_ (.A1(net161),
    .A2(_0663_),
    .A3(_0719_),
    .ZN(_0729_));
 NOR2_X1 _2799_ (.A1(\channel_state[2][3] ),
    .A2(_0356_),
    .ZN(_0730_));
 AOI21_X1 _2800_ (.A(_0712_),
    .B1(_0729_),
    .B2(_0730_),
    .ZN(_0051_));
 NAND3_X1 _2801_ (.A1(net162),
    .A2(_0667_),
    .A3(_0722_),
    .ZN(_0731_));
 NOR2_X1 _2802_ (.A1(\channel_state[3][3] ),
    .A2(_0505_),
    .ZN(_0732_));
 AOI21_X1 _2803_ (.A(_0712_),
    .B1(_0731_),
    .B2(_0732_),
    .ZN(_0052_));
 NAND2_X1 _2804_ (.A1(_1759_),
    .A2(_0368_),
    .ZN(_0733_));
 CLKBUF_X3 _2805_ (.A(_0338_),
    .Z(_0734_));
 NAND3_X1 _2806_ (.A1(\transfer_count[0][0] ),
    .A2(_0285_),
    .A3(_0734_),
    .ZN(_0735_));
 AOI21_X1 _2807_ (.A(_0712_),
    .B1(_0733_),
    .B2(_0735_),
    .ZN(_0053_));
 NAND2_X2 _2808_ (.A1(_0284_),
    .A2(_0338_),
    .ZN(_0736_));
 CLKBUF_X3 _2809_ (.A(_0338_),
    .Z(_0737_));
 OAI21_X1 _2810_ (.A(_0736_),
    .B1(_0601_),
    .B2(_0737_),
    .ZN(_0738_));
 NAND2_X1 _2811_ (.A1(_0245_),
    .A2(_0738_),
    .ZN(_0739_));
 NAND3_X1 _2812_ (.A1(_0602_),
    .A2(_0368_),
    .A3(_0601_),
    .ZN(_0740_));
 AOI21_X1 _2813_ (.A(_0712_),
    .B1(_0739_),
    .B2(_0740_),
    .ZN(_0054_));
 NAND3_X1 _2814_ (.A1(_0236_),
    .A2(_0285_),
    .A3(_0737_),
    .ZN(_0741_));
 OAI21_X1 _2815_ (.A(_0741_),
    .B1(_0734_),
    .B2(_1723_),
    .ZN(_0742_));
 AND2_X1 _2816_ (.A1(_0724_),
    .A2(_0742_),
    .ZN(_0055_));
 BUF_X4 _2817_ (.A(_1205_),
    .Z(_0743_));
 NOR2_X4 _2818_ (.A1(_0374_),
    .A2(_0368_),
    .ZN(_0744_));
 AND2_X1 _2819_ (.A1(_0368_),
    .A2(_0614_),
    .ZN(_0745_));
 OAI21_X1 _2820_ (.A(_0235_),
    .B1(_0744_),
    .B2(_0745_),
    .ZN(_0746_));
 OR3_X1 _2821_ (.A1(_0235_),
    .A2(_0338_),
    .A3(_0614_),
    .ZN(_0747_));
 AOI21_X1 _2822_ (.A(_0743_),
    .B1(_0746_),
    .B2(_0747_),
    .ZN(_0056_));
 OAI21_X1 _2823_ (.A(_0736_),
    .B1(_0737_),
    .B2(_0275_),
    .ZN(_0748_));
 NOR2_X1 _2824_ (.A1(_0234_),
    .A2(_0737_),
    .ZN(_0749_));
 AOI22_X1 _2825_ (.A1(_0234_),
    .A2(_0748_),
    .B1(_0749_),
    .B2(_0275_),
    .ZN(_0750_));
 NOR2_X1 _2826_ (.A1(_0349_),
    .A2(_0750_),
    .ZN(_0057_));
 AOI21_X1 _2827_ (.A(_0744_),
    .B1(_0606_),
    .B2(_0368_),
    .ZN(_0751_));
 NOR2_X1 _2828_ (.A1(_0612_),
    .A2(_0751_),
    .ZN(_0752_));
 NOR3_X1 _2829_ (.A1(_0231_),
    .A2(_0734_),
    .A3(_0606_),
    .ZN(_0753_));
 OAI21_X1 _2830_ (.A(_0380_),
    .B1(_0752_),
    .B2(_0753_),
    .ZN(_0754_));
 INV_X1 _2831_ (.A(_0754_),
    .ZN(_0058_));
 NAND2_X2 _2832_ (.A1(_1087_),
    .A2(_0744_),
    .ZN(_0755_));
 CLKBUF_X3 _2833_ (.A(_0755_),
    .Z(_0756_));
 OAI22_X1 _2834_ (.A1(_1711_),
    .A2(_0370_),
    .B1(_0756_),
    .B2(_0272_),
    .ZN(_0059_));
 OAI21_X1 _2835_ (.A(_0756_),
    .B1(_0613_),
    .B2(_0370_),
    .ZN(_0757_));
 NAND2_X1 _2836_ (.A1(_0230_),
    .A2(_0757_),
    .ZN(_0758_));
 NAND2_X1 _2837_ (.A1(_0340_),
    .A2(_0613_),
    .ZN(_0759_));
 OAI21_X1 _2838_ (.A(_0758_),
    .B1(_0759_),
    .B2(_0230_),
    .ZN(_0060_));
 OAI22_X1 _2839_ (.A1(_0370_),
    .A2(_1705_),
    .B1(_0756_),
    .B2(_0610_),
    .ZN(_0061_));
 OAI21_X1 _2840_ (.A(_0756_),
    .B1(_0609_),
    .B2(_0370_),
    .ZN(_0760_));
 NAND2_X1 _2841_ (.A1(_0229_),
    .A2(_0760_),
    .ZN(_0761_));
 NAND2_X1 _2842_ (.A1(_0340_),
    .A2(_0609_),
    .ZN(_0762_));
 OAI21_X1 _2843_ (.A(_0761_),
    .B1(_0762_),
    .B2(_0229_),
    .ZN(_0062_));
 OAI21_X1 _2844_ (.A(_0756_),
    .B1(_0370_),
    .B2(_0271_),
    .ZN(_0763_));
 CLKBUF_X3 _2845_ (.A(_0369_),
    .Z(_0764_));
 NOR2_X1 _2846_ (.A1(_0228_),
    .A2(_0764_),
    .ZN(_0765_));
 AOI22_X1 _2847_ (.A1(_0228_),
    .A2(_0763_),
    .B1(_0765_),
    .B2(_0271_),
    .ZN(_0766_));
 INV_X1 _2848_ (.A(_0766_),
    .ZN(_0063_));
 NAND2_X1 _2849_ (.A1(_1754_),
    .A2(_0368_),
    .ZN(_0767_));
 NAND3_X1 _2850_ (.A1(\transfer_count[0][1] ),
    .A2(_0285_),
    .A3(_0734_),
    .ZN(_0768_));
 AOI21_X1 _2851_ (.A(_0743_),
    .B1(_0767_),
    .B2(_0768_),
    .ZN(_0064_));
 OAI21_X1 _2852_ (.A(_0756_),
    .B1(_0607_),
    .B2(_0370_),
    .ZN(_0769_));
 NAND2_X1 _2853_ (.A1(_0227_),
    .A2(_0769_),
    .ZN(_0770_));
 NAND2_X1 _2854_ (.A1(_0340_),
    .A2(_0607_),
    .ZN(_0771_));
 OAI21_X1 _2855_ (.A(_0770_),
    .B1(_0771_),
    .B2(_0227_),
    .ZN(_0065_));
 NAND4_X1 _2856_ (.A1(_0269_),
    .A2(_0589_),
    .A3(_0270_),
    .A4(_0340_),
    .ZN(_0772_));
 AOI22_X1 _2857_ (.A1(_0266_),
    .A2(_0340_),
    .B1(_0744_),
    .B2(_0677_),
    .ZN(_0773_));
 OAI21_X1 _2858_ (.A(_0772_),
    .B1(_0773_),
    .B2(_0269_),
    .ZN(_0066_));
 OR4_X1 _2859_ (.A1(_1205_),
    .A2(_0257_),
    .A3(_0338_),
    .A4(_0604_),
    .ZN(_0774_));
 NAND2_X1 _2860_ (.A1(_0677_),
    .A2(_0257_),
    .ZN(_0775_));
 AOI21_X1 _2861_ (.A(_0744_),
    .B1(_0604_),
    .B2(_0368_),
    .ZN(_0776_));
 OAI21_X1 _2862_ (.A(_0774_),
    .B1(_0775_),
    .B2(_0776_),
    .ZN(_0067_));
 AOI21_X1 _2863_ (.A(_0255_),
    .B1(_0268_),
    .B2(_0340_),
    .ZN(_0777_));
 AOI21_X1 _2864_ (.A(_0598_),
    .B1(_0744_),
    .B2(_0677_),
    .ZN(_0778_));
 OAI21_X1 _2865_ (.A(_0340_),
    .B1(_0266_),
    .B2(_0265_),
    .ZN(_0779_));
 AOI21_X1 _2866_ (.A(_0777_),
    .B1(_0778_),
    .B2(_0779_),
    .ZN(_0068_));
 NOR3_X1 _2867_ (.A1(_0598_),
    .A2(_0764_),
    .A3(_0592_),
    .ZN(_0780_));
 OAI21_X1 _2868_ (.A(_0756_),
    .B1(_0599_),
    .B2(_0764_),
    .ZN(_0781_));
 MUX2_X1 _2869_ (.A(_0780_),
    .B(_0781_),
    .S(_0254_),
    .Z(_0069_));
 AOI21_X1 _2870_ (.A(_0253_),
    .B1(_0267_),
    .B2(_0340_),
    .ZN(_0782_));
 AND2_X1 _2871_ (.A1(_0253_),
    .A2(_0756_),
    .ZN(_0783_));
 OR2_X1 _2872_ (.A1(_0267_),
    .A2(_0764_),
    .ZN(_0784_));
 AOI21_X1 _2873_ (.A(_0782_),
    .B1(_0783_),
    .B2(_0784_),
    .ZN(_0070_));
 NOR3_X1 _2874_ (.A1(_0596_),
    .A2(_0764_),
    .A3(_0592_),
    .ZN(_0785_));
 OAI21_X1 _2875_ (.A(_0755_),
    .B1(_0597_),
    .B2(_0764_),
    .ZN(_0786_));
 MUX2_X1 _2876_ (.A(_0785_),
    .B(_0786_),
    .S(\transfer_count[0][26] ),
    .Z(_0071_));
 OAI21_X1 _2877_ (.A(_0756_),
    .B1(_0370_),
    .B2(_0263_),
    .ZN(_0787_));
 NAND2_X1 _2878_ (.A1(_0252_),
    .A2(_0787_),
    .ZN(_0788_));
 NAND2_X1 _2879_ (.A1(_0263_),
    .A2(_0340_),
    .ZN(_0789_));
 OAI21_X1 _2880_ (.A(_0788_),
    .B1(_0789_),
    .B2(_0252_),
    .ZN(_0072_));
 NOR3_X1 _2881_ (.A1(_0594_),
    .A2(_0369_),
    .A3(_0592_),
    .ZN(_0790_));
 OAI21_X1 _2882_ (.A(_0755_),
    .B1(_0595_),
    .B2(_0764_),
    .ZN(_0791_));
 MUX2_X1 _2883_ (.A(_0790_),
    .B(_0791_),
    .S(_0251_),
    .Z(_0073_));
 AND2_X1 _2884_ (.A1(_0261_),
    .A2(_0339_),
    .ZN(_0792_));
 OAI21_X1 _2885_ (.A(_0755_),
    .B1(_0764_),
    .B2(_0261_),
    .ZN(_0793_));
 MUX2_X1 _2886_ (.A(_0792_),
    .B(_0793_),
    .S(_0226_),
    .Z(_0074_));
 OR2_X1 _2887_ (.A1(_0734_),
    .A2(_1750_),
    .ZN(_0794_));
 NAND3_X1 _2888_ (.A1(_0239_),
    .A2(_0285_),
    .A3(_0734_),
    .ZN(_0795_));
 AOI21_X1 _2889_ (.A(_0743_),
    .B1(_0794_),
    .B2(_0795_),
    .ZN(_0075_));
 NOR3_X1 _2890_ (.A1(_0764_),
    .A2(_0588_),
    .A3(_0592_),
    .ZN(_0796_));
 OAI21_X1 _2891_ (.A(_0755_),
    .B1(_0593_),
    .B2(_0764_),
    .ZN(_0797_));
 MUX2_X1 _2892_ (.A(_0796_),
    .B(_0797_),
    .S(\transfer_count[0][30] ),
    .Z(_0076_));
 OAI22_X1 _2893_ (.A1(_0370_),
    .A2(_1663_),
    .B1(_0756_),
    .B2(_0586_),
    .ZN(_0077_));
 NAND3_X1 _2894_ (.A1(_0238_),
    .A2(_0285_),
    .A3(_0737_),
    .ZN(_0798_));
 OAI21_X1 _2895_ (.A(_0798_),
    .B1(_0734_),
    .B2(_1747_),
    .ZN(_0799_));
 AND2_X1 _2896_ (.A1(_0724_),
    .A2(_0799_),
    .ZN(_0078_));
 AND2_X1 _2897_ (.A1(_0368_),
    .A2(_0590_),
    .ZN(_0800_));
 OAI21_X1 _2898_ (.A(_0243_),
    .B1(_0744_),
    .B2(_0800_),
    .ZN(_0801_));
 OR3_X1 _2899_ (.A1(_0243_),
    .A2(_0338_),
    .A3(_0590_),
    .ZN(_0802_));
 AOI21_X1 _2900_ (.A(_0743_),
    .B1(_0801_),
    .B2(_0802_),
    .ZN(_0079_));
 NAND3_X1 _2901_ (.A1(_0242_),
    .A2(_0285_),
    .A3(_0737_),
    .ZN(_0803_));
 OAI21_X1 _2902_ (.A(_0803_),
    .B1(_0734_),
    .B2(_1741_),
    .ZN(_0804_));
 AND2_X1 _2903_ (.A1(_0724_),
    .A2(_0804_),
    .ZN(_0080_));
 OAI21_X1 _2904_ (.A(_0736_),
    .B1(_0618_),
    .B2(_0737_),
    .ZN(_0805_));
 NOR2_X1 _2905_ (.A1(_0241_),
    .A2(_0338_),
    .ZN(_0806_));
 AOI22_X1 _2906_ (.A1(_0241_),
    .A2(_0805_),
    .B1(_0806_),
    .B2(_0618_),
    .ZN(_0807_));
 NOR2_X1 _2907_ (.A1(_0349_),
    .A2(_0807_),
    .ZN(_0081_));
 NAND3_X1 _2908_ (.A1(_0248_),
    .A2(_0285_),
    .A3(_0737_),
    .ZN(_0808_));
 OAI21_X1 _2909_ (.A(_0808_),
    .B1(_0734_),
    .B2(_1735_),
    .ZN(_0809_));
 AND2_X1 _2910_ (.A1(_0724_),
    .A2(_0809_),
    .ZN(_0082_));
 NAND3_X1 _2911_ (.A1(_0247_),
    .A2(_0285_),
    .A3(_0737_),
    .ZN(_0810_));
 OAI21_X1 _2912_ (.A(_0810_),
    .B1(_1732_),
    .B2(_0734_),
    .ZN(_0811_));
 AND2_X1 _2913_ (.A1(_0724_),
    .A2(_0811_),
    .ZN(_0083_));
 OAI21_X1 _2914_ (.A(_0736_),
    .B1(_0737_),
    .B2(_0277_),
    .ZN(_0812_));
 NOR2_X1 _2915_ (.A1(_0246_),
    .A2(_0338_),
    .ZN(_0813_));
 AOI22_X1 _2916_ (.A1(_0246_),
    .A2(_0812_),
    .B1(_0813_),
    .B2(_0277_),
    .ZN(_0814_));
 NOR2_X1 _2917_ (.A1(_0349_),
    .A2(_0814_),
    .ZN(_0084_));
 NAND2_X1 _2918_ (.A1(_1660_),
    .A2(_0686_),
    .ZN(_0815_));
 BUF_X4 _2919_ (.A(_0221_),
    .Z(_0816_));
 CLKBUF_X3 _2920_ (.A(_0816_),
    .Z(_0817_));
 NAND3_X1 _2921_ (.A1(\transfer_count[1][0] ),
    .A2(_0817_),
    .A3(_0220_),
    .ZN(_0818_));
 AOI21_X1 _2922_ (.A(_0743_),
    .B1(_0815_),
    .B2(_0818_),
    .ZN(_0085_));
 CLKBUF_X3 _2923_ (.A(_0221_),
    .Z(_0819_));
 NAND3_X1 _2924_ (.A1(\transfer_count[1][10] ),
    .A2(_0819_),
    .A3(_0220_),
    .ZN(_0820_));
 OAI21_X1 _2925_ (.A(_0820_),
    .B1(_1627_),
    .B2(_0817_),
    .ZN(_0821_));
 AND2_X1 _2926_ (.A1(_0724_),
    .A2(_0821_),
    .ZN(_0086_));
 NAND2_X4 _2927_ (.A1(_0221_),
    .A2(_0220_),
    .ZN(_0822_));
 OAI21_X1 _2928_ (.A(_0822_),
    .B1(_0819_),
    .B2(_1253_),
    .ZN(_0823_));
 NOR2_X1 _2929_ (.A1(_1239_),
    .A2(_0819_),
    .ZN(_0824_));
 AOI22_X1 _2930_ (.A1(_1239_),
    .A2(_0823_),
    .B1(_0824_),
    .B2(_1253_),
    .ZN(_0825_));
 NOR2_X1 _2931_ (.A1(_0349_),
    .A2(_0825_),
    .ZN(_0087_));
 INV_X1 _2932_ (.A(_1238_),
    .ZN(_0826_));
 OAI22_X1 _2933_ (.A1(_0817_),
    .A2(_1621_),
    .B1(_0822_),
    .B2(_0826_),
    .ZN(_0827_));
 AND2_X1 _2934_ (.A1(_0724_),
    .A2(_0827_),
    .ZN(_0088_));
 NOR2_X1 _2935_ (.A1(_1254_),
    .A2(_0817_),
    .ZN(_0828_));
 NAND2_X1 _2936_ (.A1(\transfer_count[1][13] ),
    .A2(_0359_),
    .ZN(_0829_));
 OAI22_X1 _2937_ (.A1(_1618_),
    .A2(_1268_),
    .B1(_0828_),
    .B2(_0829_),
    .ZN(_0089_));
 NOR3_X1 _2938_ (.A1(_1222_),
    .A2(_0816_),
    .A3(_0563_),
    .ZN(_0830_));
 OAI21_X1 _2939_ (.A(_0822_),
    .B1(_0571_),
    .B2(_0817_),
    .ZN(_0831_));
 AOI21_X1 _2940_ (.A(_0830_),
    .B1(_0831_),
    .B2(_1222_),
    .ZN(_0832_));
 NOR2_X1 _2941_ (.A1(_0349_),
    .A2(_0832_),
    .ZN(_0090_));
 NOR2_X1 _2942_ (.A1(_1252_),
    .A2(_0819_),
    .ZN(_0833_));
 NAND2_X1 _2943_ (.A1(_1221_),
    .A2(_0822_),
    .ZN(_0834_));
 AOI21_X1 _2944_ (.A(_0819_),
    .B1(_1249_),
    .B2(_1222_),
    .ZN(_0835_));
 OAI221_X1 _2945_ (.A(_0380_),
    .B1(_1221_),
    .B2(_0833_),
    .C1(_0834_),
    .C2(_0835_),
    .ZN(_0836_));
 INV_X1 _2946_ (.A(_0836_),
    .ZN(_0091_));
 OAI21_X1 _2947_ (.A(_0822_),
    .B1(_0578_),
    .B2(_0819_),
    .ZN(_0837_));
 NOR2_X1 _2948_ (.A1(_1220_),
    .A2(_0816_),
    .ZN(_0838_));
 AOI22_X1 _2949_ (.A1(_1220_),
    .A2(_0837_),
    .B1(_0838_),
    .B2(_0578_),
    .ZN(_0839_));
 NOR2_X1 _2950_ (.A1(_0349_),
    .A2(_0839_),
    .ZN(_0092_));
 NOR2_X2 _2951_ (.A1(_1266_),
    .A2(_0358_),
    .ZN(_0840_));
 AOI21_X1 _2952_ (.A(_0816_),
    .B1(_1249_),
    .B2(_0576_),
    .ZN(_0841_));
 OAI21_X1 _2953_ (.A(\transfer_count[1][17] ),
    .B1(_0840_),
    .B2(_0841_),
    .ZN(_0842_));
 NAND4_X1 _2954_ (.A1(_0575_),
    .A2(_0576_),
    .A3(_1249_),
    .A4(_1266_),
    .ZN(_0843_));
 AOI21_X1 _2955_ (.A(_0743_),
    .B1(_0842_),
    .B2(_0843_),
    .ZN(_0093_));
 OAI21_X1 _2956_ (.A(_0822_),
    .B1(_0574_),
    .B2(_0817_),
    .ZN(_0844_));
 NAND2_X1 _2957_ (.A1(_1224_),
    .A2(_0844_),
    .ZN(_0845_));
 INV_X1 _2958_ (.A(_1224_),
    .ZN(_0846_));
 NAND3_X1 _2959_ (.A1(_0846_),
    .A2(_0686_),
    .A3(_0574_),
    .ZN(_0847_));
 AOI21_X1 _2960_ (.A(_0743_),
    .B1(_0845_),
    .B2(_0847_),
    .ZN(_0094_));
 INV_X1 _2961_ (.A(\transfer_count[1][19] ),
    .ZN(_0848_));
 NAND3_X1 _2962_ (.A1(_0848_),
    .A2(_1251_),
    .A3(_0223_),
    .ZN(_0849_));
 NAND2_X1 _2963_ (.A1(\transfer_count[1][19] ),
    .A2(_0222_),
    .ZN(_0850_));
 NAND2_X4 _2964_ (.A1(_0816_),
    .A2(_0359_),
    .ZN(_0851_));
 OAI221_X1 _2965_ (.A(_0849_),
    .B1(_0850_),
    .B2(_1251_),
    .C1(_0848_),
    .C2(_0851_),
    .ZN(_0095_));
 NAND2_X1 _2966_ (.A1(_1655_),
    .A2(_0686_),
    .ZN(_0852_));
 NAND3_X1 _2967_ (.A1(\transfer_count[1][1] ),
    .A2(_0817_),
    .A3(_0220_),
    .ZN(_0853_));
 AOI21_X1 _2968_ (.A(_0743_),
    .B1(_0852_),
    .B2(_0853_),
    .ZN(_0096_));
 OR4_X1 _2969_ (.A1(_1205_),
    .A2(_1219_),
    .A3(_0816_),
    .A4(_0573_),
    .ZN(_0854_));
 NAND2_X1 _2970_ (.A1(_0677_),
    .A2(_1219_),
    .ZN(_0855_));
 AOI21_X1 _2971_ (.A(_0840_),
    .B1(_0573_),
    .B2(_0686_),
    .ZN(_0856_));
 OAI21_X1 _2972_ (.A(_0854_),
    .B1(_0855_),
    .B2(_0856_),
    .ZN(_0097_));
 NOR2_X1 _2973_ (.A1(_1242_),
    .A2(_0816_),
    .ZN(_0857_));
 NOR2_X1 _2974_ (.A1(_1217_),
    .A2(_0857_),
    .ZN(_0858_));
 NAND2_X1 _2975_ (.A1(_1217_),
    .A2(_0822_),
    .ZN(_0859_));
 AOI21_X1 _2976_ (.A(_0859_),
    .B1(_1266_),
    .B2(_1242_),
    .ZN(_0860_));
 NOR3_X1 _2977_ (.A1(_0219_),
    .A2(_0858_),
    .A3(_0860_),
    .ZN(_0098_));
 OAI21_X1 _2978_ (.A(_0851_),
    .B1(_0572_),
    .B2(_1268_),
    .ZN(_0861_));
 NAND2_X1 _2979_ (.A1(_1216_),
    .A2(_0861_),
    .ZN(_0862_));
 NAND2_X1 _2980_ (.A1(_0223_),
    .A2(_0572_),
    .ZN(_0863_));
 OAI21_X1 _2981_ (.A(_0862_),
    .B1(_0863_),
    .B2(_1216_),
    .ZN(_0099_));
 OAI21_X1 _2982_ (.A(_0822_),
    .B1(_0817_),
    .B2(_1244_),
    .ZN(_0864_));
 NAND2_X1 _2983_ (.A1(_1213_),
    .A2(_0864_),
    .ZN(_0865_));
 NAND3_X1 _2984_ (.A1(_0569_),
    .A2(_1244_),
    .A3(_0686_),
    .ZN(_0866_));
 AOI21_X1 _2985_ (.A(_0743_),
    .B1(_0865_),
    .B2(_0866_),
    .ZN(_0100_));
 OAI21_X1 _2986_ (.A(_0851_),
    .B1(_0570_),
    .B2(_1268_),
    .ZN(_0867_));
 NAND2_X1 _2987_ (.A1(_1212_),
    .A2(_0867_),
    .ZN(_0868_));
 NAND2_X1 _2988_ (.A1(_0223_),
    .A2(_0570_),
    .ZN(_0869_));
 OAI21_X1 _2989_ (.A(_0868_),
    .B1(_0869_),
    .B2(_1212_),
    .ZN(_0101_));
 NOR3_X1 _2990_ (.A1(_1246_),
    .A2(_0558_),
    .A3(_1267_),
    .ZN(_0870_));
 OAI21_X1 _2991_ (.A(_0851_),
    .B1(_1268_),
    .B2(_1247_),
    .ZN(_0871_));
 MUX2_X1 _2992_ (.A(_0870_),
    .B(_0871_),
    .S(_1211_),
    .Z(_0102_));
 OAI21_X1 _2993_ (.A(_0851_),
    .B1(_0568_),
    .B2(_1268_),
    .ZN(_0872_));
 NAND2_X1 _2994_ (.A1(_1210_),
    .A2(_0872_),
    .ZN(_0873_));
 NAND2_X1 _2995_ (.A1(_0223_),
    .A2(_0568_),
    .ZN(_0874_));
 OAI21_X1 _2996_ (.A(_0873_),
    .B1(_0874_),
    .B2(_1210_),
    .ZN(_0103_));
 NOR3_X2 _2997_ (.A1(_1205_),
    .A2(_1266_),
    .A3(_0358_),
    .ZN(_0875_));
 AOI21_X1 _2998_ (.A(_1267_),
    .B1(_1244_),
    .B2(_1214_),
    .ZN(_0876_));
 OAI21_X1 _2999_ (.A(_1209_),
    .B1(_0875_),
    .B2(_0876_),
    .ZN(_0877_));
 NAND3_X1 _3000_ (.A1(_1214_),
    .A2(_1244_),
    .A3(_0223_),
    .ZN(_0878_));
 OAI21_X1 _3001_ (.A(_0877_),
    .B1(_0878_),
    .B2(_1209_),
    .ZN(_0104_));
 OAI21_X1 _3002_ (.A(_0851_),
    .B1(_0566_),
    .B2(_1268_),
    .ZN(_0879_));
 NAND2_X1 _3003_ (.A1(_1208_),
    .A2(_0879_),
    .ZN(_0880_));
 NAND2_X1 _3004_ (.A1(_0223_),
    .A2(_0566_),
    .ZN(_0881_));
 OAI21_X1 _3005_ (.A(_0880_),
    .B1(_0881_),
    .B2(_1208_),
    .ZN(_0105_));
 NOR3_X1 _3006_ (.A1(_1215_),
    .A2(_0558_),
    .A3(_1267_),
    .ZN(_0882_));
 OAI21_X1 _3007_ (.A(_0851_),
    .B1(_1268_),
    .B2(_1243_),
    .ZN(_0883_));
 MUX2_X1 _3008_ (.A(_0882_),
    .B(_0883_),
    .S(\transfer_count[1][29] ),
    .Z(_0106_));
 NOR2_X1 _3009_ (.A1(_0561_),
    .A2(_0819_),
    .ZN(_0884_));
 OAI21_X1 _3010_ (.A(_1232_),
    .B1(_0840_),
    .B2(_0884_),
    .ZN(_0885_));
 INV_X1 _3011_ (.A(_1232_),
    .ZN(_0886_));
 NAND3_X1 _3012_ (.A1(_0886_),
    .A2(_0561_),
    .A3(_0686_),
    .ZN(_0887_));
 AOI21_X1 _3013_ (.A(_0743_),
    .B1(_0885_),
    .B2(_0887_),
    .ZN(_0107_));
 OAI21_X1 _3014_ (.A(_0851_),
    .B1(_0564_),
    .B2(_1268_),
    .ZN(_0888_));
 NAND2_X1 _3015_ (.A1(\transfer_count[1][30] ),
    .A2(_0888_),
    .ZN(_0889_));
 NAND3_X1 _3016_ (.A1(_0556_),
    .A2(_0223_),
    .A3(_0564_),
    .ZN(_0890_));
 NAND2_X1 _3017_ (.A1(_0889_),
    .A2(_0890_),
    .ZN(_0108_));
 OR3_X1 _3018_ (.A1(\transfer_count[1][31] ),
    .A2(_1267_),
    .A3(_0560_),
    .ZN(_0891_));
 AOI21_X1 _3019_ (.A(_0875_),
    .B1(_0560_),
    .B2(_0223_),
    .ZN(_0892_));
 OAI21_X1 _3020_ (.A(_0891_),
    .B1(_0892_),
    .B2(_0555_),
    .ZN(_0109_));
 BUF_X4 _3021_ (.A(_1205_),
    .Z(_0893_));
 AND2_X1 _3022_ (.A1(_1259_),
    .A2(_1266_),
    .ZN(_0894_));
 OAI21_X1 _3023_ (.A(_1231_),
    .B1(_0840_),
    .B2(_0894_),
    .ZN(_0895_));
 OR3_X1 _3024_ (.A1(_1231_),
    .A2(_1259_),
    .A3(_0816_),
    .ZN(_0896_));
 AOI21_X1 _3025_ (.A(_0893_),
    .B1(_0895_),
    .B2(_0896_),
    .ZN(_0110_));
 NOR2_X1 _3026_ (.A1(_0817_),
    .A2(_0584_),
    .ZN(_0897_));
 OAI21_X1 _3027_ (.A(_1229_),
    .B1(_0840_),
    .B2(_0897_),
    .ZN(_0898_));
 NAND3_X1 _3028_ (.A1(_1257_),
    .A2(_0686_),
    .A3(_0584_),
    .ZN(_0899_));
 AOI21_X1 _3029_ (.A(_0893_),
    .B1(_0898_),
    .B2(_0899_),
    .ZN(_0111_));
 AOI21_X1 _3030_ (.A(_0223_),
    .B1(_0359_),
    .B2(_1228_),
    .ZN(_0900_));
 AOI21_X1 _3031_ (.A(_0900_),
    .B1(_0686_),
    .B2(_1642_),
    .ZN(_0112_));
 OAI21_X1 _3032_ (.A(_0822_),
    .B1(_0585_),
    .B2(_0819_),
    .ZN(_0901_));
 NOR2_X1 _3033_ (.A1(_1227_),
    .A2(_0816_),
    .ZN(_0902_));
 AOI22_X1 _3034_ (.A1(_1227_),
    .A2(_0901_),
    .B1(_0902_),
    .B2(_0585_),
    .ZN(_0903_));
 NOR2_X1 _3035_ (.A1(_0349_),
    .A2(_0903_),
    .ZN(_0113_));
 OAI21_X1 _3036_ (.A(_0822_),
    .B1(_0819_),
    .B2(_1255_),
    .ZN(_0904_));
 NOR2_X1 _3037_ (.A1(_1236_),
    .A2(_0816_),
    .ZN(_0905_));
 AOI22_X1 _3038_ (.A1(_1236_),
    .A2(_0904_),
    .B1(_0905_),
    .B2(_1255_),
    .ZN(_0906_));
 NOR2_X1 _3039_ (.A1(_0349_),
    .A2(_0906_),
    .ZN(_0114_));
 AOI21_X1 _3040_ (.A(_0222_),
    .B1(_0359_),
    .B2(_1235_),
    .ZN(_0907_));
 AOI21_X1 _3041_ (.A(_0907_),
    .B1(_1633_),
    .B2(_0686_),
    .ZN(_0115_));
 NAND3_X1 _3042_ (.A1(\transfer_count[1][9] ),
    .A2(_0819_),
    .A3(_0220_),
    .ZN(_0908_));
 OAI21_X1 _3043_ (.A(_0908_),
    .B1(_0817_),
    .B2(_1630_),
    .ZN(_0909_));
 AND2_X1 _3044_ (.A1(_0724_),
    .A2(_0909_),
    .ZN(_0116_));
 NAND2_X1 _3045_ (.A1(_1466_),
    .A2(_0515_),
    .ZN(_0910_));
 NAND3_X1 _3046_ (.A1(\transfer_count[2][0] ),
    .A2(_1207_),
    .A3(_0693_),
    .ZN(_0911_));
 AOI21_X1 _3047_ (.A(_0893_),
    .B1(_0910_),
    .B2(_0911_),
    .ZN(_0117_));
 CLKBUF_X3 _3048_ (.A(_0516_),
    .Z(_0912_));
 NAND2_X1 _3049_ (.A1(_1180_),
    .A2(_0354_),
    .ZN(_0913_));
 CLKBUF_X3 _3050_ (.A(_0913_),
    .Z(_0914_));
 OAI22_X1 _3051_ (.A1(_0912_),
    .A2(_1507_),
    .B1(_0914_),
    .B2(_1110_),
    .ZN(_0118_));
 NAND2_X2 _3052_ (.A1(_1207_),
    .A2(_1180_),
    .ZN(_0915_));
 OAI22_X1 _3053_ (.A1(_0693_),
    .A2(_1504_),
    .B1(_0915_),
    .B2(_1107_),
    .ZN(_0916_));
 AND2_X1 _3054_ (.A1(_0724_),
    .A2(_0916_),
    .ZN(_0119_));
 NOR3_X1 _3055_ (.A1(_1105_),
    .A2(_1180_),
    .A3(_0522_),
    .ZN(_0917_));
 INV_X1 _3056_ (.A(_0522_),
    .ZN(_0918_));
 OAI21_X1 _3057_ (.A(_0915_),
    .B1(_0918_),
    .B2(_0691_),
    .ZN(_0919_));
 AOI21_X1 _3058_ (.A(_0917_),
    .B1(_0919_),
    .B2(_1105_),
    .ZN(_0920_));
 NOR2_X1 _3059_ (.A1(_0219_),
    .A2(_0920_),
    .ZN(_0120_));
 OR4_X1 _3060_ (.A1(\transfer_count[2][13] ),
    .A2(_1106_),
    .A3(_1120_),
    .A4(_0516_),
    .ZN(_0921_));
 NOR3_X4 _3061_ (.A1(_1178_),
    .A2(_0353_),
    .A3(_0515_),
    .ZN(_0922_));
 CLKBUF_X3 _3062_ (.A(_1181_),
    .Z(_0923_));
 AOI21_X1 _3063_ (.A(_0922_),
    .B1(_0923_),
    .B2(_1116_),
    .ZN(_0924_));
 OAI21_X1 _3064_ (.A(_0921_),
    .B1(_0924_),
    .B2(_1104_),
    .ZN(_0121_));
 OAI21_X1 _3065_ (.A(_0914_),
    .B1(_0523_),
    .B2(_0912_),
    .ZN(_0925_));
 NAND2_X1 _3066_ (.A1(_1131_),
    .A2(_0925_),
    .ZN(_0926_));
 NAND2_X1 _3067_ (.A1(_0923_),
    .A2(_0523_),
    .ZN(_0927_));
 OAI21_X1 _3068_ (.A(_0926_),
    .B1(_0927_),
    .B2(_1131_),
    .ZN(_0122_));
 OAI21_X1 _3069_ (.A(_0914_),
    .B1(_0533_),
    .B2(_0912_),
    .ZN(_0928_));
 NAND2_X1 _3070_ (.A1(\transfer_count[2][15] ),
    .A2(_0928_),
    .ZN(_0929_));
 NAND3_X1 _3071_ (.A1(_0553_),
    .A2(_0923_),
    .A3(_0533_),
    .ZN(_0930_));
 NAND2_X1 _3072_ (.A1(_0929_),
    .A2(_0930_),
    .ZN(_0123_));
 OAI21_X1 _3073_ (.A(_0914_),
    .B1(_0554_),
    .B2(_0912_),
    .ZN(_0931_));
 NAND2_X1 _3074_ (.A1(_1130_),
    .A2(_0931_),
    .ZN(_0932_));
 NAND2_X1 _3075_ (.A1(_0923_),
    .A2(_0554_),
    .ZN(_0933_));
 OAI21_X1 _3076_ (.A(_0932_),
    .B1(_0933_),
    .B2(_1130_),
    .ZN(_0124_));
 OAI21_X1 _3077_ (.A(_0914_),
    .B1(_0912_),
    .B2(_1144_),
    .ZN(_0934_));
 NAND2_X1 _3078_ (.A1(_1134_),
    .A2(_0934_),
    .ZN(_0935_));
 NAND3_X1 _3079_ (.A1(_0551_),
    .A2(_1144_),
    .A3(_0923_),
    .ZN(_0936_));
 NAND2_X1 _3080_ (.A1(_0935_),
    .A2(_0936_),
    .ZN(_0125_));
 OAI21_X1 _3081_ (.A(_0914_),
    .B1(_0552_),
    .B2(_0912_),
    .ZN(_0937_));
 NAND2_X1 _3082_ (.A1(_1133_),
    .A2(_0937_),
    .ZN(_0938_));
 NAND2_X1 _3083_ (.A1(_0923_),
    .A2(_0552_),
    .ZN(_0939_));
 OAI21_X1 _3084_ (.A(_0938_),
    .B1(_0939_),
    .B2(_1133_),
    .ZN(_0126_));
 AND2_X1 _3085_ (.A1(_1181_),
    .A2(_0550_),
    .ZN(_0940_));
 OAI21_X1 _3086_ (.A(_0913_),
    .B1(_0550_),
    .B2(_0518_),
    .ZN(_0941_));
 MUX2_X1 _3087_ (.A(_0940_),
    .B(_0941_),
    .S(\transfer_count[2][19] ),
    .Z(_0127_));
 NAND2_X1 _3088_ (.A1(_1470_),
    .A2(_0515_),
    .ZN(_0942_));
 NAND3_X1 _3089_ (.A1(\transfer_count[2][1] ),
    .A2(_1207_),
    .A3(_0693_),
    .ZN(_0943_));
 AOI21_X1 _3090_ (.A(_0893_),
    .B1(_0942_),
    .B2(_0943_),
    .ZN(_0128_));
 OR3_X1 _3091_ (.A1(_1127_),
    .A2(_0691_),
    .A3(_0542_),
    .ZN(_0944_));
 OAI21_X1 _3092_ (.A(_0515_),
    .B1(_0522_),
    .B2(_1136_),
    .ZN(_0945_));
 NAND2_X1 _3093_ (.A1(_0915_),
    .A2(_0945_),
    .ZN(_0946_));
 NAND2_X1 _3094_ (.A1(_1127_),
    .A2(_0946_),
    .ZN(_0947_));
 AOI21_X1 _3095_ (.A(_0893_),
    .B1(_0944_),
    .B2(_0947_),
    .ZN(_0129_));
 AOI21_X1 _3096_ (.A(_0518_),
    .B1(_1140_),
    .B2(_1127_),
    .ZN(_0948_));
 OAI21_X1 _3097_ (.A(_1126_),
    .B1(_0922_),
    .B2(_0948_),
    .ZN(_0949_));
 NAND3_X1 _3098_ (.A1(_1127_),
    .A2(_1140_),
    .A3(_1181_),
    .ZN(_0950_));
 OAI21_X1 _3099_ (.A(_0949_),
    .B1(_0950_),
    .B2(_1126_),
    .ZN(_0130_));
 NOR3_X1 _3100_ (.A1(_0548_),
    .A2(_0691_),
    .A3(_0542_),
    .ZN(_0951_));
 NAND2_X1 _3101_ (.A1(\transfer_count[2][22] ),
    .A2(_0354_),
    .ZN(_0952_));
 OAI22_X1 _3102_ (.A1(_0912_),
    .A2(_1543_),
    .B1(_0951_),
    .B2(_0952_),
    .ZN(_0131_));
 AOI21_X1 _3103_ (.A(_0518_),
    .B1(_1140_),
    .B2(_0546_),
    .ZN(_0953_));
 OAI21_X1 _3104_ (.A(\transfer_count[2][23] ),
    .B1(_0922_),
    .B2(_0953_),
    .ZN(_0954_));
 NAND3_X1 _3105_ (.A1(_0546_),
    .A2(_1140_),
    .A3(_1181_),
    .ZN(_0955_));
 OAI21_X1 _3106_ (.A(_0954_),
    .B1(_0955_),
    .B2(\transfer_count[2][23] ),
    .ZN(_0132_));
 OAI21_X1 _3107_ (.A(_0914_),
    .B1(_0545_),
    .B2(_0518_),
    .ZN(_0956_));
 NAND2_X1 _3108_ (.A1(_1125_),
    .A2(_0956_),
    .ZN(_0957_));
 NAND2_X1 _3109_ (.A1(_0923_),
    .A2(_0545_),
    .ZN(_0958_));
 OAI21_X1 _3110_ (.A(_0957_),
    .B1(_0958_),
    .B2(_1125_),
    .ZN(_0133_));
 NAND4_X1 _3111_ (.A1(_1138_),
    .A2(_1139_),
    .A3(_1140_),
    .A4(_1181_),
    .ZN(_0959_));
 AOI21_X1 _3112_ (.A(_0922_),
    .B1(_1181_),
    .B2(_1141_),
    .ZN(_0960_));
 OAI21_X1 _3113_ (.A(_0959_),
    .B1(_0960_),
    .B2(_1138_),
    .ZN(_0134_));
 NOR3_X1 _3114_ (.A1(_1129_),
    .A2(_0518_),
    .A3(_0542_),
    .ZN(_0961_));
 OAI21_X1 _3115_ (.A(_0913_),
    .B1(_0543_),
    .B2(_0518_),
    .ZN(_0962_));
 MUX2_X1 _3116_ (.A(_0961_),
    .B(_0962_),
    .S(_1123_),
    .Z(_0135_));
 OR3_X1 _3117_ (.A1(_1122_),
    .A2(_0518_),
    .A3(_0541_),
    .ZN(_0963_));
 AOI21_X1 _3118_ (.A(_0922_),
    .B1(_0541_),
    .B2(_1181_),
    .ZN(_0964_));
 OAI21_X1 _3119_ (.A(_0963_),
    .B1(_0964_),
    .B2(_0540_),
    .ZN(_0136_));
 OAI21_X1 _3120_ (.A(_0914_),
    .B1(_0539_),
    .B2(_0518_),
    .ZN(_0965_));
 NAND2_X1 _3121_ (.A1(_1121_),
    .A2(_0965_),
    .ZN(_0966_));
 NAND2_X1 _3122_ (.A1(_0923_),
    .A2(_0539_),
    .ZN(_0967_));
 OAI21_X1 _3123_ (.A(_0966_),
    .B1(_0967_),
    .B2(_1121_),
    .ZN(_0137_));
 OAI21_X1 _3124_ (.A(_0914_),
    .B1(_0912_),
    .B2(_1137_),
    .ZN(_0968_));
 NAND2_X1 _3125_ (.A1(_1118_),
    .A2(_0968_),
    .ZN(_0969_));
 NAND2_X1 _3126_ (.A1(_1137_),
    .A2(_0923_),
    .ZN(_0970_));
 OAI21_X1 _3127_ (.A(_0969_),
    .B1(_0970_),
    .B2(_1118_),
    .ZN(_0138_));
 OR2_X1 _3128_ (.A1(_0691_),
    .A2(_1477_),
    .ZN(_0971_));
 NAND3_X1 _3129_ (.A1(_1100_),
    .A2(_1207_),
    .A3(_0693_),
    .ZN(_0972_));
 AOI21_X1 _3130_ (.A(_0893_),
    .B1(_0971_),
    .B2(_0972_),
    .ZN(_0139_));
 OAI21_X1 _3131_ (.A(_0914_),
    .B1(_0537_),
    .B2(_0912_),
    .ZN(_0973_));
 NAND2_X1 _3132_ (.A1(\transfer_count[2][30] ),
    .A2(_0973_),
    .ZN(_0974_));
 NAND3_X1 _3133_ (.A1(_0524_),
    .A2(_0923_),
    .A3(_0537_),
    .ZN(_0975_));
 NAND2_X1 _3134_ (.A1(_0974_),
    .A2(_0975_),
    .ZN(_0140_));
 NOR2_X1 _3135_ (.A1(\transfer_count[2][31] ),
    .A2(_0912_),
    .ZN(_0976_));
 OAI21_X1 _3136_ (.A(_0913_),
    .B1(_0527_),
    .B2(_0518_),
    .ZN(_0977_));
 AOI22_X1 _3137_ (.A1(_0527_),
    .A2(_0976_),
    .B1(_0977_),
    .B2(\transfer_count[2][31] ),
    .ZN(_0978_));
 INV_X1 _3138_ (.A(_0978_),
    .ZN(_0141_));
 NAND3_X1 _3139_ (.A1(_1098_),
    .A2(_1207_),
    .A3(_0691_),
    .ZN(_0979_));
 OAI21_X1 _3140_ (.A(_0979_),
    .B1(_1474_),
    .B2(_0693_),
    .ZN(_0980_));
 AND2_X1 _3141_ (.A1(_0372_),
    .A2(_0980_),
    .ZN(_0142_));
 AOI21_X1 _3142_ (.A(_1181_),
    .B1(_0354_),
    .B2(_1099_),
    .ZN(_0981_));
 AOI21_X1 _3143_ (.A(_0981_),
    .B1(_1489_),
    .B2(_0515_),
    .ZN(_0143_));
 NAND3_X1 _3144_ (.A1(_1097_),
    .A2(_1207_),
    .A3(_0691_),
    .ZN(_0982_));
 OAI21_X1 _3145_ (.A(_0982_),
    .B1(_0693_),
    .B2(_1486_),
    .ZN(_0983_));
 AND2_X1 _3146_ (.A1(_0372_),
    .A2(_0983_),
    .ZN(_0144_));
 NAND3_X1 _3147_ (.A1(\transfer_count[2][6] ),
    .A2(_1207_),
    .A3(_0691_),
    .ZN(_0984_));
 OAI21_X1 _3148_ (.A(_0984_),
    .B1(_1483_),
    .B2(_0693_),
    .ZN(_0985_));
 AND2_X1 _3149_ (.A1(_0372_),
    .A2(_0985_),
    .ZN(_0145_));
 INV_X1 _3150_ (.A(_1108_),
    .ZN(_0986_));
 OAI22_X1 _3151_ (.A1(_0693_),
    .A2(_1480_),
    .B1(_0915_),
    .B2(_0986_),
    .ZN(_0987_));
 AND2_X1 _3152_ (.A1(_0372_),
    .A2(_0987_),
    .ZN(_0146_));
 OAI21_X1 _3153_ (.A(_0915_),
    .B1(_0536_),
    .B2(_0691_),
    .ZN(_0988_));
 NOR2_X1 _3154_ (.A1(_1112_),
    .A2(_0691_),
    .ZN(_0989_));
 AOI22_X1 _3155_ (.A1(_1112_),
    .A2(_0988_),
    .B1(_0989_),
    .B2(_0536_),
    .ZN(_0990_));
 NOR2_X1 _3156_ (.A1(_0219_),
    .A2(_0990_),
    .ZN(_0147_));
 OAI22_X1 _3157_ (.A1(_1510_),
    .A2(_0693_),
    .B1(_0915_),
    .B2(_1111_),
    .ZN(_0991_));
 AND2_X1 _3158_ (.A1(_0372_),
    .A2(_0991_),
    .ZN(_0148_));
 CLKBUF_X3 _3159_ (.A(_0492_),
    .Z(_0992_));
 NAND2_X1 _3160_ (.A1(_1763_),
    .A2(_0992_),
    .ZN(_0993_));
 NAND3_X1 _3161_ (.A1(\transfer_count[3][0] ),
    .A2(_0697_),
    .A3(_0503_),
    .ZN(_0994_));
 AOI21_X1 _3162_ (.A(_0893_),
    .B1(_0993_),
    .B2(_0994_),
    .ZN(_0149_));
 NOR2_X4 _3163_ (.A1(_0492_),
    .A2(_0508_),
    .ZN(_0995_));
 CLKBUF_X3 _3164_ (.A(_0995_),
    .Z(_0996_));
 AOI21_X1 _3165_ (.A(_0695_),
    .B1(_0626_),
    .B2(_0400_),
    .ZN(_0997_));
 OAI21_X1 _3166_ (.A(_0399_),
    .B1(_0996_),
    .B2(_0997_),
    .ZN(_0998_));
 CLKBUF_X3 _3167_ (.A(_0438_),
    .Z(_0999_));
 OR3_X1 _3168_ (.A1(_0399_),
    .A2(_0999_),
    .A3(_0630_),
    .ZN(_1000_));
 AOI21_X1 _3169_ (.A(_0893_),
    .B1(_0998_),
    .B2(_1000_),
    .ZN(_0150_));
 AND2_X1 _3170_ (.A1(_0992_),
    .A2(_0629_),
    .ZN(_1001_));
 OAI21_X1 _3171_ (.A(_0398_),
    .B1(_0996_),
    .B2(_1001_),
    .ZN(_1002_));
 OR3_X1 _3172_ (.A1(_0398_),
    .A2(_0999_),
    .A3(_0629_),
    .ZN(_1003_));
 AOI21_X1 _3173_ (.A(_0893_),
    .B1(_1002_),
    .B2(_1003_),
    .ZN(_0151_));
 AND2_X1 _3174_ (.A1(_0992_),
    .A2(_0628_),
    .ZN(_1004_));
 OAI21_X1 _3175_ (.A(\transfer_count[3][12] ),
    .B1(_0996_),
    .B2(_1004_),
    .ZN(_1005_));
 OR3_X1 _3176_ (.A1(\transfer_count[3][12] ),
    .A2(_0999_),
    .A3(_0628_),
    .ZN(_1006_));
 AOI21_X1 _3177_ (.A(_0893_),
    .B1(_1005_),
    .B2(_1006_),
    .ZN(_0152_));
 AOI21_X1 _3178_ (.A(_0999_),
    .B1(_0406_),
    .B2(_0401_),
    .ZN(_1007_));
 OAI21_X1 _3179_ (.A(_0397_),
    .B1(_0996_),
    .B2(_1007_),
    .ZN(_1008_));
 OR3_X1 _3180_ (.A1(_0397_),
    .A2(_0407_),
    .A3(_0999_),
    .ZN(_1009_));
 AOI21_X1 _3181_ (.A(_1206_),
    .B1(_1008_),
    .B2(_1009_),
    .ZN(_0153_));
 BUF_X2 _3182_ (.A(_0493_),
    .Z(_1010_));
 OR3_X1 _3183_ (.A1(\transfer_count[3][14] ),
    .A2(_1010_),
    .A3(_0627_),
    .ZN(_1011_));
 AOI22_X1 _3184_ (.A1(_0498_),
    .A2(_0627_),
    .B1(_0996_),
    .B2(_1089_),
    .ZN(_1012_));
 OAI21_X1 _3185_ (.A(_1011_),
    .B1(_1012_),
    .B2(_0625_),
    .ZN(_0154_));
 AOI21_X1 _3186_ (.A(\transfer_count[3][15] ),
    .B1(_0992_),
    .B2(_0624_),
    .ZN(_1013_));
 INV_X1 _3187_ (.A(\transfer_count[3][15] ),
    .ZN(_1014_));
 NOR2_X1 _3188_ (.A1(_0438_),
    .A2(_0624_),
    .ZN(_1015_));
 NOR3_X1 _3189_ (.A1(_1014_),
    .A2(_0995_),
    .A3(_1015_),
    .ZN(_1016_));
 NOR3_X1 _3190_ (.A1(_0219_),
    .A2(_1013_),
    .A3(_1016_),
    .ZN(_0155_));
 AND2_X1 _3191_ (.A1(_0992_),
    .A2(_0656_),
    .ZN(_1017_));
 NAND2_X2 _3192_ (.A1(_0438_),
    .A2(_0503_),
    .ZN(_1018_));
 NAND2_X1 _3193_ (.A1(_0421_),
    .A2(_1018_),
    .ZN(_1019_));
 NOR2_X1 _3194_ (.A1(_0697_),
    .A2(_0656_),
    .ZN(_1020_));
 OAI221_X1 _3195_ (.A(_0677_),
    .B1(_0421_),
    .B2(_1017_),
    .C1(_1019_),
    .C2(_1020_),
    .ZN(_1021_));
 INV_X1 _3196_ (.A(_1021_),
    .ZN(_0156_));
 OAI21_X1 _3197_ (.A(_1018_),
    .B1(_0695_),
    .B2(_0431_),
    .ZN(_1022_));
 NOR2_X1 _3198_ (.A1(_0418_),
    .A2(_0695_),
    .ZN(_1023_));
 AOI22_X1 _3199_ (.A1(_0418_),
    .A2(_1022_),
    .B1(_1023_),
    .B2(_0431_),
    .ZN(_1024_));
 NOR2_X1 _3200_ (.A1(_0219_),
    .A2(_1024_),
    .ZN(_0157_));
 NAND4_X1 _3201_ (.A1(_0653_),
    .A2(_0418_),
    .A3(_0498_),
    .A4(_0654_),
    .ZN(_1025_));
 AOI22_X1 _3202_ (.A1(_0498_),
    .A2(_0655_),
    .B1(_0996_),
    .B2(_1089_),
    .ZN(_1026_));
 OAI21_X1 _3203_ (.A(_1025_),
    .B1(_1026_),
    .B2(_0653_),
    .ZN(_0158_));
 NAND2_X2 _3204_ (.A1(_1088_),
    .A2(_0995_),
    .ZN(_1027_));
 OAI21_X1 _3205_ (.A(_1027_),
    .B1(_0652_),
    .B2(_1010_),
    .ZN(_1028_));
 NOR2_X1 _3206_ (.A1(_0417_),
    .A2(_1010_),
    .ZN(_1029_));
 AOI22_X1 _3207_ (.A1(_0417_),
    .A2(_1028_),
    .B1(_1029_),
    .B2(_0652_),
    .ZN(_1030_));
 INV_X1 _3208_ (.A(_1030_),
    .ZN(_0159_));
 NAND2_X1 _3209_ (.A1(_1767_),
    .A2(_0992_),
    .ZN(_1031_));
 NAND3_X1 _3210_ (.A1(\transfer_count[3][1] ),
    .A2(_0697_),
    .A3(_0503_),
    .ZN(_1032_));
 AOI21_X1 _3211_ (.A(_1206_),
    .B1(_1031_),
    .B2(_1032_),
    .ZN(_0160_));
 AND2_X1 _3212_ (.A1(_0992_),
    .A2(_0651_),
    .ZN(_1033_));
 OAI21_X1 _3213_ (.A(_0416_),
    .B1(_0996_),
    .B2(_1033_),
    .ZN(_1034_));
 OR3_X1 _3214_ (.A1(_0416_),
    .A2(_0999_),
    .A3(_0651_),
    .ZN(_1035_));
 AOI21_X1 _3215_ (.A(_1206_),
    .B1(_1034_),
    .B2(_1035_),
    .ZN(_0161_));
 OAI21_X1 _3216_ (.A(_1027_),
    .B1(_1010_),
    .B2(_0429_),
    .ZN(_1036_));
 NOR2_X1 _3217_ (.A1(_0415_),
    .A2(_1010_),
    .ZN(_1037_));
 AOI22_X1 _3218_ (.A1(_0415_),
    .A2(_1036_),
    .B1(_1037_),
    .B2(_0429_),
    .ZN(_1038_));
 INV_X1 _3219_ (.A(_1038_),
    .ZN(_0162_));
 OAI21_X1 _3220_ (.A(_1027_),
    .B1(_0650_),
    .B2(_1010_),
    .ZN(_1039_));
 NAND2_X1 _3221_ (.A1(_0414_),
    .A2(_1039_),
    .ZN(_1040_));
 NAND2_X1 _3222_ (.A1(_0498_),
    .A2(_0650_),
    .ZN(_1041_));
 OAI21_X1 _3223_ (.A(_1040_),
    .B1(_1041_),
    .B2(_0414_),
    .ZN(_0163_));
 OAI21_X1 _3224_ (.A(_1018_),
    .B1(_0697_),
    .B2(_0634_),
    .ZN(_1042_));
 NAND2_X1 _3225_ (.A1(_0408_),
    .A2(_1042_),
    .ZN(_1043_));
 INV_X1 _3226_ (.A(_0408_),
    .ZN(_1044_));
 NAND3_X1 _3227_ (.A1(_1044_),
    .A2(_0424_),
    .A3(_0992_),
    .ZN(_1045_));
 AOI21_X1 _3228_ (.A(_1206_),
    .B1(_1043_),
    .B2(_1045_),
    .ZN(_0164_));
 AOI221_X1 _3229_ (.A(_0646_),
    .B1(_0439_),
    .B2(_0647_),
    .C1(_0995_),
    .C2(_1088_),
    .ZN(_1046_));
 NAND3_X1 _3230_ (.A1(_0408_),
    .A2(_0498_),
    .A3(_0639_),
    .ZN(_1047_));
 AOI21_X1 _3231_ (.A(_1046_),
    .B1(_1047_),
    .B2(_0646_),
    .ZN(_0165_));
 NAND4_X1 _3232_ (.A1(_0426_),
    .A2(_0409_),
    .A3(_0424_),
    .A4(_0498_),
    .ZN(_1048_));
 AOI22_X1 _3233_ (.A1(_0427_),
    .A2(_0498_),
    .B1(_0996_),
    .B2(_1089_),
    .ZN(_1049_));
 OAI21_X1 _3234_ (.A(_1048_),
    .B1(_1049_),
    .B2(_0426_),
    .ZN(_0166_));
 AOI221_X1 _3235_ (.A(_0644_),
    .B1(_0439_),
    .B2(_0645_),
    .C1(_0995_),
    .C2(_1088_),
    .ZN(_1050_));
 OR2_X1 _3236_ (.A1(_1010_),
    .A2(_0645_),
    .ZN(_1051_));
 AOI21_X1 _3237_ (.A(_1050_),
    .B1(_1051_),
    .B2(_0644_),
    .ZN(_0167_));
 NAND4_X1 _3238_ (.A1(_0409_),
    .A2(_0410_),
    .A3(_0634_),
    .A4(_1018_),
    .ZN(_1052_));
 NAND2_X1 _3239_ (.A1(_0697_),
    .A2(_0508_),
    .ZN(_1053_));
 NAND3_X1 _3240_ (.A1(\transfer_count[3][27] ),
    .A2(_1052_),
    .A3(_1053_),
    .ZN(_1054_));
 OR3_X1 _3241_ (.A1(\transfer_count[3][27] ),
    .A2(_0999_),
    .A3(_0643_),
    .ZN(_1055_));
 AOI21_X1 _3242_ (.A(_1206_),
    .B1(_1054_),
    .B2(_1055_),
    .ZN(_0168_));
 OR3_X1 _3243_ (.A1(\transfer_count[3][28] ),
    .A2(_1010_),
    .A3(_0642_),
    .ZN(_1056_));
 AOI22_X1 _3244_ (.A1(_0498_),
    .A2(_0642_),
    .B1(_0995_),
    .B2(_1089_),
    .ZN(_1057_));
 OAI21_X1 _3245_ (.A(_1056_),
    .B1(_1057_),
    .B2(_0641_),
    .ZN(_0169_));
 AND2_X1 _3246_ (.A1(_0425_),
    .A2(_0439_),
    .ZN(_1058_));
 OAI21_X1 _3247_ (.A(_1027_),
    .B1(_1010_),
    .B2(_0425_),
    .ZN(_1059_));
 MUX2_X1 _3248_ (.A(_1058_),
    .B(_1059_),
    .S(\transfer_count[3][29] ),
    .Z(_0170_));
 NOR2_X1 _3249_ (.A1(_0619_),
    .A2(_0695_),
    .ZN(_1060_));
 OAI21_X1 _3250_ (.A(_0393_),
    .B1(_0996_),
    .B2(_1060_),
    .ZN(_1061_));
 INV_X1 _3251_ (.A(_0393_),
    .ZN(_1062_));
 NAND3_X1 _3252_ (.A1(_1062_),
    .A2(_0619_),
    .A3(_0992_),
    .ZN(_1063_));
 AOI21_X1 _3253_ (.A(_1206_),
    .B1(_1061_),
    .B2(_1063_),
    .ZN(_0171_));
 OR3_X1 _3254_ (.A1(\transfer_count[3][30] ),
    .A2(_0493_),
    .A3(_0640_),
    .ZN(_1064_));
 AOI22_X1 _3255_ (.A1(_0498_),
    .A2(_0640_),
    .B1(_0995_),
    .B2(_1089_),
    .ZN(_1065_));
 OAI21_X1 _3256_ (.A(_1064_),
    .B1(_1065_),
    .B2(_0637_),
    .ZN(_0172_));
 AOI221_X1 _3257_ (.A(_0633_),
    .B1(_0439_),
    .B2(_0636_),
    .C1(_0995_),
    .C2(_1088_),
    .ZN(_1066_));
 OR2_X1 _3258_ (.A1(_1010_),
    .A2(_0636_),
    .ZN(_1067_));
 AOI21_X1 _3259_ (.A(_1066_),
    .B1(_1067_),
    .B2(_0633_),
    .ZN(_0173_));
 NOR3_X1 _3260_ (.A1(_0391_),
    .A2(_0412_),
    .A3(_0999_),
    .ZN(_1068_));
 OAI21_X1 _3261_ (.A(_1018_),
    .B1(_0695_),
    .B2(_0395_),
    .ZN(_1069_));
 AOI21_X1 _3262_ (.A(_1068_),
    .B1(_1069_),
    .B2(_0391_),
    .ZN(_1070_));
 NOR2_X1 _3263_ (.A1(_0219_),
    .A2(_1070_),
    .ZN(_0174_));
 AOI21_X1 _3264_ (.A(_0999_),
    .B1(_0621_),
    .B2(_0391_),
    .ZN(_1071_));
 OAI21_X1 _3265_ (.A(_0392_),
    .B1(_0996_),
    .B2(_1071_),
    .ZN(_1072_));
 OR3_X1 _3266_ (.A1(_0392_),
    .A2(_0999_),
    .A3(_0623_),
    .ZN(_1073_));
 AOI21_X1 _3267_ (.A(_1206_),
    .B1(_1072_),
    .B2(_1073_),
    .ZN(_0175_));
 NAND3_X1 _3268_ (.A1(_0390_),
    .A2(_0695_),
    .A3(_0503_),
    .ZN(_1074_));
 OAI21_X1 _3269_ (.A(_1074_),
    .B1(_0697_),
    .B2(_1783_),
    .ZN(_1075_));
 AND2_X1 _3270_ (.A1(_0372_),
    .A2(_1075_),
    .ZN(_0176_));
 NAND3_X1 _3271_ (.A1(\transfer_count[3][6] ),
    .A2(_0695_),
    .A3(_0503_),
    .ZN(_1076_));
 OAI21_X1 _3272_ (.A(_1076_),
    .B1(_1780_),
    .B2(_0697_),
    .ZN(_1077_));
 AND2_X1 _3273_ (.A1(_0372_),
    .A2(_1077_),
    .ZN(_0177_));
 NAND3_X1 _3274_ (.A1(_0402_),
    .A2(_0695_),
    .A3(_0503_),
    .ZN(_1078_));
 OAI21_X1 _3275_ (.A(_1078_),
    .B1(_1777_),
    .B2(_0697_),
    .ZN(_1079_));
 AND2_X1 _3276_ (.A1(_0372_),
    .A2(_1079_),
    .ZN(_0178_));
 AOI21_X1 _3277_ (.A(_0995_),
    .B1(_0632_),
    .B2(_0992_),
    .ZN(_1080_));
 NOR2_X1 _3278_ (.A1(_0631_),
    .A2(_1080_),
    .ZN(_1081_));
 NOR3_X1 _3279_ (.A1(_0403_),
    .A2(_0697_),
    .A3(_0632_),
    .ZN(_1082_));
 OAI21_X1 _3280_ (.A(_0380_),
    .B1(_1081_),
    .B2(_1082_),
    .ZN(_1083_));
 INV_X1 _3281_ (.A(_1083_),
    .ZN(_0179_));
 NOR3_X1 _3282_ (.A1(_0400_),
    .A2(_0430_),
    .A3(_0438_),
    .ZN(_1084_));
 OAI21_X1 _3283_ (.A(_1018_),
    .B1(_0695_),
    .B2(_0406_),
    .ZN(_1085_));
 AOI21_X1 _3284_ (.A(_1084_),
    .B1(_1085_),
    .B2(_0400_),
    .ZN(_1086_));
 NOR2_X1 _3285_ (.A1(_0219_),
    .A2(_1086_),
    .ZN(_0180_));
 HA_X1 _3286_ (.A(_1465_),
    .B(_1466_),
    .CO(_1467_),
    .S(_1468_));
 HA_X1 _3287_ (.A(\transfer_count[2][0] ),
    .B(\transfer_count[2][1] ),
    .CO(_1469_),
    .S(_1470_));
 HA_X1 _3288_ (.A(net90),
    .B(_1471_),
    .CO(_1472_),
    .S(_1473_));
 HA_X1 _3289_ (.A(net92),
    .B(_1474_),
    .CO(_1475_),
    .S(_1476_));
 HA_X1 _3290_ (.A(net91),
    .B(_1477_),
    .CO(_1478_),
    .S(_1479_));
 HA_X1 _3291_ (.A(net97),
    .B(_1480_),
    .CO(_1481_),
    .S(_1482_));
 HA_X1 _3292_ (.A(net96),
    .B(_1483_),
    .CO(_1484_),
    .S(_1485_));
 HA_X1 _3293_ (.A(net94),
    .B(_1486_),
    .CO(_1487_),
    .S(_1488_));
 HA_X1 _3294_ (.A(net93),
    .B(_1489_),
    .CO(_1490_),
    .S(_1491_));
 HA_X1 _3295_ (.A(net105),
    .B(_1492_),
    .CO(_1493_),
    .S(_1494_));
 HA_X1 _3296_ (.A(_1495_),
    .B(net104),
    .CO(_1496_),
    .S(_1497_));
 HA_X1 _3297_ (.A(_1498_),
    .B(net103),
    .CO(_1499_),
    .S(_1500_));
 HA_X1 _3298_ (.A(_1501_),
    .B(net102),
    .CO(_1502_),
    .S(_1503_));
 HA_X1 _3299_ (.A(net101),
    .B(_1504_),
    .CO(_1505_),
    .S(_1506_));
 HA_X1 _3300_ (.A(net100),
    .B(_1507_),
    .CO(_1508_),
    .S(_1509_));
 HA_X1 _3301_ (.A(net99),
    .B(_1510_),
    .CO(_1511_),
    .S(_1512_));
 HA_X1 _3302_ (.A(net98),
    .B(_1513_),
    .CO(_1514_),
    .S(_1515_));
 HA_X1 _3303_ (.A(net123),
    .B(_1516_),
    .CO(_1517_),
    .S(_1518_));
 HA_X1 _3304_ (.A(net122),
    .B(_1519_),
    .CO(_1520_),
    .S(_1521_));
 HA_X1 _3305_ (.A(net121),
    .B(_1522_),
    .CO(_1523_),
    .S(_1524_));
 HA_X1 _3306_ (.A(net120),
    .B(_1525_),
    .CO(_1526_),
    .S(_1527_));
 HA_X1 _3307_ (.A(net119),
    .B(_1528_),
    .CO(_1529_),
    .S(_1530_));
 HA_X1 _3308_ (.A(net118),
    .B(_1531_),
    .CO(_1532_),
    .S(_1533_));
 HA_X1 _3309_ (.A(net116),
    .B(_1534_),
    .CO(_1535_),
    .S(_1536_));
 HA_X1 _3310_ (.A(net115),
    .B(_1537_),
    .CO(_1538_),
    .S(_1539_));
 HA_X1 _3311_ (.A(net114),
    .B(_1540_),
    .CO(_1541_),
    .S(_1542_));
 HA_X1 _3312_ (.A(net113),
    .B(_1543_),
    .CO(_1544_),
    .S(_1545_));
 HA_X1 _3313_ (.A(net112),
    .B(_1546_),
    .CO(_1547_),
    .S(_1548_));
 HA_X1 _3314_ (.A(net111),
    .B(_1549_),
    .CO(_1550_),
    .S(_1551_));
 HA_X1 _3315_ (.A(net110),
    .B(_1552_),
    .CO(_1553_),
    .S(_1554_));
 HA_X1 _3316_ (.A(net109),
    .B(_1555_),
    .CO(_1556_),
    .S(_1557_));
 HA_X1 _3317_ (.A(net108),
    .B(_1558_),
    .CO(_1559_),
    .S(_1560_));
 HA_X1 _3318_ (.A(net107),
    .B(_1561_),
    .CO(_1562_),
    .S(_1563_));
 HA_X1 _3319_ (.A(net88),
    .B(_1564_),
    .CO(_1565_),
    .S(_1566_));
 HA_X1 _3320_ (.A(net87),
    .B(_1567_),
    .CO(_1568_),
    .S(_1569_));
 HA_X1 _3321_ (.A(net86),
    .B(_1570_),
    .CO(_1571_),
    .S(_1572_));
 HA_X1 _3322_ (.A(net85),
    .B(_1573_),
    .CO(_1574_),
    .S(_1575_));
 HA_X1 _3323_ (.A(net83),
    .B(_1576_),
    .CO(_1577_),
    .S(_1578_));
 HA_X1 _3324_ (.A(net82),
    .B(_1579_),
    .CO(_1580_),
    .S(_1581_));
 HA_X1 _3325_ (.A(net81),
    .B(_1582_),
    .CO(_1583_),
    .S(_1584_));
 HA_X1 _3326_ (.A(net80),
    .B(_1585_),
    .CO(_1586_),
    .S(_1587_));
 HA_X1 _3327_ (.A(net79),
    .B(_1588_),
    .CO(_1589_),
    .S(_1590_));
 HA_X1 _3328_ (.A(net78),
    .B(_1591_),
    .CO(_1592_),
    .S(_1593_));
 HA_X1 _3329_ (.A(net77),
    .B(_1594_),
    .CO(_1595_),
    .S(_1596_));
 HA_X1 _3330_ (.A(net76),
    .B(_1597_),
    .CO(_1598_),
    .S(_1599_));
 HA_X1 _3331_ (.A(net75),
    .B(_1600_),
    .CO(_1601_),
    .S(_1602_));
 HA_X1 _3332_ (.A(net74),
    .B(_1603_),
    .CO(_1604_),
    .S(_1605_));
 HA_X1 _3333_ (.A(net72),
    .B(_1606_),
    .CO(_1607_),
    .S(_1608_));
 HA_X1 _3334_ (.A(net71),
    .B(_1609_),
    .CO(_1610_),
    .S(_1611_));
 HA_X1 _3335_ (.A(net70),
    .B(_1612_),
    .CO(_1613_),
    .S(_1614_));
 HA_X1 _3336_ (.A(net69),
    .B(_1615_),
    .CO(_1616_),
    .S(_1617_));
 HA_X1 _3337_ (.A(net68),
    .B(_1618_),
    .CO(_1619_),
    .S(_1620_));
 HA_X1 _3338_ (.A(net67),
    .B(_1621_),
    .CO(_1622_),
    .S(_1623_));
 HA_X1 _3339_ (.A(net66),
    .B(_1624_),
    .CO(_1625_),
    .S(_1626_));
 HA_X1 _3340_ (.A(net65),
    .B(_1627_),
    .CO(_1628_),
    .S(_1629_));
 HA_X1 _3341_ (.A(net64),
    .B(_1630_),
    .CO(_1631_),
    .S(_1632_));
 HA_X1 _3342_ (.A(net63),
    .B(_1633_),
    .CO(_1634_),
    .S(_1635_));
 HA_X1 _3343_ (.A(net61),
    .B(_1636_),
    .CO(_1637_),
    .S(_1638_));
 HA_X1 _3344_ (.A(net60),
    .B(_1639_),
    .CO(_1640_),
    .S(_1641_));
 HA_X1 _3345_ (.A(net59),
    .B(_1642_),
    .CO(_1643_),
    .S(_1644_));
 HA_X1 _3346_ (.A(net58),
    .B(_1645_),
    .CO(_1646_),
    .S(_1647_));
 HA_X1 _3347_ (.A(net57),
    .B(_1648_),
    .CO(_1649_),
    .S(_1650_));
 HA_X1 _3348_ (.A(net56),
    .B(_1651_),
    .CO(_1652_),
    .S(_1653_));
 HA_X1 _3349_ (.A(\transfer_count[1][0] ),
    .B(\transfer_count[1][1] ),
    .CO(_1654_),
    .S(_1655_));
 HA_X1 _3350_ (.A(net55),
    .B(_1656_),
    .CO(_1657_),
    .S(_1658_));
 HA_X1 _3351_ (.A(_1659_),
    .B(_1660_),
    .CO(_1661_),
    .S(_1662_));
 HA_X1 _3352_ (.A(net53),
    .B(_1663_),
    .CO(_1664_),
    .S(_1665_));
 HA_X1 _3353_ (.A(net52),
    .B(_1666_),
    .CO(_1667_),
    .S(_1668_));
 HA_X1 _3354_ (.A(net50),
    .B(_1669_),
    .CO(_1670_),
    .S(_1671_));
 HA_X1 _3355_ (.A(net49),
    .B(_1672_),
    .CO(_1673_),
    .S(_1674_));
 HA_X1 _3356_ (.A(net48),
    .B(_1675_),
    .CO(_1676_),
    .S(_1677_));
 HA_X1 _3357_ (.A(net47),
    .B(_1678_),
    .CO(_1679_),
    .S(_1680_));
 HA_X1 _3358_ (.A(net46),
    .B(_1681_),
    .CO(_1682_),
    .S(_1683_));
 HA_X1 _3359_ (.A(net45),
    .B(_1684_),
    .CO(_1685_),
    .S(_1686_));
 HA_X1 _3360_ (.A(net44),
    .B(_1687_),
    .CO(_1688_),
    .S(_1689_));
 HA_X1 _3361_ (.A(net43),
    .B(_1690_),
    .CO(_1691_),
    .S(_1692_));
 HA_X1 _3362_ (.A(net42),
    .B(_1693_),
    .CO(_1694_),
    .S(_1695_));
 HA_X1 _3363_ (.A(net41),
    .B(_1696_),
    .CO(_1697_),
    .S(_1698_));
 HA_X1 _3364_ (.A(net39),
    .B(_1699_),
    .CO(_1700_),
    .S(_1701_));
 HA_X1 _3365_ (.A(net38),
    .B(_1702_),
    .CO(_1703_),
    .S(_1704_));
 HA_X1 _3366_ (.A(net37),
    .B(_1705_),
    .CO(_1706_),
    .S(_1707_));
 HA_X1 _3367_ (.A(net36),
    .B(_1708_),
    .CO(_1709_),
    .S(_1710_));
 HA_X1 _3368_ (.A(net35),
    .B(_1711_),
    .CO(_1712_),
    .S(_1713_));
 HA_X1 _3369_ (.A(net34),
    .B(_1714_),
    .CO(_1715_),
    .S(_1716_));
 HA_X1 _3370_ (.A(net33),
    .B(_1717_),
    .CO(_1718_),
    .S(_1719_));
 HA_X1 _3371_ (.A(net32),
    .B(_1720_),
    .CO(_1721_),
    .S(_1722_));
 HA_X1 _3372_ (.A(net23),
    .B(_1723_),
    .CO(_1724_),
    .S(_1725_));
 HA_X1 _3373_ (.A(net12),
    .B(_1726_),
    .CO(_1727_),
    .S(_1728_));
 HA_X1 _3374_ (.A(net128),
    .B(_1729_),
    .CO(_1730_),
    .S(_1731_));
 HA_X1 _3375_ (.A(net117),
    .B(_1732_),
    .CO(_1733_),
    .S(_1734_));
 HA_X1 _3376_ (.A(net106),
    .B(_1735_),
    .CO(_1736_),
    .S(_1737_));
 HA_X1 _3377_ (.A(net95),
    .B(_1738_),
    .CO(_1739_),
    .S(_1740_));
 HA_X1 _3378_ (.A(net84),
    .B(_1741_),
    .CO(_1742_),
    .S(_1743_));
 HA_X1 _3379_ (.A(net73),
    .B(_1744_),
    .CO(_1745_),
    .S(_1746_));
 HA_X1 _3380_ (.A(net62),
    .B(_1747_),
    .CO(_1748_),
    .S(_1749_));
 HA_X1 _3381_ (.A(net51),
    .B(_1750_),
    .CO(_1751_),
    .S(_1752_));
 HA_X1 _3382_ (.A(\transfer_count[0][0] ),
    .B(\transfer_count[0][1] ),
    .CO(_1753_),
    .S(_1754_));
 HA_X1 _3383_ (.A(net40),
    .B(_1755_),
    .CO(_1756_),
    .S(_1757_));
 HA_X1 _3384_ (.A(_1758_),
    .B(_1759_),
    .CO(_1760_),
    .S(_1761_));
 HA_X1 _3385_ (.A(_1762_),
    .B(_1763_),
    .CO(_1764_),
    .S(_1765_));
 HA_X1 _3386_ (.A(\transfer_count[3][0] ),
    .B(\transfer_count[3][1] ),
    .CO(_1766_),
    .S(_1767_));
 HA_X1 _3387_ (.A(net125),
    .B(_1768_),
    .CO(_1769_),
    .S(_1770_));
 HA_X1 _3388_ (.A(net127),
    .B(_1771_),
    .CO(_1772_),
    .S(_1773_));
 HA_X1 _3389_ (.A(net126),
    .B(_1774_),
    .CO(_1775_),
    .S(_1776_));
 HA_X1 _3390_ (.A(net5),
    .B(_1777_),
    .CO(_1778_),
    .S(_1779_));
 HA_X1 _3391_ (.A(net4),
    .B(_1780_),
    .CO(_1781_),
    .S(_1782_));
 HA_X1 _3392_ (.A(net3),
    .B(_1783_),
    .CO(_1784_),
    .S(_1785_));
 HA_X1 _3393_ (.A(net2),
    .B(_1786_),
    .CO(_1787_),
    .S(_1788_));
 HA_X1 _3394_ (.A(net14),
    .B(_1789_),
    .CO(_1790_),
    .S(_1791_));
 HA_X1 _3395_ (.A(net13),
    .B(_1792_),
    .CO(_1793_),
    .S(_1794_));
 HA_X1 _3396_ (.A(net11),
    .B(_1795_),
    .CO(_1796_),
    .S(_1797_));
 HA_X1 _3397_ (.A(net10),
    .B(_1798_),
    .CO(_1799_),
    .S(_1800_));
 HA_X1 _3398_ (.A(net9),
    .B(_1801_),
    .CO(_1802_),
    .S(_1803_));
 HA_X1 _3399_ (.A(net8),
    .B(_1804_),
    .CO(_1805_),
    .S(_1806_));
 HA_X1 _3400_ (.A(net7),
    .B(_1807_),
    .CO(_1808_),
    .S(_1809_));
 HA_X1 _3401_ (.A(net6),
    .B(_1810_),
    .CO(_1811_),
    .S(_1812_));
 HA_X1 _3402_ (.A(net31),
    .B(_1813_),
    .CO(_1814_),
    .S(_1815_));
 HA_X1 _3403_ (.A(net30),
    .B(_1816_),
    .CO(_1817_),
    .S(_1818_));
 HA_X1 _3404_ (.A(net29),
    .B(_1819_),
    .CO(_1820_),
    .S(_1821_));
 HA_X1 _3405_ (.A(net28),
    .B(_1822_),
    .CO(_1823_),
    .S(_1824_));
 HA_X1 _3406_ (.A(net27),
    .B(_1825_),
    .CO(_1826_),
    .S(_1827_));
 HA_X1 _3407_ (.A(net26),
    .B(_1828_),
    .CO(_1829_),
    .S(_1830_));
 HA_X1 _3408_ (.A(net25),
    .B(_1831_),
    .CO(_1832_),
    .S(_1833_));
 HA_X1 _3409_ (.A(net24),
    .B(_1834_),
    .CO(_1835_),
    .S(_1836_));
 HA_X1 _3410_ (.A(net22),
    .B(_1837_),
    .CO(_1838_),
    .S(_1839_));
 HA_X1 _3411_ (.A(net21),
    .B(_1840_),
    .CO(_1841_),
    .S(_1842_));
 HA_X1 _3412_ (.A(net20),
    .B(_1843_),
    .CO(_1844_),
    .S(_1845_));
 HA_X1 _3413_ (.A(net19),
    .B(_1846_),
    .CO(_1847_),
    .S(_1848_));
 HA_X1 _3414_ (.A(net18),
    .B(_1849_),
    .CO(_1850_),
    .S(_1851_));
 HA_X1 _3415_ (.A(net17),
    .B(_1852_),
    .CO(_1853_),
    .S(_1854_));
 HA_X1 _3416_ (.A(net16),
    .B(_1855_),
    .CO(_1856_),
    .S(_1857_));
 HA_X1 _3417_ (.A(net15),
    .B(_1858_),
    .CO(_1859_),
    .S(_1860_));
 HA_X1 _3418_ (.A(_1861_),
    .B(_1862_),
    .CO(_1863_),
    .S(_1864_));
 HA_X1 _3419_ (.A(\active_channel_count[0] ),
    .B(\active_channel_count[1] ),
    .CO(_1865_),
    .S(_1866_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X1 _3421_ (.A(net163),
    .Z(channel_error[0]));
 BUF_X1 _3422_ (.A(net164),
    .Z(channel_error[1]));
 BUF_X1 _3423_ (.A(net165),
    .Z(channel_error[2]));
 BUF_X1 _3424_ (.A(net166),
    .Z(channel_error[3]));
 BUF_X1 _3425_ (.A(net167),
    .Z(debug_channel_state[0]));
 BUF_X1 _3426_ (.A(net168),
    .Z(debug_channel_state[1]));
 BUF_X1 _3427_ (.A(net169),
    .Z(debug_channel_state[2]));
 BUF_X1 _3428_ (.A(net170),
    .Z(debug_channel_state[3]));
 BUF_X1 _3429_ (.A(net171),
    .Z(debug_channel_state[4]));
 BUF_X1 _3430_ (.A(net172),
    .Z(debug_channel_state[5]));
 BUF_X1 _3431_ (.A(net173),
    .Z(debug_channel_state[6]));
 BUF_X1 _3432_ (.A(net174),
    .Z(debug_channel_state[7]));
 BUF_X1 _3433_ (.A(net175),
    .Z(debug_channel_state[8]));
 BUF_X1 _3434_ (.A(net176),
    .Z(debug_channel_state[9]));
 BUF_X1 _3435_ (.A(net177),
    .Z(debug_channel_state[10]));
 BUF_X1 _3436_ (.A(net178),
    .Z(debug_channel_state[11]));
 BUF_X1 _3437_ (.A(net179),
    .Z(debug_transfer_count[0]));
 BUF_X1 _3438_ (.A(net180),
    .Z(debug_transfer_count[1]));
 BUF_X1 _3439_ (.A(net181),
    .Z(debug_transfer_count[2]));
 BUF_X1 _3440_ (.A(net182),
    .Z(debug_transfer_count[3]));
 BUF_X1 _3441_ (.A(net183),
    .Z(debug_transfer_count[4]));
 BUF_X1 _3442_ (.A(net184),
    .Z(debug_transfer_count[5]));
 BUF_X1 _3443_ (.A(net185),
    .Z(debug_transfer_count[6]));
 BUF_X1 _3444_ (.A(net186),
    .Z(debug_transfer_count[7]));
 BUF_X1 _3445_ (.A(net187),
    .Z(debug_transfer_count[8]));
 BUF_X1 _3446_ (.A(net188),
    .Z(debug_transfer_count[9]));
 BUF_X1 _3447_ (.A(net189),
    .Z(debug_transfer_count[10]));
 BUF_X1 _3448_ (.A(net190),
    .Z(debug_transfer_count[11]));
 BUF_X1 _3449_ (.A(net191),
    .Z(debug_transfer_count[12]));
 BUF_X1 _3450_ (.A(net192),
    .Z(debug_transfer_count[13]));
 BUF_X1 _3451_ (.A(net193),
    .Z(debug_transfer_count[14]));
 BUF_X1 _3452_ (.A(net194),
    .Z(debug_transfer_count[15]));
 BUF_X1 _3453_ (.A(net195),
    .Z(debug_transfer_count[16]));
 BUF_X1 _3454_ (.A(net196),
    .Z(debug_transfer_count[17]));
 BUF_X1 _3455_ (.A(net197),
    .Z(debug_transfer_count[18]));
 BUF_X1 _3456_ (.A(net198),
    .Z(debug_transfer_count[19]));
 BUF_X1 _3457_ (.A(net199),
    .Z(debug_transfer_count[20]));
 BUF_X1 _3458_ (.A(net200),
    .Z(debug_transfer_count[21]));
 BUF_X1 _3459_ (.A(net201),
    .Z(debug_transfer_count[22]));
 BUF_X1 _3460_ (.A(net202),
    .Z(debug_transfer_count[23]));
 BUF_X1 _3461_ (.A(net203),
    .Z(debug_transfer_count[24]));
 BUF_X1 _3462_ (.A(net204),
    .Z(debug_transfer_count[25]));
 BUF_X1 _3463_ (.A(net205),
    .Z(debug_transfer_count[26]));
 BUF_X1 _3464_ (.A(net206),
    .Z(debug_transfer_count[27]));
 BUF_X1 _3465_ (.A(net207),
    .Z(debug_transfer_count[28]));
 BUF_X1 _3466_ (.A(net208),
    .Z(debug_transfer_count[29]));
 BUF_X1 _3467_ (.A(net209),
    .Z(debug_transfer_count[30]));
 BUF_X1 _3468_ (.A(net210),
    .Z(debug_transfer_count[31]));
 BUF_X1 _3469_ (.A(net211),
    .Z(debug_transfer_count[32]));
 BUF_X1 _3470_ (.A(net212),
    .Z(debug_transfer_count[33]));
 BUF_X1 _3471_ (.A(net213),
    .Z(debug_transfer_count[34]));
 BUF_X1 _3472_ (.A(net214),
    .Z(debug_transfer_count[35]));
 BUF_X1 _3473_ (.A(net215),
    .Z(debug_transfer_count[36]));
 BUF_X1 _3474_ (.A(net216),
    .Z(debug_transfer_count[37]));
 BUF_X1 _3475_ (.A(net217),
    .Z(debug_transfer_count[38]));
 BUF_X1 _3476_ (.A(net218),
    .Z(debug_transfer_count[39]));
 BUF_X1 _3477_ (.A(net219),
    .Z(debug_transfer_count[40]));
 BUF_X1 _3478_ (.A(net220),
    .Z(debug_transfer_count[41]));
 BUF_X1 _3479_ (.A(net221),
    .Z(debug_transfer_count[42]));
 BUF_X1 _3480_ (.A(net222),
    .Z(debug_transfer_count[43]));
 BUF_X1 _3481_ (.A(net223),
    .Z(debug_transfer_count[44]));
 BUF_X1 _3482_ (.A(net224),
    .Z(debug_transfer_count[45]));
 BUF_X1 _3483_ (.A(net225),
    .Z(debug_transfer_count[46]));
 BUF_X1 _3484_ (.A(net226),
    .Z(debug_transfer_count[47]));
 BUF_X1 _3485_ (.A(net227),
    .Z(debug_transfer_count[48]));
 BUF_X1 _3486_ (.A(net228),
    .Z(debug_transfer_count[49]));
 BUF_X1 _3487_ (.A(net229),
    .Z(debug_transfer_count[50]));
 BUF_X1 _3488_ (.A(net230),
    .Z(debug_transfer_count[51]));
 BUF_X1 _3489_ (.A(net231),
    .Z(debug_transfer_count[52]));
 BUF_X1 _3490_ (.A(net232),
    .Z(debug_transfer_count[53]));
 BUF_X1 _3491_ (.A(net233),
    .Z(debug_transfer_count[54]));
 BUF_X1 _3492_ (.A(net234),
    .Z(debug_transfer_count[55]));
 BUF_X1 _3493_ (.A(net235),
    .Z(debug_transfer_count[56]));
 BUF_X1 _3494_ (.A(net236),
    .Z(debug_transfer_count[57]));
 BUF_X1 _3495_ (.A(net237),
    .Z(debug_transfer_count[58]));
 BUF_X1 _3496_ (.A(net238),
    .Z(debug_transfer_count[59]));
 BUF_X1 _3497_ (.A(net239),
    .Z(debug_transfer_count[60]));
 BUF_X1 _3498_ (.A(net240),
    .Z(debug_transfer_count[61]));
 BUF_X1 _3499_ (.A(net241),
    .Z(debug_transfer_count[62]));
 BUF_X1 _3500_ (.A(net242),
    .Z(debug_transfer_count[63]));
 BUF_X1 _3501_ (.A(net243),
    .Z(debug_transfer_count[64]));
 BUF_X1 _3502_ (.A(net244),
    .Z(debug_transfer_count[65]));
 BUF_X1 _3503_ (.A(net245),
    .Z(debug_transfer_count[66]));
 BUF_X1 _3504_ (.A(net246),
    .Z(debug_transfer_count[67]));
 BUF_X1 _3505_ (.A(net247),
    .Z(debug_transfer_count[68]));
 BUF_X1 _3506_ (.A(net248),
    .Z(debug_transfer_count[69]));
 BUF_X1 _3507_ (.A(net249),
    .Z(debug_transfer_count[70]));
 BUF_X1 _3508_ (.A(net250),
    .Z(debug_transfer_count[71]));
 BUF_X1 _3509_ (.A(net251),
    .Z(debug_transfer_count[72]));
 BUF_X1 _3510_ (.A(net252),
    .Z(debug_transfer_count[73]));
 BUF_X1 _3511_ (.A(net253),
    .Z(debug_transfer_count[74]));
 BUF_X1 _3512_ (.A(net254),
    .Z(debug_transfer_count[75]));
 BUF_X1 _3513_ (.A(net255),
    .Z(debug_transfer_count[76]));
 BUF_X1 _3514_ (.A(net256),
    .Z(debug_transfer_count[77]));
 BUF_X1 _3515_ (.A(net257),
    .Z(debug_transfer_count[78]));
 BUF_X1 _3516_ (.A(net258),
    .Z(debug_transfer_count[79]));
 BUF_X1 _3517_ (.A(net259),
    .Z(debug_transfer_count[80]));
 BUF_X1 _3518_ (.A(net260),
    .Z(debug_transfer_count[81]));
 BUF_X1 _3519_ (.A(net261),
    .Z(debug_transfer_count[82]));
 BUF_X1 _3520_ (.A(net262),
    .Z(debug_transfer_count[83]));
 BUF_X1 _3521_ (.A(net263),
    .Z(debug_transfer_count[84]));
 BUF_X1 _3522_ (.A(net264),
    .Z(debug_transfer_count[85]));
 BUF_X1 _3523_ (.A(net265),
    .Z(debug_transfer_count[86]));
 BUF_X1 _3524_ (.A(net266),
    .Z(debug_transfer_count[87]));
 BUF_X1 _3525_ (.A(net267),
    .Z(debug_transfer_count[88]));
 BUF_X1 _3526_ (.A(net268),
    .Z(debug_transfer_count[89]));
 BUF_X1 _3527_ (.A(net269),
    .Z(debug_transfer_count[90]));
 BUF_X1 _3528_ (.A(net270),
    .Z(debug_transfer_count[91]));
 BUF_X1 _3529_ (.A(net271),
    .Z(debug_transfer_count[92]));
 BUF_X1 _3530_ (.A(net272),
    .Z(debug_transfer_count[93]));
 BUF_X1 _3531_ (.A(net273),
    .Z(debug_transfer_count[94]));
 BUF_X1 _3532_ (.A(net274),
    .Z(debug_transfer_count[95]));
 BUF_X1 _3533_ (.A(net275),
    .Z(debug_transfer_count[96]));
 BUF_X1 _3534_ (.A(net276),
    .Z(debug_transfer_count[97]));
 BUF_X1 _3535_ (.A(net277),
    .Z(debug_transfer_count[98]));
 BUF_X1 _3536_ (.A(net278),
    .Z(debug_transfer_count[99]));
 BUF_X1 _3537_ (.A(net279),
    .Z(debug_transfer_count[100]));
 BUF_X1 _3538_ (.A(net280),
    .Z(debug_transfer_count[101]));
 BUF_X1 _3539_ (.A(net281),
    .Z(debug_transfer_count[102]));
 BUF_X1 _3540_ (.A(net282),
    .Z(debug_transfer_count[103]));
 BUF_X1 _3541_ (.A(net283),
    .Z(debug_transfer_count[104]));
 BUF_X1 _3542_ (.A(net284),
    .Z(debug_transfer_count[105]));
 BUF_X1 _3543_ (.A(net285),
    .Z(debug_transfer_count[106]));
 BUF_X1 _3544_ (.A(net286),
    .Z(debug_transfer_count[107]));
 BUF_X1 _3545_ (.A(net287),
    .Z(debug_transfer_count[108]));
 BUF_X1 _3546_ (.A(net288),
    .Z(debug_transfer_count[109]));
 BUF_X1 _3547_ (.A(net289),
    .Z(debug_transfer_count[110]));
 BUF_X1 _3548_ (.A(net290),
    .Z(debug_transfer_count[111]));
 BUF_X1 _3549_ (.A(net291),
    .Z(debug_transfer_count[112]));
 BUF_X1 _3550_ (.A(net292),
    .Z(debug_transfer_count[113]));
 BUF_X1 _3551_ (.A(net293),
    .Z(debug_transfer_count[114]));
 BUF_X1 _3552_ (.A(net294),
    .Z(debug_transfer_count[115]));
 BUF_X1 _3553_ (.A(net295),
    .Z(debug_transfer_count[116]));
 BUF_X1 _3554_ (.A(net296),
    .Z(debug_transfer_count[117]));
 BUF_X1 _3555_ (.A(net297),
    .Z(debug_transfer_count[118]));
 BUF_X1 _3556_ (.A(net298),
    .Z(debug_transfer_count[119]));
 BUF_X1 _3557_ (.A(net299),
    .Z(debug_transfer_count[120]));
 BUF_X1 _3558_ (.A(net300),
    .Z(debug_transfer_count[121]));
 BUF_X1 _3559_ (.A(net301),
    .Z(debug_transfer_count[122]));
 BUF_X1 _3560_ (.A(net302),
    .Z(debug_transfer_count[123]));
 BUF_X1 _3561_ (.A(net303),
    .Z(debug_transfer_count[124]));
 BUF_X1 _3562_ (.A(net304),
    .Z(debug_transfer_count[125]));
 BUF_X1 _3563_ (.A(net305),
    .Z(debug_transfer_count[126]));
 BUF_X1 _3564_ (.A(net306),
    .Z(debug_transfer_count[127]));
 BUF_X1 _3565_ (.A(net307),
    .Z(dst_addr[0]));
 BUF_X1 _3566_ (.A(net308),
    .Z(dst_addr[1]));
 BUF_X1 _3567_ (.A(net309),
    .Z(dst_addr[2]));
 BUF_X1 _3568_ (.A(net310),
    .Z(dst_addr[3]));
 BUF_X1 _3569_ (.A(net311),
    .Z(dst_addr[4]));
 BUF_X1 _3570_ (.A(net312),
    .Z(dst_addr[5]));
 BUF_X1 _3571_ (.A(net313),
    .Z(dst_addr[6]));
 BUF_X1 _3572_ (.A(net314),
    .Z(dst_addr[7]));
 BUF_X1 _3573_ (.A(net315),
    .Z(dst_addr[8]));
 BUF_X1 _3574_ (.A(net316),
    .Z(dst_addr[9]));
 BUF_X1 _3575_ (.A(net317),
    .Z(dst_addr[10]));
 BUF_X1 _3576_ (.A(net318),
    .Z(dst_addr[11]));
 BUF_X1 _3577_ (.A(net319),
    .Z(dst_addr[12]));
 BUF_X1 _3578_ (.A(net320),
    .Z(dst_addr[13]));
 BUF_X1 _3579_ (.A(net321),
    .Z(dst_addr[14]));
 BUF_X1 _3580_ (.A(net322),
    .Z(dst_addr[15]));
 BUF_X1 _3581_ (.A(net323),
    .Z(dst_addr[16]));
 BUF_X1 _3582_ (.A(net324),
    .Z(dst_addr[17]));
 BUF_X1 _3583_ (.A(net325),
    .Z(dst_addr[18]));
 BUF_X1 _3584_ (.A(net326),
    .Z(dst_addr[19]));
 BUF_X1 _3585_ (.A(net327),
    .Z(dst_addr[20]));
 BUF_X1 _3586_ (.A(net328),
    .Z(dst_addr[21]));
 BUF_X1 _3587_ (.A(net329),
    .Z(dst_addr[22]));
 BUF_X1 _3588_ (.A(net330),
    .Z(dst_addr[23]));
 BUF_X1 _3589_ (.A(net331),
    .Z(dst_addr[24]));
 BUF_X1 _3590_ (.A(net332),
    .Z(dst_addr[25]));
 BUF_X1 _3591_ (.A(net333),
    .Z(dst_addr[26]));
 BUF_X1 _3592_ (.A(net334),
    .Z(dst_addr[27]));
 BUF_X1 _3593_ (.A(net335),
    .Z(dst_addr[28]));
 BUF_X1 _3594_ (.A(net336),
    .Z(dst_addr[29]));
 BUF_X1 _3595_ (.A(net337),
    .Z(dst_addr[30]));
 BUF_X1 _3596_ (.A(net338),
    .Z(dst_addr[31]));
 BUF_X1 _3597_ (.A(net339),
    .Z(dst_addr[32]));
 BUF_X1 _3598_ (.A(net340),
    .Z(dst_addr[33]));
 BUF_X1 _3599_ (.A(net341),
    .Z(dst_addr[34]));
 BUF_X1 _3600_ (.A(net342),
    .Z(dst_addr[35]));
 BUF_X1 _3601_ (.A(net343),
    .Z(dst_addr[36]));
 BUF_X1 _3602_ (.A(net344),
    .Z(dst_addr[37]));
 BUF_X1 _3603_ (.A(net345),
    .Z(dst_addr[38]));
 BUF_X1 _3604_ (.A(net346),
    .Z(dst_addr[39]));
 BUF_X1 _3605_ (.A(net347),
    .Z(dst_addr[40]));
 BUF_X1 _3606_ (.A(net348),
    .Z(dst_addr[41]));
 BUF_X1 _3607_ (.A(net349),
    .Z(dst_addr[42]));
 BUF_X1 _3608_ (.A(net350),
    .Z(dst_addr[43]));
 BUF_X1 _3609_ (.A(net351),
    .Z(dst_addr[44]));
 BUF_X1 _3610_ (.A(net352),
    .Z(dst_addr[45]));
 BUF_X1 _3611_ (.A(net353),
    .Z(dst_addr[46]));
 BUF_X1 _3612_ (.A(net354),
    .Z(dst_addr[47]));
 BUF_X1 _3613_ (.A(net355),
    .Z(dst_addr[48]));
 BUF_X1 _3614_ (.A(net356),
    .Z(dst_addr[49]));
 BUF_X1 _3615_ (.A(net357),
    .Z(dst_addr[50]));
 BUF_X1 _3616_ (.A(net358),
    .Z(dst_addr[51]));
 BUF_X1 _3617_ (.A(net359),
    .Z(dst_addr[52]));
 BUF_X1 _3618_ (.A(net360),
    .Z(dst_addr[53]));
 BUF_X1 _3619_ (.A(net361),
    .Z(dst_addr[54]));
 BUF_X1 _3620_ (.A(net362),
    .Z(dst_addr[55]));
 BUF_X1 _3621_ (.A(net363),
    .Z(dst_addr[56]));
 BUF_X1 _3622_ (.A(net364),
    .Z(dst_addr[57]));
 BUF_X1 _3623_ (.A(net365),
    .Z(dst_addr[58]));
 BUF_X1 _3624_ (.A(net366),
    .Z(dst_addr[59]));
 BUF_X1 _3625_ (.A(net367),
    .Z(dst_addr[60]));
 BUF_X1 _3626_ (.A(net368),
    .Z(dst_addr[61]));
 BUF_X1 _3627_ (.A(net369),
    .Z(dst_addr[62]));
 BUF_X1 _3628_ (.A(net370),
    .Z(dst_addr[63]));
 BUF_X1 _3629_ (.A(net371),
    .Z(dst_addr[64]));
 BUF_X1 _3630_ (.A(net372),
    .Z(dst_addr[65]));
 BUF_X1 _3631_ (.A(net373),
    .Z(dst_addr[66]));
 BUF_X1 _3632_ (.A(net374),
    .Z(dst_addr[67]));
 BUF_X1 _3633_ (.A(net375),
    .Z(dst_addr[68]));
 BUF_X1 _3634_ (.A(net376),
    .Z(dst_addr[69]));
 BUF_X1 _3635_ (.A(net377),
    .Z(dst_addr[70]));
 BUF_X1 _3636_ (.A(net378),
    .Z(dst_addr[71]));
 BUF_X1 _3637_ (.A(net379),
    .Z(dst_addr[72]));
 BUF_X1 _3638_ (.A(net380),
    .Z(dst_addr[73]));
 BUF_X1 _3639_ (.A(net381),
    .Z(dst_addr[74]));
 BUF_X1 _3640_ (.A(net382),
    .Z(dst_addr[75]));
 BUF_X1 _3641_ (.A(net383),
    .Z(dst_addr[76]));
 BUF_X1 _3642_ (.A(net384),
    .Z(dst_addr[77]));
 BUF_X1 _3643_ (.A(net385),
    .Z(dst_addr[78]));
 BUF_X1 _3644_ (.A(net386),
    .Z(dst_addr[79]));
 BUF_X1 _3645_ (.A(net387),
    .Z(dst_addr[80]));
 BUF_X1 _3646_ (.A(net388),
    .Z(dst_addr[81]));
 BUF_X1 _3647_ (.A(net389),
    .Z(dst_addr[82]));
 BUF_X1 _3648_ (.A(net390),
    .Z(dst_addr[83]));
 BUF_X1 _3649_ (.A(net391),
    .Z(dst_addr[84]));
 BUF_X1 _3650_ (.A(net392),
    .Z(dst_addr[85]));
 BUF_X1 _3651_ (.A(net393),
    .Z(dst_addr[86]));
 BUF_X1 _3652_ (.A(net394),
    .Z(dst_addr[87]));
 BUF_X1 _3653_ (.A(net395),
    .Z(dst_addr[88]));
 BUF_X1 _3654_ (.A(net396),
    .Z(dst_addr[89]));
 BUF_X1 _3655_ (.A(net397),
    .Z(dst_addr[90]));
 BUF_X1 _3656_ (.A(net398),
    .Z(dst_addr[91]));
 BUF_X1 _3657_ (.A(net399),
    .Z(dst_addr[92]));
 BUF_X1 _3658_ (.A(net400),
    .Z(dst_addr[93]));
 BUF_X1 _3659_ (.A(net401),
    .Z(dst_addr[94]));
 BUF_X1 _3660_ (.A(net402),
    .Z(dst_addr[95]));
 BUF_X1 _3661_ (.A(net403),
    .Z(dst_addr[96]));
 BUF_X1 _3662_ (.A(net404),
    .Z(dst_addr[97]));
 BUF_X1 _3663_ (.A(net405),
    .Z(dst_addr[98]));
 BUF_X1 _3664_ (.A(net406),
    .Z(dst_addr[99]));
 BUF_X1 _3665_ (.A(net407),
    .Z(dst_addr[100]));
 BUF_X1 _3666_ (.A(net408),
    .Z(dst_addr[101]));
 BUF_X1 _3667_ (.A(net409),
    .Z(dst_addr[102]));
 BUF_X1 _3668_ (.A(net410),
    .Z(dst_addr[103]));
 BUF_X1 _3669_ (.A(net411),
    .Z(dst_addr[104]));
 BUF_X1 _3670_ (.A(net412),
    .Z(dst_addr[105]));
 BUF_X1 _3671_ (.A(net413),
    .Z(dst_addr[106]));
 BUF_X1 _3672_ (.A(net414),
    .Z(dst_addr[107]));
 BUF_X1 _3673_ (.A(net415),
    .Z(dst_addr[108]));
 BUF_X1 _3674_ (.A(net416),
    .Z(dst_addr[109]));
 BUF_X1 _3675_ (.A(net417),
    .Z(dst_addr[110]));
 BUF_X1 _3676_ (.A(net418),
    .Z(dst_addr[111]));
 BUF_X1 _3677_ (.A(net419),
    .Z(dst_addr[112]));
 BUF_X1 _3678_ (.A(net420),
    .Z(dst_addr[113]));
 BUF_X1 _3679_ (.A(net421),
    .Z(dst_addr[114]));
 BUF_X1 _3680_ (.A(net422),
    .Z(dst_addr[115]));
 BUF_X1 _3681_ (.A(net423),
    .Z(dst_addr[116]));
 BUF_X1 _3682_ (.A(net424),
    .Z(dst_addr[117]));
 BUF_X1 _3683_ (.A(net425),
    .Z(dst_addr[118]));
 BUF_X1 _3684_ (.A(net426),
    .Z(dst_addr[119]));
 BUF_X1 _3685_ (.A(net427),
    .Z(dst_addr[120]));
 BUF_X1 _3686_ (.A(net428),
    .Z(dst_addr[121]));
 BUF_X1 _3687_ (.A(net429),
    .Z(dst_addr[122]));
 BUF_X1 _3688_ (.A(net430),
    .Z(dst_addr[123]));
 BUF_X1 _3689_ (.A(net431),
    .Z(dst_addr[124]));
 BUF_X1 _3690_ (.A(net432),
    .Z(dst_addr[125]));
 BUF_X1 _3691_ (.A(net433),
    .Z(dst_addr[126]));
 BUF_X1 _3692_ (.A(net434),
    .Z(dst_addr[127]));
 BUF_X1 _3693_ (.A(net435),
    .Z(dst_wdata[0]));
 BUF_X1 _3694_ (.A(net436),
    .Z(dst_wdata[1]));
 BUF_X1 _3695_ (.A(net437),
    .Z(dst_wdata[2]));
 BUF_X1 _3696_ (.A(net438),
    .Z(dst_wdata[3]));
 BUF_X1 _3697_ (.A(net439),
    .Z(dst_wdata[4]));
 BUF_X1 _3698_ (.A(net440),
    .Z(dst_wdata[5]));
 BUF_X1 _3699_ (.A(net441),
    .Z(dst_wdata[6]));
 BUF_X1 _3700_ (.A(net442),
    .Z(dst_wdata[7]));
 BUF_X1 _3701_ (.A(net443),
    .Z(dst_wdata[8]));
 BUF_X1 _3702_ (.A(net444),
    .Z(dst_wdata[9]));
 BUF_X1 _3703_ (.A(net445),
    .Z(dst_wdata[10]));
 BUF_X1 _3704_ (.A(net446),
    .Z(dst_wdata[11]));
 BUF_X1 _3705_ (.A(net447),
    .Z(dst_wdata[12]));
 BUF_X1 _3706_ (.A(net448),
    .Z(dst_wdata[13]));
 BUF_X1 _3707_ (.A(net449),
    .Z(dst_wdata[14]));
 BUF_X1 _3708_ (.A(net450),
    .Z(dst_wdata[15]));
 BUF_X1 _3709_ (.A(net451),
    .Z(dst_wdata[16]));
 BUF_X1 _3710_ (.A(net452),
    .Z(dst_wdata[17]));
 BUF_X1 _3711_ (.A(net453),
    .Z(dst_wdata[18]));
 BUF_X1 _3712_ (.A(net454),
    .Z(dst_wdata[19]));
 BUF_X1 _3713_ (.A(net455),
    .Z(dst_wdata[20]));
 BUF_X1 _3714_ (.A(net456),
    .Z(dst_wdata[21]));
 BUF_X1 _3715_ (.A(net457),
    .Z(dst_wdata[22]));
 BUF_X1 _3716_ (.A(net458),
    .Z(dst_wdata[23]));
 BUF_X1 _3717_ (.A(net459),
    .Z(dst_wdata[24]));
 BUF_X1 _3718_ (.A(net460),
    .Z(dst_wdata[25]));
 BUF_X1 _3719_ (.A(net461),
    .Z(dst_wdata[26]));
 BUF_X1 _3720_ (.A(net462),
    .Z(dst_wdata[27]));
 BUF_X1 _3721_ (.A(net463),
    .Z(dst_wdata[28]));
 BUF_X1 _3722_ (.A(net464),
    .Z(dst_wdata[29]));
 BUF_X1 _3723_ (.A(net465),
    .Z(dst_wdata[30]));
 BUF_X1 _3724_ (.A(net466),
    .Z(dst_wdata[31]));
 BUF_X1 _3725_ (.A(net467),
    .Z(dst_wdata[32]));
 BUF_X1 _3726_ (.A(net468),
    .Z(dst_wdata[33]));
 BUF_X1 _3727_ (.A(net469),
    .Z(dst_wdata[34]));
 BUF_X1 _3728_ (.A(net470),
    .Z(dst_wdata[35]));
 BUF_X1 _3729_ (.A(net471),
    .Z(dst_wdata[36]));
 BUF_X1 _3730_ (.A(net472),
    .Z(dst_wdata[37]));
 BUF_X1 _3731_ (.A(net473),
    .Z(dst_wdata[38]));
 BUF_X1 _3732_ (.A(net474),
    .Z(dst_wdata[39]));
 BUF_X1 _3733_ (.A(net475),
    .Z(dst_wdata[40]));
 BUF_X1 _3734_ (.A(net476),
    .Z(dst_wdata[41]));
 BUF_X1 _3735_ (.A(net477),
    .Z(dst_wdata[42]));
 BUF_X1 _3736_ (.A(net478),
    .Z(dst_wdata[43]));
 BUF_X1 _3737_ (.A(net479),
    .Z(dst_wdata[44]));
 BUF_X1 _3738_ (.A(net480),
    .Z(dst_wdata[45]));
 BUF_X1 _3739_ (.A(net481),
    .Z(dst_wdata[46]));
 BUF_X1 _3740_ (.A(net482),
    .Z(dst_wdata[47]));
 BUF_X1 _3741_ (.A(net483),
    .Z(dst_wdata[48]));
 BUF_X1 _3742_ (.A(net484),
    .Z(dst_wdata[49]));
 BUF_X1 _3743_ (.A(net485),
    .Z(dst_wdata[50]));
 BUF_X1 _3744_ (.A(net486),
    .Z(dst_wdata[51]));
 BUF_X1 _3745_ (.A(net487),
    .Z(dst_wdata[52]));
 BUF_X1 _3746_ (.A(net488),
    .Z(dst_wdata[53]));
 BUF_X1 _3747_ (.A(net489),
    .Z(dst_wdata[54]));
 BUF_X1 _3748_ (.A(net490),
    .Z(dst_wdata[55]));
 BUF_X1 _3749_ (.A(net491),
    .Z(dst_wdata[56]));
 BUF_X1 _3750_ (.A(net492),
    .Z(dst_wdata[57]));
 BUF_X1 _3751_ (.A(net493),
    .Z(dst_wdata[58]));
 BUF_X1 _3752_ (.A(net494),
    .Z(dst_wdata[59]));
 BUF_X1 _3753_ (.A(net495),
    .Z(dst_wdata[60]));
 BUF_X1 _3754_ (.A(net496),
    .Z(dst_wdata[61]));
 BUF_X1 _3755_ (.A(net497),
    .Z(dst_wdata[62]));
 BUF_X1 _3756_ (.A(net498),
    .Z(dst_wdata[63]));
 BUF_X1 _3757_ (.A(net499),
    .Z(dst_wdata[64]));
 BUF_X1 _3758_ (.A(net500),
    .Z(dst_wdata[65]));
 BUF_X1 _3759_ (.A(net501),
    .Z(dst_wdata[66]));
 BUF_X1 _3760_ (.A(net502),
    .Z(dst_wdata[67]));
 BUF_X1 _3761_ (.A(net503),
    .Z(dst_wdata[68]));
 BUF_X1 _3762_ (.A(net504),
    .Z(dst_wdata[69]));
 BUF_X1 _3763_ (.A(net505),
    .Z(dst_wdata[70]));
 BUF_X1 _3764_ (.A(net506),
    .Z(dst_wdata[71]));
 BUF_X1 _3765_ (.A(net507),
    .Z(dst_wdata[72]));
 BUF_X1 _3766_ (.A(net508),
    .Z(dst_wdata[73]));
 BUF_X1 _3767_ (.A(net509),
    .Z(dst_wdata[74]));
 BUF_X1 _3768_ (.A(net510),
    .Z(dst_wdata[75]));
 BUF_X1 _3769_ (.A(net511),
    .Z(dst_wdata[76]));
 BUF_X1 _3770_ (.A(net512),
    .Z(dst_wdata[77]));
 BUF_X1 _3771_ (.A(net513),
    .Z(dst_wdata[78]));
 BUF_X1 _3772_ (.A(net514),
    .Z(dst_wdata[79]));
 BUF_X1 _3773_ (.A(net515),
    .Z(dst_wdata[80]));
 BUF_X1 _3774_ (.A(net516),
    .Z(dst_wdata[81]));
 BUF_X1 _3775_ (.A(net517),
    .Z(dst_wdata[82]));
 BUF_X1 _3776_ (.A(net518),
    .Z(dst_wdata[83]));
 BUF_X1 _3777_ (.A(net519),
    .Z(dst_wdata[84]));
 BUF_X1 _3778_ (.A(net520),
    .Z(dst_wdata[85]));
 BUF_X1 _3779_ (.A(net521),
    .Z(dst_wdata[86]));
 BUF_X1 _3780_ (.A(net522),
    .Z(dst_wdata[87]));
 BUF_X1 _3781_ (.A(net523),
    .Z(dst_wdata[88]));
 BUF_X1 _3782_ (.A(net524),
    .Z(dst_wdata[89]));
 BUF_X1 _3783_ (.A(net525),
    .Z(dst_wdata[90]));
 BUF_X1 _3784_ (.A(net526),
    .Z(dst_wdata[91]));
 BUF_X1 _3785_ (.A(net527),
    .Z(dst_wdata[92]));
 BUF_X1 _3786_ (.A(net528),
    .Z(dst_wdata[93]));
 BUF_X1 _3787_ (.A(net529),
    .Z(dst_wdata[94]));
 BUF_X1 _3788_ (.A(net530),
    .Z(dst_wdata[95]));
 BUF_X1 _3789_ (.A(net531),
    .Z(dst_wdata[96]));
 BUF_X1 _3790_ (.A(net532),
    .Z(dst_wdata[97]));
 BUF_X1 _3791_ (.A(net533),
    .Z(dst_wdata[98]));
 BUF_X1 _3792_ (.A(net534),
    .Z(dst_wdata[99]));
 BUF_X1 _3793_ (.A(net535),
    .Z(dst_wdata[100]));
 BUF_X1 _3794_ (.A(net536),
    .Z(dst_wdata[101]));
 BUF_X1 _3795_ (.A(net537),
    .Z(dst_wdata[102]));
 BUF_X1 _3796_ (.A(net538),
    .Z(dst_wdata[103]));
 BUF_X1 _3797_ (.A(net539),
    .Z(dst_wdata[104]));
 BUF_X1 _3798_ (.A(net540),
    .Z(dst_wdata[105]));
 BUF_X1 _3799_ (.A(net541),
    .Z(dst_wdata[106]));
 BUF_X1 _3800_ (.A(net542),
    .Z(dst_wdata[107]));
 BUF_X1 _3801_ (.A(net543),
    .Z(dst_wdata[108]));
 BUF_X1 _3802_ (.A(net544),
    .Z(dst_wdata[109]));
 BUF_X1 _3803_ (.A(net545),
    .Z(dst_wdata[110]));
 BUF_X1 _3804_ (.A(net546),
    .Z(dst_wdata[111]));
 BUF_X1 _3805_ (.A(net547),
    .Z(dst_wdata[112]));
 BUF_X1 _3806_ (.A(net548),
    .Z(dst_wdata[113]));
 BUF_X1 _3807_ (.A(net549),
    .Z(dst_wdata[114]));
 BUF_X1 _3808_ (.A(net550),
    .Z(dst_wdata[115]));
 BUF_X1 _3809_ (.A(net551),
    .Z(dst_wdata[116]));
 BUF_X1 _3810_ (.A(net552),
    .Z(dst_wdata[117]));
 BUF_X1 _3811_ (.A(net553),
    .Z(dst_wdata[118]));
 BUF_X1 _3812_ (.A(net554),
    .Z(dst_wdata[119]));
 BUF_X1 _3813_ (.A(net555),
    .Z(dst_wdata[120]));
 BUF_X1 _3814_ (.A(net556),
    .Z(dst_wdata[121]));
 BUF_X1 _3815_ (.A(net557),
    .Z(dst_wdata[122]));
 BUF_X1 _3816_ (.A(net558),
    .Z(dst_wdata[123]));
 BUF_X1 _3817_ (.A(net559),
    .Z(dst_wdata[124]));
 BUF_X1 _3818_ (.A(net560),
    .Z(dst_wdata[125]));
 BUF_X1 _3819_ (.A(net561),
    .Z(dst_wdata[126]));
 BUF_X1 _3820_ (.A(net562),
    .Z(dst_wdata[127]));
 BUF_X1 _3821_ (.A(net563),
    .Z(dst_wstrb[0]));
 BUF_X1 _3822_ (.A(net564),
    .Z(dst_wstrb[1]));
 BUF_X1 _3823_ (.A(net565),
    .Z(dst_wstrb[2]));
 BUF_X1 _3824_ (.A(net566),
    .Z(dst_wstrb[3]));
 BUF_X1 _3825_ (.A(net567),
    .Z(dst_wstrb[4]));
 BUF_X1 _3826_ (.A(net568),
    .Z(dst_wstrb[5]));
 BUF_X1 _3827_ (.A(net569),
    .Z(dst_wstrb[6]));
 BUF_X1 _3828_ (.A(net570),
    .Z(dst_wstrb[7]));
 BUF_X1 _3829_ (.A(net571),
    .Z(dst_wstrb[8]));
 BUF_X1 _3830_ (.A(net572),
    .Z(dst_wstrb[9]));
 BUF_X1 _3831_ (.A(net573),
    .Z(dst_wstrb[10]));
 BUF_X1 _3832_ (.A(net574),
    .Z(dst_wstrb[11]));
 BUF_X1 _3833_ (.A(net575),
    .Z(dst_wstrb[12]));
 BUF_X1 _3834_ (.A(net576),
    .Z(dst_wstrb[13]));
 BUF_X1 _3835_ (.A(net577),
    .Z(dst_wstrb[14]));
 BUF_X1 _3836_ (.A(net578),
    .Z(dst_wstrb[15]));
 BUF_X1 _3837_ (.A(net579),
    .Z(src_addr[0]));
 BUF_X1 _3838_ (.A(net580),
    .Z(src_addr[1]));
 BUF_X1 _3839_ (.A(net581),
    .Z(src_addr[2]));
 BUF_X1 _3840_ (.A(net582),
    .Z(src_addr[3]));
 BUF_X1 _3841_ (.A(net583),
    .Z(src_addr[4]));
 BUF_X1 _3842_ (.A(net584),
    .Z(src_addr[5]));
 BUF_X1 _3843_ (.A(net585),
    .Z(src_addr[6]));
 BUF_X1 _3844_ (.A(net586),
    .Z(src_addr[7]));
 BUF_X1 _3845_ (.A(net587),
    .Z(src_addr[8]));
 BUF_X1 _3846_ (.A(net588),
    .Z(src_addr[9]));
 BUF_X1 _3847_ (.A(net589),
    .Z(src_addr[10]));
 BUF_X1 _3848_ (.A(net590),
    .Z(src_addr[11]));
 BUF_X1 _3849_ (.A(net591),
    .Z(src_addr[12]));
 BUF_X1 _3850_ (.A(net592),
    .Z(src_addr[13]));
 BUF_X1 _3851_ (.A(net593),
    .Z(src_addr[14]));
 BUF_X1 _3852_ (.A(net594),
    .Z(src_addr[15]));
 BUF_X1 _3853_ (.A(net595),
    .Z(src_addr[16]));
 BUF_X1 _3854_ (.A(net596),
    .Z(src_addr[17]));
 BUF_X1 _3855_ (.A(net597),
    .Z(src_addr[18]));
 BUF_X1 _3856_ (.A(net598),
    .Z(src_addr[19]));
 BUF_X1 _3857_ (.A(net599),
    .Z(src_addr[20]));
 BUF_X1 _3858_ (.A(net600),
    .Z(src_addr[21]));
 BUF_X1 _3859_ (.A(net601),
    .Z(src_addr[22]));
 BUF_X1 _3860_ (.A(net602),
    .Z(src_addr[23]));
 BUF_X1 _3861_ (.A(net603),
    .Z(src_addr[24]));
 BUF_X1 _3862_ (.A(net604),
    .Z(src_addr[25]));
 BUF_X1 _3863_ (.A(net605),
    .Z(src_addr[26]));
 BUF_X1 _3864_ (.A(net606),
    .Z(src_addr[27]));
 BUF_X1 _3865_ (.A(net607),
    .Z(src_addr[28]));
 BUF_X1 _3866_ (.A(net608),
    .Z(src_addr[29]));
 BUF_X1 _3867_ (.A(net609),
    .Z(src_addr[30]));
 BUF_X1 _3868_ (.A(net610),
    .Z(src_addr[31]));
 BUF_X1 _3869_ (.A(net611),
    .Z(src_addr[32]));
 BUF_X1 _3870_ (.A(net612),
    .Z(src_addr[33]));
 BUF_X1 _3871_ (.A(net613),
    .Z(src_addr[34]));
 BUF_X1 _3872_ (.A(net614),
    .Z(src_addr[35]));
 BUF_X1 _3873_ (.A(net615),
    .Z(src_addr[36]));
 BUF_X1 _3874_ (.A(net616),
    .Z(src_addr[37]));
 BUF_X1 _3875_ (.A(net617),
    .Z(src_addr[38]));
 BUF_X1 _3876_ (.A(net618),
    .Z(src_addr[39]));
 BUF_X1 _3877_ (.A(net619),
    .Z(src_addr[40]));
 BUF_X1 _3878_ (.A(net620),
    .Z(src_addr[41]));
 BUF_X1 _3879_ (.A(net621),
    .Z(src_addr[42]));
 BUF_X1 _3880_ (.A(net622),
    .Z(src_addr[43]));
 BUF_X1 _3881_ (.A(net623),
    .Z(src_addr[44]));
 BUF_X1 _3882_ (.A(net624),
    .Z(src_addr[45]));
 BUF_X1 _3883_ (.A(net625),
    .Z(src_addr[46]));
 BUF_X1 _3884_ (.A(net626),
    .Z(src_addr[47]));
 BUF_X1 _3885_ (.A(net627),
    .Z(src_addr[48]));
 BUF_X1 _3886_ (.A(net628),
    .Z(src_addr[49]));
 BUF_X1 _3887_ (.A(net629),
    .Z(src_addr[50]));
 BUF_X1 _3888_ (.A(net630),
    .Z(src_addr[51]));
 BUF_X1 _3889_ (.A(net631),
    .Z(src_addr[52]));
 BUF_X1 _3890_ (.A(net632),
    .Z(src_addr[53]));
 BUF_X1 _3891_ (.A(net633),
    .Z(src_addr[54]));
 BUF_X1 _3892_ (.A(net634),
    .Z(src_addr[55]));
 BUF_X1 _3893_ (.A(net635),
    .Z(src_addr[56]));
 BUF_X1 _3894_ (.A(net636),
    .Z(src_addr[57]));
 BUF_X1 _3895_ (.A(net637),
    .Z(src_addr[58]));
 BUF_X1 _3896_ (.A(net638),
    .Z(src_addr[59]));
 BUF_X1 _3897_ (.A(net639),
    .Z(src_addr[60]));
 BUF_X1 _3898_ (.A(net640),
    .Z(src_addr[61]));
 BUF_X1 _3899_ (.A(net641),
    .Z(src_addr[62]));
 BUF_X1 _3900_ (.A(net642),
    .Z(src_addr[63]));
 BUF_X1 _3901_ (.A(net643),
    .Z(src_addr[64]));
 BUF_X1 _3902_ (.A(net644),
    .Z(src_addr[65]));
 BUF_X1 _3903_ (.A(net645),
    .Z(src_addr[66]));
 BUF_X1 _3904_ (.A(net646),
    .Z(src_addr[67]));
 BUF_X1 _3905_ (.A(net647),
    .Z(src_addr[68]));
 BUF_X1 _3906_ (.A(net648),
    .Z(src_addr[69]));
 BUF_X1 _3907_ (.A(net649),
    .Z(src_addr[70]));
 BUF_X1 _3908_ (.A(net650),
    .Z(src_addr[71]));
 BUF_X1 _3909_ (.A(net651),
    .Z(src_addr[72]));
 BUF_X1 _3910_ (.A(net652),
    .Z(src_addr[73]));
 BUF_X1 _3911_ (.A(net653),
    .Z(src_addr[74]));
 BUF_X1 _3912_ (.A(net654),
    .Z(src_addr[75]));
 BUF_X1 _3913_ (.A(net655),
    .Z(src_addr[76]));
 BUF_X1 _3914_ (.A(net656),
    .Z(src_addr[77]));
 BUF_X1 _3915_ (.A(net657),
    .Z(src_addr[78]));
 BUF_X1 _3916_ (.A(net658),
    .Z(src_addr[79]));
 BUF_X1 _3917_ (.A(net659),
    .Z(src_addr[80]));
 BUF_X1 _3918_ (.A(net660),
    .Z(src_addr[81]));
 BUF_X1 _3919_ (.A(net661),
    .Z(src_addr[82]));
 BUF_X1 _3920_ (.A(net662),
    .Z(src_addr[83]));
 BUF_X1 _3921_ (.A(net663),
    .Z(src_addr[84]));
 BUF_X1 _3922_ (.A(net664),
    .Z(src_addr[85]));
 BUF_X1 _3923_ (.A(net665),
    .Z(src_addr[86]));
 BUF_X1 _3924_ (.A(net666),
    .Z(src_addr[87]));
 BUF_X1 _3925_ (.A(net667),
    .Z(src_addr[88]));
 BUF_X1 _3926_ (.A(net668),
    .Z(src_addr[89]));
 BUF_X1 _3927_ (.A(net669),
    .Z(src_addr[90]));
 BUF_X1 _3928_ (.A(net670),
    .Z(src_addr[91]));
 BUF_X1 _3929_ (.A(net671),
    .Z(src_addr[92]));
 BUF_X1 _3930_ (.A(net672),
    .Z(src_addr[93]));
 BUF_X1 _3931_ (.A(net673),
    .Z(src_addr[94]));
 BUF_X1 _3932_ (.A(net674),
    .Z(src_addr[95]));
 BUF_X1 _3933_ (.A(net675),
    .Z(src_addr[96]));
 BUF_X1 _3934_ (.A(net676),
    .Z(src_addr[97]));
 BUF_X1 _3935_ (.A(net677),
    .Z(src_addr[98]));
 BUF_X1 _3936_ (.A(net678),
    .Z(src_addr[99]));
 BUF_X1 _3937_ (.A(net679),
    .Z(src_addr[100]));
 BUF_X1 _3938_ (.A(net680),
    .Z(src_addr[101]));
 BUF_X1 _3939_ (.A(net681),
    .Z(src_addr[102]));
 BUF_X1 _3940_ (.A(net682),
    .Z(src_addr[103]));
 BUF_X1 _3941_ (.A(net683),
    .Z(src_addr[104]));
 BUF_X1 _3942_ (.A(net684),
    .Z(src_addr[105]));
 BUF_X1 _3943_ (.A(net685),
    .Z(src_addr[106]));
 BUF_X1 _3944_ (.A(net686),
    .Z(src_addr[107]));
 BUF_X1 _3945_ (.A(net687),
    .Z(src_addr[108]));
 BUF_X1 _3946_ (.A(net688),
    .Z(src_addr[109]));
 BUF_X1 _3947_ (.A(net689),
    .Z(src_addr[110]));
 BUF_X1 _3948_ (.A(net690),
    .Z(src_addr[111]));
 BUF_X1 _3949_ (.A(net691),
    .Z(src_addr[112]));
 BUF_X1 _3950_ (.A(net692),
    .Z(src_addr[113]));
 BUF_X1 _3951_ (.A(net693),
    .Z(src_addr[114]));
 BUF_X1 _3952_ (.A(net694),
    .Z(src_addr[115]));
 BUF_X1 _3953_ (.A(net695),
    .Z(src_addr[116]));
 BUF_X1 _3954_ (.A(net696),
    .Z(src_addr[117]));
 BUF_X1 _3955_ (.A(net697),
    .Z(src_addr[118]));
 BUF_X1 _3956_ (.A(net698),
    .Z(src_addr[119]));
 BUF_X1 _3957_ (.A(net699),
    .Z(src_addr[120]));
 BUF_X1 _3958_ (.A(net700),
    .Z(src_addr[121]));
 BUF_X1 _3959_ (.A(net701),
    .Z(src_addr[122]));
 BUF_X1 _3960_ (.A(net702),
    .Z(src_addr[123]));
 BUF_X1 _3961_ (.A(net703),
    .Z(src_addr[124]));
 BUF_X1 _3962_ (.A(net704),
    .Z(src_addr[125]));
 BUF_X1 _3963_ (.A(net705),
    .Z(src_addr[126]));
 BUF_X1 _3964_ (.A(net706),
    .Z(src_addr[127]));
 DFF_X2 \active_channel_count[0]$_SDFF_PN0_  (.D(_0024_),
    .CK(clknet_4_6_0_clk),
    .Q(\active_channel_count[0] ),
    .QN(_1861_));
 DFF_X1 \active_channel_count[1]$_SDFF_PN0_  (.D(_0025_),
    .CK(clknet_4_7_0_clk),
    .Q(\active_channel_count[1] ),
    .QN(_1862_));
 DFF_X1 \active_channel_count[2]$_SDFF_PN0_  (.D(_0026_),
    .CK(clknet_4_7_0_clk),
    .Q(\active_channel_count[2] ),
    .QN(_1440_));
 DFF_X1 \active_channel_count[3]$_SDFF_PN0_  (.D(_0027_),
    .CK(clknet_4_7_0_clk),
    .Q(\active_channel_count[3] ),
    .QN(_1439_));
 DFF_X2 \channel_busy[0]$_SDFF_PN0_  (.D(_0028_),
    .CK(clknet_4_7_0_clk),
    .Q(net138),
    .QN(_1438_));
 DFF_X2 \channel_busy[1]$_SDFF_PN0_  (.D(_0029_),
    .CK(clknet_4_0_0_clk),
    .Q(net139),
    .QN(_1437_));
 DFF_X2 \channel_busy[2]$_SDFF_PN0_  (.D(_0030_),
    .CK(clknet_4_15_0_clk),
    .Q(net140),
    .QN(_1436_));
 DFF_X2 \channel_busy[3]$_SDFF_PN0_  (.D(_0031_),
    .CK(clknet_4_8_0_clk),
    .Q(net141),
    .QN(_1435_));
 DFF_X1 \channel_done[0]$_SDFF_PN0_  (.D(_0032_),
    .CK(clknet_4_7_0_clk),
    .Q(net142),
    .QN(_1434_));
 DFF_X1 \channel_done[1]$_SDFF_PN0_  (.D(_0033_),
    .CK(clknet_4_0_0_clk),
    .Q(net143),
    .QN(_1433_));
 DFF_X2 \channel_done[2]$_SDFF_PN0_  (.D(_0034_),
    .CK(clknet_4_9_0_clk),
    .Q(net144),
    .QN(_1432_));
 DFF_X2 \channel_done[3]$_SDFF_PN0_  (.D(_0035_),
    .CK(clknet_4_10_0_clk),
    .Q(net145),
    .QN(_1441_));
 DFF_X1 \channel_state[0][0]$_DFF_P_  (.D(_0004_),
    .CK(clknet_4_7_0_clk),
    .Q(\channel_state[0][0] ),
    .QN(_1442_));
 DFF_X1 \channel_state[0][1]$_DFF_P_  (.D(_0005_),
    .CK(clknet_4_7_0_clk),
    .Q(\channel_state[0][1] ),
    .QN(_1443_));
 DFF_X1 \channel_state[0][2]$_DFF_P_  (.D(_0006_),
    .CK(clknet_4_7_0_clk),
    .Q(\channel_state[0][2] ),
    .QN(_1444_));
 DFF_X1 \channel_state[0][3]$_DFF_P_  (.D(_0007_),
    .CK(clknet_4_7_0_clk),
    .Q(\channel_state[0][3] ),
    .QN(_1445_));
 DFF_X1 \channel_state[0][4]$_DFF_P_  (.D(_0008_),
    .CK(clknet_4_7_0_clk),
    .Q(\channel_state[0][4] ),
    .QN(_1446_));
 DFF_X1 \channel_state[0][5]$_DFF_P_  (.D(_0000_),
    .CK(clknet_4_7_0_clk),
    .Q(\channel_state[0][5] ),
    .QN(_1447_));
 DFF_X1 \channel_state[1][0]$_DFF_P_  (.D(_0009_),
    .CK(clknet_4_3_0_clk),
    .Q(\channel_state[1][0] ),
    .QN(_1448_));
 DFF_X2 \channel_state[1][1]$_DFF_P_  (.D(_0010_),
    .CK(clknet_4_2_0_clk),
    .Q(\channel_state[1][1] ),
    .QN(_1449_));
 DFF_X1 \channel_state[1][2]$_DFF_P_  (.D(_0011_),
    .CK(clknet_4_3_0_clk),
    .Q(\channel_state[1][2] ),
    .QN(_1450_));
 DFF_X1 \channel_state[1][3]$_DFF_P_  (.D(_0012_),
    .CK(clknet_4_0_0_clk),
    .Q(\channel_state[1][3] ),
    .QN(_1451_));
 DFF_X1 \channel_state[1][4]$_DFF_P_  (.D(_0013_),
    .CK(clknet_4_3_0_clk),
    .Q(\channel_state[1][4] ),
    .QN(_1452_));
 DFF_X1 \channel_state[1][5]$_DFF_P_  (.D(_0001_),
    .CK(clknet_4_3_0_clk),
    .Q(\channel_state[1][5] ),
    .QN(_1453_));
 DFF_X1 \channel_state[2][0]$_DFF_P_  (.D(_0014_),
    .CK(clknet_4_6_0_clk),
    .Q(\channel_state[2][0] ),
    .QN(_1454_));
 DFF_X1 \channel_state[2][1]$_DFF_P_  (.D(_0015_),
    .CK(clknet_4_9_0_clk),
    .Q(\channel_state[2][1] ),
    .QN(_1455_));
 DFF_X2 \channel_state[2][2]$_DFF_P_  (.D(_0016_),
    .CK(clknet_4_6_0_clk),
    .Q(\channel_state[2][2] ),
    .QN(_1456_));
 DFF_X2 \channel_state[2][3]$_DFF_P_  (.D(_0017_),
    .CK(clknet_4_15_0_clk),
    .Q(\channel_state[2][3] ),
    .QN(_1457_));
 DFF_X2 \channel_state[2][4]$_DFF_P_  (.D(_0018_),
    .CK(clknet_4_9_0_clk),
    .Q(\channel_state[2][4] ),
    .QN(_1458_));
 DFF_X1 \channel_state[2][5]$_DFF_P_  (.D(_0002_),
    .CK(clknet_4_6_0_clk),
    .Q(\channel_state[2][5] ),
    .QN(_1459_));
 DFF_X1 \channel_state[3][0]$_DFF_P_  (.D(_0019_),
    .CK(clknet_4_8_0_clk),
    .Q(\channel_state[3][0] ),
    .QN(_1460_));
 DFF_X1 \channel_state[3][1]$_DFF_P_  (.D(_0020_),
    .CK(clknet_4_8_0_clk),
    .Q(\channel_state[3][1] ),
    .QN(_1461_));
 DFF_X1 \channel_state[3][2]$_DFF_P_  (.D(_0021_),
    .CK(clknet_4_8_0_clk),
    .Q(\channel_state[3][2] ),
    .QN(_1462_));
 DFF_X1 \channel_state[3][3]$_DFF_P_  (.D(_0022_),
    .CK(clknet_4_8_0_clk),
    .Q(\channel_state[3][3] ),
    .QN(_1463_));
 DFF_X1 \channel_state[3][4]$_DFF_P_  (.D(_0023_),
    .CK(clknet_4_8_0_clk),
    .Q(\channel_state[3][4] ),
    .QN(_1464_));
 DFF_X1 \channel_state[3][5]$_DFF_P_  (.D(_0003_),
    .CK(clknet_4_8_0_clk),
    .Q(\channel_state[3][5] ),
    .QN(_1431_));
 DFF_X1 \debug_active_channels[0]$_SDFF_PN0_  (.D(_0036_),
    .CK(clknet_4_7_0_clk),
    .Q(net146),
    .QN(_1430_));
 DFF_X1 \debug_active_channels[1]$_SDFF_PN0_  (.D(_0037_),
    .CK(clknet_4_7_0_clk),
    .Q(net147),
    .QN(_1429_));
 DFF_X1 \debug_active_channels[2]$_SDFF_PN0_  (.D(_0038_),
    .CK(clknet_4_7_0_clk),
    .Q(net148),
    .QN(_1428_));
 DFF_X1 \debug_active_channels[3]$_SDFF_PN0_  (.D(_0039_),
    .CK(clknet_4_7_0_clk),
    .Q(net149),
    .QN(_1427_));
 DFF_X1 \debug_has_active_channels$_SDFF_PN0_  (.D(_0040_),
    .CK(clknet_4_7_0_clk),
    .Q(net150),
    .QN(_1426_));
 DFF_X1 \dst_write[0]$_SDFFE_PN0P_  (.D(_0041_),
    .CK(clknet_4_7_0_clk),
    .Q(net151),
    .QN(_1425_));
 DFF_X2 \dst_write[1]$_SDFFE_PN0P_  (.D(_0042_),
    .CK(clknet_4_3_0_clk),
    .Q(net152),
    .QN(_1424_));
 DFF_X1 \dst_write[2]$_SDFFE_PN0P_  (.D(_0043_),
    .CK(clknet_4_6_0_clk),
    .Q(net153),
    .QN(_1423_));
 DFF_X2 \dst_write[3]$_SDFFE_PN0P_  (.D(_0044_),
    .CK(clknet_4_9_0_clk),
    .Q(net154),
    .QN(_1422_));
 DFF_X1 \src_read[0]$_SDFF_PN0_  (.D(_0045_),
    .CK(clknet_4_7_0_clk),
    .Q(net155),
    .QN(_1421_));
 DFF_X1 \src_read[1]$_SDFF_PN0_  (.D(_0046_),
    .CK(clknet_4_2_0_clk),
    .Q(net156),
    .QN(_1420_));
 DFF_X1 \src_read[2]$_SDFF_PN0_  (.D(_0047_),
    .CK(clknet_4_6_0_clk),
    .Q(net157),
    .QN(_1419_));
 DFF_X1 \src_read[3]$_SDFF_PN0_  (.D(_0048_),
    .CK(clknet_4_7_0_clk),
    .Q(net158),
    .QN(_1418_));
 DFF_X1 \src_rready[0]$_SDFFE_PN0P_  (.D(_0049_),
    .CK(clknet_4_7_0_clk),
    .Q(net159),
    .QN(_1417_));
 DFF_X2 \src_rready[1]$_SDFFE_PN0P_  (.D(_0050_),
    .CK(clknet_4_3_0_clk),
    .Q(net160),
    .QN(_1416_));
 DFF_X1 \src_rready[2]$_SDFFE_PN0P_  (.D(_0051_),
    .CK(clknet_4_6_0_clk),
    .Q(net161),
    .QN(_1415_));
 DFF_X2 \src_rready[3]$_SDFFE_PN0P_  (.D(_0052_),
    .CK(clknet_4_8_0_clk),
    .Q(net162),
    .QN(_1414_));
 DFF_X2 \transfer_count[0][0]$_SDFF_PN0_  (.D(_0053_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][0] ),
    .QN(_1759_));
 DFF_X1 \transfer_count[0][10]$_SDFF_PN0_  (.D(_0054_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][10] ),
    .QN(_1413_));
 DFF_X1 \transfer_count[0][11]$_SDFF_PN0_  (.D(_0055_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][11] ),
    .QN(_1412_));
 DFF_X1 \transfer_count[0][12]$_SDFF_PN0_  (.D(_0056_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][12] ),
    .QN(_1411_));
 DFF_X1 \transfer_count[0][13]$_SDFF_PN0_  (.D(_0057_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][13] ),
    .QN(_1410_));
 DFF_X1 \transfer_count[0][14]$_SDFF_PN0_  (.D(_0058_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][14] ),
    .QN(_1409_));
 DFF_X1 \transfer_count[0][15]$_SDFF_PN0_  (.D(_0059_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][15] ),
    .QN(_1408_));
 DFF_X1 \transfer_count[0][16]$_SDFF_PN0_  (.D(_0060_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][16] ),
    .QN(_1407_));
 DFF_X1 \transfer_count[0][17]$_SDFF_PN0_  (.D(_0061_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][17] ),
    .QN(_1406_));
 DFF_X1 \transfer_count[0][18]$_SDFF_PN0_  (.D(_0062_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][18] ),
    .QN(_1405_));
 DFF_X1 \transfer_count[0][19]$_SDFF_PN0_  (.D(_0063_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][19] ),
    .QN(_1404_));
 DFF_X2 \transfer_count[0][1]$_SDFF_PN0_  (.D(_0064_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][1] ),
    .QN(_1403_));
 DFF_X1 \transfer_count[0][20]$_SDFF_PN0_  (.D(_0065_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][20] ),
    .QN(_1402_));
 DFF_X1 \transfer_count[0][21]$_SDFF_PN0_  (.D(_0066_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][21] ),
    .QN(_1401_));
 DFF_X1 \transfer_count[0][22]$_SDFF_PN0_  (.D(_0067_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][22] ),
    .QN(_1400_));
 DFF_X1 \transfer_count[0][23]$_SDFF_PN0_  (.D(_0068_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][23] ),
    .QN(_1399_));
 DFF_X1 \transfer_count[0][24]$_SDFF_PN0_  (.D(_0069_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][24] ),
    .QN(_1398_));
 DFF_X1 \transfer_count[0][25]$_SDFF_PN0_  (.D(_0070_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][25] ),
    .QN(_1397_));
 DFF_X1 \transfer_count[0][26]$_SDFF_PN0_  (.D(_0071_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][26] ),
    .QN(_1396_));
 DFF_X1 \transfer_count[0][27]$_SDFF_PN0_  (.D(_0072_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][27] ),
    .QN(_1395_));
 DFF_X1 \transfer_count[0][28]$_SDFF_PN0_  (.D(_0073_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][28] ),
    .QN(_1394_));
 DFF_X1 \transfer_count[0][29]$_SDFF_PN0_  (.D(_0074_),
    .CK(clknet_4_6_0_clk),
    .Q(\transfer_count[0][29] ),
    .QN(_1393_));
 DFF_X1 \transfer_count[0][2]$_SDFF_PN0_  (.D(_0075_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][2] ),
    .QN(_1392_));
 DFF_X1 \transfer_count[0][30]$_SDFF_PN0_  (.D(_0076_),
    .CK(clknet_4_7_0_clk),
    .Q(\transfer_count[0][30] ),
    .QN(_1391_));
 DFF_X1 \transfer_count[0][31]$_SDFF_PN0_  (.D(_0077_),
    .CK(clknet_4_4_0_clk),
    .Q(\transfer_count[0][31] ),
    .QN(_1390_));
 DFF_X1 \transfer_count[0][3]$_SDFF_PN0_  (.D(_0078_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][3] ),
    .QN(_1389_));
 DFF_X1 \transfer_count[0][4]$_SDFF_PN0_  (.D(_0079_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][4] ),
    .QN(_1388_));
 DFF_X1 \transfer_count[0][5]$_SDFF_PN0_  (.D(_0080_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][5] ),
    .QN(_1387_));
 DFF_X1 \transfer_count[0][6]$_SDFF_PN0_  (.D(_0081_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][6] ),
    .QN(_1386_));
 DFF_X1 \transfer_count[0][7]$_SDFF_PN0_  (.D(_0082_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][7] ),
    .QN(_1385_));
 DFF_X1 \transfer_count[0][8]$_SDFF_PN0_  (.D(_0083_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][8] ),
    .QN(_1384_));
 DFF_X1 \transfer_count[0][9]$_SDFF_PN0_  (.D(_0084_),
    .CK(clknet_4_5_0_clk),
    .Q(\transfer_count[0][9] ),
    .QN(_1383_));
 DFF_X2 \transfer_count[1][0]$_SDFF_PN0_  (.D(_0085_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][0] ),
    .QN(_1660_));
 DFF_X2 \transfer_count[1][10]$_SDFF_PN0_  (.D(_0086_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][10] ),
    .QN(_1382_));
 DFF_X1 \transfer_count[1][11]$_SDFF_PN0_  (.D(_0087_),
    .CK(clknet_4_0_0_clk),
    .Q(\transfer_count[1][11] ),
    .QN(_1381_));
 DFF_X1 \transfer_count[1][12]$_SDFF_PN0_  (.D(_0088_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][12] ),
    .QN(_1380_));
 DFF_X2 \transfer_count[1][13]$_SDFF_PN0_  (.D(_0089_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][13] ),
    .QN(_1379_));
 DFF_X1 \transfer_count[1][14]$_SDFF_PN0_  (.D(_0090_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][14] ),
    .QN(_1378_));
 DFF_X1 \transfer_count[1][15]$_SDFF_PN0_  (.D(_0091_),
    .CK(clknet_4_0_0_clk),
    .Q(\transfer_count[1][15] ),
    .QN(_1377_));
 DFF_X1 \transfer_count[1][16]$_SDFF_PN0_  (.D(_0092_),
    .CK(clknet_4_0_0_clk),
    .Q(\transfer_count[1][16] ),
    .QN(_1376_));
 DFF_X1 \transfer_count[1][17]$_SDFF_PN0_  (.D(_0093_),
    .CK(clknet_4_0_0_clk),
    .Q(\transfer_count[1][17] ),
    .QN(_1375_));
 DFF_X1 \transfer_count[1][18]$_SDFF_PN0_  (.D(_0094_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][18] ),
    .QN(_1374_));
 DFF_X2 \transfer_count[1][19]$_SDFF_PN0_  (.D(_0095_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][19] ),
    .QN(_1373_));
 DFF_X2 \transfer_count[1][1]$_SDFF_PN0_  (.D(_0096_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][1] ),
    .QN(_1372_));
 DFF_X1 \transfer_count[1][20]$_SDFF_PN0_  (.D(_0097_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][20] ),
    .QN(_1371_));
 DFF_X1 \transfer_count[1][21]$_SDFF_PN0_  (.D(_0098_),
    .CK(clknet_4_0_0_clk),
    .Q(\transfer_count[1][21] ),
    .QN(_1370_));
 DFF_X1 \transfer_count[1][22]$_SDFF_PN0_  (.D(_0099_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][22] ),
    .QN(_1369_));
 DFF_X1 \transfer_count[1][23]$_SDFF_PN0_  (.D(_0100_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][23] ),
    .QN(_1368_));
 DFF_X1 \transfer_count[1][24]$_SDFF_PN0_  (.D(_0101_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][24] ),
    .QN(_1367_));
 DFF_X1 \transfer_count[1][25]$_SDFF_PN0_  (.D(_0102_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][25] ),
    .QN(_1366_));
 DFF_X1 \transfer_count[1][26]$_SDFF_PN0_  (.D(_0103_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][26] ),
    .QN(_1365_));
 DFF_X1 \transfer_count[1][27]$_SDFF_PN0_  (.D(_0104_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][27] ),
    .QN(_1364_));
 DFF_X1 \transfer_count[1][28]$_SDFF_PN0_  (.D(_0105_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][28] ),
    .QN(_1363_));
 DFF_X2 \transfer_count[1][29]$_SDFF_PN0_  (.D(_0106_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][29] ),
    .QN(_1362_));
 DFF_X1 \transfer_count[1][2]$_SDFF_PN0_  (.D(_0107_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][2] ),
    .QN(_1361_));
 DFF_X1 \transfer_count[1][30]$_SDFF_PN0_  (.D(_0108_),
    .CK(clknet_4_3_0_clk),
    .Q(\transfer_count[1][30] ),
    .QN(_1360_));
 DFF_X1 \transfer_count[1][31]$_SDFF_PN0_  (.D(_0109_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][31] ),
    .QN(_1359_));
 DFF_X1 \transfer_count[1][3]$_SDFF_PN0_  (.D(_0110_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][3] ),
    .QN(_1358_));
 DFF_X1 \transfer_count[1][4]$_SDFF_PN0_  (.D(_0111_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][4] ),
    .QN(_1357_));
 DFF_X1 \transfer_count[1][5]$_SDFF_PN0_  (.D(_0112_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][5] ),
    .QN(_1356_));
 DFF_X1 \transfer_count[1][6]$_SDFF_PN0_  (.D(_0113_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][6] ),
    .QN(_1355_));
 DFF_X1 \transfer_count[1][7]$_SDFF_PN0_  (.D(_0114_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][7] ),
    .QN(_1354_));
 DFF_X1 \transfer_count[1][8]$_SDFF_PN0_  (.D(_0115_),
    .CK(clknet_4_1_0_clk),
    .Q(\transfer_count[1][8] ),
    .QN(_1353_));
 DFF_X2 \transfer_count[1][9]$_SDFF_PN0_  (.D(_0116_),
    .CK(clknet_4_2_0_clk),
    .Q(\transfer_count[1][9] ),
    .QN(_1352_));
 DFF_X2 \transfer_count[2][0]$_SDFF_PN0_  (.D(_0117_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][0] ),
    .QN(_1466_));
 DFF_X1 \transfer_count[2][10]$_SDFF_PN0_  (.D(_0118_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][10] ),
    .QN(_1351_));
 DFF_X2 \transfer_count[2][11]$_SDFF_PN0_  (.D(_0119_),
    .CK(clknet_4_13_0_clk),
    .Q(\transfer_count[2][11] ),
    .QN(_1350_));
 DFF_X1 \transfer_count[2][12]$_SDFF_PN0_  (.D(_0120_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][12] ),
    .QN(_1349_));
 DFF_X1 \transfer_count[2][13]$_SDFF_PN0_  (.D(_0121_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][13] ),
    .QN(_1348_));
 DFF_X1 \transfer_count[2][14]$_SDFF_PN0_  (.D(_0122_),
    .CK(clknet_4_13_0_clk),
    .Q(\transfer_count[2][14] ),
    .QN(_1347_));
 DFF_X1 \transfer_count[2][15]$_SDFF_PN0_  (.D(_0123_),
    .CK(clknet_4_13_0_clk),
    .Q(\transfer_count[2][15] ),
    .QN(_1346_));
 DFF_X1 \transfer_count[2][16]$_SDFF_PN0_  (.D(_0124_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][16] ),
    .QN(_1345_));
 DFF_X1 \transfer_count[2][17]$_SDFF_PN0_  (.D(_0125_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][17] ),
    .QN(_1344_));
 DFF_X1 \transfer_count[2][18]$_SDFF_PN0_  (.D(_0126_),
    .CK(clknet_4_13_0_clk),
    .Q(\transfer_count[2][18] ),
    .QN(_1343_));
 DFF_X1 \transfer_count[2][19]$_SDFF_PN0_  (.D(_0127_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][19] ),
    .QN(_1342_));
 DFF_X2 \transfer_count[2][1]$_SDFF_PN0_  (.D(_0128_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][1] ),
    .QN(_1341_));
 DFF_X1 \transfer_count[2][20]$_SDFF_PN0_  (.D(_0129_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][20] ),
    .QN(_1340_));
 DFF_X1 \transfer_count[2][21]$_SDFF_PN0_  (.D(_0130_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][21] ),
    .QN(_1339_));
 DFF_X2 \transfer_count[2][22]$_SDFF_PN0_  (.D(_0131_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][22] ),
    .QN(_1338_));
 DFF_X2 \transfer_count[2][23]$_SDFF_PN0_  (.D(_0132_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][23] ),
    .QN(_1337_));
 DFF_X1 \transfer_count[2][24]$_SDFF_PN0_  (.D(_0133_),
    .CK(clknet_4_14_0_clk),
    .Q(\transfer_count[2][24] ),
    .QN(_1336_));
 DFF_X2 \transfer_count[2][25]$_SDFF_PN0_  (.D(_0134_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][25] ),
    .QN(_1335_));
 DFF_X1 \transfer_count[2][26]$_SDFF_PN0_  (.D(_0135_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][26] ),
    .QN(_1334_));
 DFF_X1 \transfer_count[2][27]$_SDFF_PN0_  (.D(_0136_),
    .CK(clknet_4_13_0_clk),
    .Q(\transfer_count[2][27] ),
    .QN(_1333_));
 DFF_X1 \transfer_count[2][28]$_SDFF_PN0_  (.D(_0137_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][28] ),
    .QN(_1332_));
 DFF_X1 \transfer_count[2][29]$_SDFF_PN0_  (.D(_0138_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][29] ),
    .QN(_1331_));
 DFF_X1 \transfer_count[2][2]$_SDFF_PN0_  (.D(_0139_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][2] ),
    .QN(_1330_));
 DFF_X1 \transfer_count[2][30]$_SDFF_PN0_  (.D(_0140_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][30] ),
    .QN(_1329_));
 DFF_X1 \transfer_count[2][31]$_SDFF_PN0_  (.D(_0141_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][31] ),
    .QN(_1328_));
 DFF_X1 \transfer_count[2][3]$_SDFF_PN0_  (.D(_0142_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][3] ),
    .QN(_1327_));
 DFF_X1 \transfer_count[2][4]$_SDFF_PN0_  (.D(_0143_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][4] ),
    .QN(_1326_));
 DFF_X1 \transfer_count[2][5]$_SDFF_PN0_  (.D(_0144_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][5] ),
    .QN(_1325_));
 DFF_X2 \transfer_count[2][6]$_SDFF_PN0_  (.D(_0145_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][6] ),
    .QN(_1324_));
 DFF_X1 \transfer_count[2][7]$_SDFF_PN0_  (.D(_0146_),
    .CK(clknet_4_12_0_clk),
    .Q(\transfer_count[2][7] ),
    .QN(_1323_));
 DFF_X1 \transfer_count[2][8]$_SDFF_PN0_  (.D(_0147_),
    .CK(clknet_4_15_0_clk),
    .Q(\transfer_count[2][8] ),
    .QN(_1322_));
 DFF_X1 \transfer_count[2][9]$_SDFF_PN0_  (.D(_0148_),
    .CK(clknet_4_13_0_clk),
    .Q(\transfer_count[2][9] ),
    .QN(_1321_));
 DFF_X1 \transfer_count[3][0]$_SDFF_PN0_  (.D(_0149_),
    .CK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][0] ),
    .QN(_1763_));
 DFF_X1 \transfer_count[3][10]$_SDFF_PN0_  (.D(_0150_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][10] ),
    .QN(_1320_));
 DFF_X1 \transfer_count[3][11]$_SDFF_PN0_  (.D(_0151_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][11] ),
    .QN(_1319_));
 DFF_X2 \transfer_count[3][12]$_SDFF_PN0_  (.D(_0152_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][12] ),
    .QN(_1318_));
 DFF_X1 \transfer_count[3][13]$_SDFF_PN0_  (.D(_0153_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][13] ),
    .QN(_1317_));
 DFF_X1 \transfer_count[3][14]$_SDFF_PN0_  (.D(_0154_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][14] ),
    .QN(_1316_));
 DFF_X1 \transfer_count[3][15]$_SDFF_PN0_  (.D(_0155_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][15] ),
    .QN(_1315_));
 DFF_X1 \transfer_count[3][16]$_SDFF_PN0_  (.D(_0156_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][16] ),
    .QN(_1314_));
 DFF_X1 \transfer_count[3][17]$_SDFF_PN0_  (.D(_0157_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][17] ),
    .QN(_1313_));
 DFF_X1 \transfer_count[3][18]$_SDFF_PN0_  (.D(_0158_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][18] ),
    .QN(_1312_));
 DFF_X1 \transfer_count[3][19]$_SDFF_PN0_  (.D(_0159_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][19] ),
    .QN(_1311_));
 DFF_X1 \transfer_count[3][1]$_SDFF_PN0_  (.D(_0160_),
    .CK(clknet_4_8_0_clk),
    .Q(\transfer_count[3][1] ),
    .QN(_1310_));
 DFF_X1 \transfer_count[3][20]$_SDFF_PN0_  (.D(_0161_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][20] ),
    .QN(_1309_));
 DFF_X1 \transfer_count[3][21]$_SDFF_PN0_  (.D(_0162_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][21] ),
    .QN(_1308_));
 DFF_X1 \transfer_count[3][22]$_SDFF_PN0_  (.D(_0163_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][22] ),
    .QN(_1307_));
 DFF_X1 \transfer_count[3][23]$_SDFF_PN0_  (.D(_0164_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][23] ),
    .QN(_1306_));
 DFF_X1 \transfer_count[3][24]$_SDFF_PN0_  (.D(_0165_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][24] ),
    .QN(_1305_));
 DFF_X1 \transfer_count[3][25]$_SDFF_PN0_  (.D(_0166_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][25] ),
    .QN(_1304_));
 DFF_X1 \transfer_count[3][26]$_SDFF_PN0_  (.D(_0167_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][26] ),
    .QN(_1303_));
 DFF_X1 \transfer_count[3][27]$_SDFF_PN0_  (.D(_0168_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][27] ),
    .QN(_1302_));
 DFF_X1 \transfer_count[3][28]$_SDFF_PN0_  (.D(_0169_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][28] ),
    .QN(_1301_));
 DFF_X1 \transfer_count[3][29]$_SDFF_PN0_  (.D(_0170_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][29] ),
    .QN(_1300_));
 DFF_X1 \transfer_count[3][2]$_SDFF_PN0_  (.D(_0171_),
    .CK(clknet_4_9_0_clk),
    .Q(\transfer_count[3][2] ),
    .QN(_1299_));
 DFF_X1 \transfer_count[3][30]$_SDFF_PN0_  (.D(_0172_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][30] ),
    .QN(_1298_));
 DFF_X1 \transfer_count[3][31]$_SDFF_PN0_  (.D(_0173_),
    .CK(clknet_4_10_0_clk),
    .Q(\transfer_count[3][31] ),
    .QN(_1297_));
 DFF_X1 \transfer_count[3][3]$_SDFF_PN0_  (.D(_0174_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][3] ),
    .QN(_1296_));
 DFF_X1 \transfer_count[3][4]$_SDFF_PN0_  (.D(_0175_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][4] ),
    .QN(_1295_));
 DFF_X1 \transfer_count[3][5]$_SDFF_PN0_  (.D(_0176_),
    .CK(clknet_4_9_0_clk),
    .Q(\transfer_count[3][5] ),
    .QN(_1294_));
 DFF_X2 \transfer_count[3][6]$_SDFF_PN0_  (.D(_0177_),
    .CK(clknet_4_9_0_clk),
    .Q(\transfer_count[3][6] ),
    .QN(_1293_));
 DFF_X1 \transfer_count[3][7]$_SDFF_PN0_  (.D(_0178_),
    .CK(clknet_4_9_0_clk),
    .Q(\transfer_count[3][7] ),
    .QN(_1292_));
 DFF_X1 \transfer_count[3][8]$_SDFF_PN0_  (.D(_0179_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][8] ),
    .QN(_1291_));
 DFF_X1 \transfer_count[3][9]$_SDFF_PN0_  (.D(_0180_),
    .CK(clknet_4_11_0_clk),
    .Q(\transfer_count[3][9] ),
    .QN(_1290_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_427 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_428 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_429 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_430 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_431 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_432 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_433 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_434 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_435 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_436 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_541 ();
 BUF_X1 input1 (.A(channel_length[0]),
    .Z(net1));
 BUF_X2 input2 (.A(channel_length[100]),
    .Z(net2));
 BUF_X2 input3 (.A(channel_length[101]),
    .Z(net3));
 BUF_X2 input4 (.A(channel_length[102]),
    .Z(net4));
 BUF_X2 input5 (.A(channel_length[103]),
    .Z(net5));
 BUF_X2 input6 (.A(channel_length[104]),
    .Z(net6));
 BUF_X2 input7 (.A(channel_length[105]),
    .Z(net7));
 BUF_X2 input8 (.A(channel_length[106]),
    .Z(net8));
 BUF_X2 input9 (.A(channel_length[107]),
    .Z(net9));
 BUF_X2 input10 (.A(channel_length[108]),
    .Z(net10));
 CLKBUF_X2 input11 (.A(channel_length[109]),
    .Z(net11));
 BUF_X1 input12 (.A(channel_length[10]),
    .Z(net12));
 CLKBUF_X2 input13 (.A(channel_length[110]),
    .Z(net13));
 BUF_X2 input14 (.A(channel_length[111]),
    .Z(net14));
 BUF_X1 input15 (.A(channel_length[112]),
    .Z(net15));
 BUF_X1 input16 (.A(channel_length[113]),
    .Z(net16));
 BUF_X1 input17 (.A(channel_length[114]),
    .Z(net17));
 BUF_X1 input18 (.A(channel_length[115]),
    .Z(net18));
 CLKBUF_X2 input19 (.A(channel_length[116]),
    .Z(net19));
 CLKBUF_X2 input20 (.A(channel_length[117]),
    .Z(net20));
 CLKBUF_X2 input21 (.A(channel_length[118]),
    .Z(net21));
 CLKBUF_X2 input22 (.A(channel_length[119]),
    .Z(net22));
 BUF_X1 input23 (.A(channel_length[11]),
    .Z(net23));
 BUF_X2 input24 (.A(channel_length[120]),
    .Z(net24));
 BUF_X2 input25 (.A(channel_length[121]),
    .Z(net25));
 BUF_X2 input26 (.A(channel_length[122]),
    .Z(net26));
 BUF_X2 input27 (.A(channel_length[123]),
    .Z(net27));
 CLKBUF_X2 input28 (.A(channel_length[124]),
    .Z(net28));
 CLKBUF_X2 input29 (.A(channel_length[125]),
    .Z(net29));
 CLKBUF_X2 input30 (.A(channel_length[126]),
    .Z(net30));
 CLKBUF_X2 input31 (.A(channel_length[127]),
    .Z(net31));
 BUF_X1 input32 (.A(channel_length[12]),
    .Z(net32));
 BUF_X1 input33 (.A(channel_length[13]),
    .Z(net33));
 BUF_X1 input34 (.A(channel_length[14]),
    .Z(net34));
 BUF_X1 input35 (.A(channel_length[15]),
    .Z(net35));
 BUF_X1 input36 (.A(channel_length[16]),
    .Z(net36));
 BUF_X1 input37 (.A(channel_length[17]),
    .Z(net37));
 BUF_X1 input38 (.A(channel_length[18]),
    .Z(net38));
 BUF_X1 input39 (.A(channel_length[19]),
    .Z(net39));
 BUF_X1 input40 (.A(channel_length[1]),
    .Z(net40));
 BUF_X1 input41 (.A(channel_length[20]),
    .Z(net41));
 BUF_X1 input42 (.A(channel_length[21]),
    .Z(net42));
 BUF_X1 input43 (.A(channel_length[22]),
    .Z(net43));
 BUF_X1 input44 (.A(channel_length[23]),
    .Z(net44));
 BUF_X1 input45 (.A(channel_length[24]),
    .Z(net45));
 BUF_X1 input46 (.A(channel_length[25]),
    .Z(net46));
 BUF_X1 input47 (.A(channel_length[26]),
    .Z(net47));
 BUF_X1 input48 (.A(channel_length[27]),
    .Z(net48));
 BUF_X1 input49 (.A(channel_length[28]),
    .Z(net49));
 BUF_X1 input50 (.A(channel_length[29]),
    .Z(net50));
 BUF_X1 input51 (.A(channel_length[2]),
    .Z(net51));
 BUF_X1 input52 (.A(channel_length[30]),
    .Z(net52));
 BUF_X1 input53 (.A(channel_length[31]),
    .Z(net53));
 BUF_X1 input54 (.A(channel_length[32]),
    .Z(net54));
 BUF_X1 input55 (.A(channel_length[33]),
    .Z(net55));
 BUF_X1 input56 (.A(channel_length[34]),
    .Z(net56));
 BUF_X1 input57 (.A(channel_length[35]),
    .Z(net57));
 BUF_X1 input58 (.A(channel_length[36]),
    .Z(net58));
 BUF_X1 input59 (.A(channel_length[37]),
    .Z(net59));
 BUF_X1 input60 (.A(channel_length[38]),
    .Z(net60));
 BUF_X1 input61 (.A(channel_length[39]),
    .Z(net61));
 BUF_X1 input62 (.A(channel_length[3]),
    .Z(net62));
 BUF_X1 input63 (.A(channel_length[40]),
    .Z(net63));
 BUF_X1 input64 (.A(channel_length[41]),
    .Z(net64));
 BUF_X1 input65 (.A(channel_length[42]),
    .Z(net65));
 BUF_X1 input66 (.A(channel_length[43]),
    .Z(net66));
 BUF_X1 input67 (.A(channel_length[44]),
    .Z(net67));
 BUF_X1 input68 (.A(channel_length[45]),
    .Z(net68));
 BUF_X1 input69 (.A(channel_length[46]),
    .Z(net69));
 BUF_X1 input70 (.A(channel_length[47]),
    .Z(net70));
 BUF_X1 input71 (.A(channel_length[48]),
    .Z(net71));
 BUF_X1 input72 (.A(channel_length[49]),
    .Z(net72));
 BUF_X1 input73 (.A(channel_length[4]),
    .Z(net73));
 BUF_X1 input74 (.A(channel_length[50]),
    .Z(net74));
 BUF_X1 input75 (.A(channel_length[51]),
    .Z(net75));
 BUF_X1 input76 (.A(channel_length[52]),
    .Z(net76));
 BUF_X1 input77 (.A(channel_length[53]),
    .Z(net77));
 BUF_X1 input78 (.A(channel_length[54]),
    .Z(net78));
 BUF_X1 input79 (.A(channel_length[55]),
    .Z(net79));
 BUF_X1 input80 (.A(channel_length[56]),
    .Z(net80));
 BUF_X1 input81 (.A(channel_length[57]),
    .Z(net81));
 BUF_X1 input82 (.A(channel_length[58]),
    .Z(net82));
 BUF_X1 input83 (.A(channel_length[59]),
    .Z(net83));
 BUF_X1 input84 (.A(channel_length[5]),
    .Z(net84));
 BUF_X1 input85 (.A(channel_length[60]),
    .Z(net85));
 BUF_X1 input86 (.A(channel_length[61]),
    .Z(net86));
 BUF_X1 input87 (.A(channel_length[62]),
    .Z(net87));
 BUF_X1 input88 (.A(channel_length[63]),
    .Z(net88));
 BUF_X1 input89 (.A(channel_length[64]),
    .Z(net89));
 BUF_X1 input90 (.A(channel_length[65]),
    .Z(net90));
 BUF_X1 input91 (.A(channel_length[66]),
    .Z(net91));
 BUF_X1 input92 (.A(channel_length[67]),
    .Z(net92));
 BUF_X1 input93 (.A(channel_length[68]),
    .Z(net93));
 BUF_X1 input94 (.A(channel_length[69]),
    .Z(net94));
 BUF_X1 input95 (.A(channel_length[6]),
    .Z(net95));
 BUF_X1 input96 (.A(channel_length[70]),
    .Z(net96));
 BUF_X1 input97 (.A(channel_length[71]),
    .Z(net97));
 BUF_X1 input98 (.A(channel_length[72]),
    .Z(net98));
 BUF_X1 input99 (.A(channel_length[73]),
    .Z(net99));
 BUF_X1 input100 (.A(channel_length[74]),
    .Z(net100));
 BUF_X1 input101 (.A(channel_length[75]),
    .Z(net101));
 BUF_X1 input102 (.A(channel_length[76]),
    .Z(net102));
 BUF_X1 input103 (.A(channel_length[77]),
    .Z(net103));
 BUF_X1 input104 (.A(channel_length[78]),
    .Z(net104));
 BUF_X1 input105 (.A(channel_length[79]),
    .Z(net105));
 BUF_X1 input106 (.A(channel_length[7]),
    .Z(net106));
 BUF_X1 input107 (.A(channel_length[80]),
    .Z(net107));
 BUF_X1 input108 (.A(channel_length[81]),
    .Z(net108));
 BUF_X1 input109 (.A(channel_length[82]),
    .Z(net109));
 BUF_X1 input110 (.A(channel_length[83]),
    .Z(net110));
 BUF_X1 input111 (.A(channel_length[84]),
    .Z(net111));
 BUF_X1 input112 (.A(channel_length[85]),
    .Z(net112));
 BUF_X1 input113 (.A(channel_length[86]),
    .Z(net113));
 BUF_X1 input114 (.A(channel_length[87]),
    .Z(net114));
 BUF_X1 input115 (.A(channel_length[88]),
    .Z(net115));
 BUF_X1 input116 (.A(channel_length[89]),
    .Z(net116));
 BUF_X1 input117 (.A(channel_length[8]),
    .Z(net117));
 BUF_X1 input118 (.A(channel_length[90]),
    .Z(net118));
 BUF_X1 input119 (.A(channel_length[91]),
    .Z(net119));
 BUF_X1 input120 (.A(channel_length[92]),
    .Z(net120));
 BUF_X2 input121 (.A(channel_length[93]),
    .Z(net121));
 BUF_X2 input122 (.A(channel_length[94]),
    .Z(net122));
 BUF_X1 input123 (.A(channel_length[95]),
    .Z(net123));
 BUF_X1 input124 (.A(channel_length[96]),
    .Z(net124));
 BUF_X2 input125 (.A(channel_length[97]),
    .Z(net125));
 BUF_X2 input126 (.A(channel_length[98]),
    .Z(net126));
 BUF_X2 input127 (.A(channel_length[99]),
    .Z(net127));
 BUF_X2 input128 (.A(channel_length[9]),
    .Z(net128));
 CLKBUF_X3 input129 (.A(channel_start[2]),
    .Z(net129));
 CLKBUF_X2 input130 (.A(dst_wready[0]),
    .Z(net130));
 BUF_X1 input131 (.A(dst_wready[1]),
    .Z(net131));
 CLKBUF_X3 input132 (.A(dst_wready[2]),
    .Z(net132));
 CLKBUF_X3 input133 (.A(dst_wready[3]),
    .Z(net133));
 BUF_X1 input134 (.A(src_rvalid[0]),
    .Z(net134));
 BUF_X1 input135 (.A(src_rvalid[1]),
    .Z(net135));
 BUF_X1 input136 (.A(src_rvalid[2]),
    .Z(net136));
 BUF_X2 input137 (.A(src_rvalid[3]),
    .Z(net137));
 BUF_X1 output138 (.A(net138),
    .Z(channel_busy[0]));
 BUF_X1 output139 (.A(net139),
    .Z(channel_busy[1]));
 BUF_X1 output140 (.A(net140),
    .Z(channel_busy[2]));
 BUF_X1 output141 (.A(net141),
    .Z(channel_busy[3]));
 BUF_X1 output142 (.A(net142),
    .Z(channel_done[0]));
 BUF_X1 output143 (.A(net143),
    .Z(channel_done[1]));
 BUF_X1 output144 (.A(net144),
    .Z(channel_done[2]));
 BUF_X1 output145 (.A(net145),
    .Z(channel_done[3]));
 BUF_X1 output146 (.A(net146),
    .Z(debug_active_channels[0]));
 BUF_X1 output147 (.A(net147),
    .Z(debug_active_channels[1]));
 BUF_X1 output148 (.A(net148),
    .Z(debug_active_channels[2]));
 BUF_X1 output149 (.A(net149),
    .Z(debug_active_channels[3]));
 BUF_X1 output150 (.A(net150),
    .Z(debug_has_active_channels));
 BUF_X1 output151 (.A(net151),
    .Z(dst_write[0]));
 BUF_X1 output152 (.A(net152),
    .Z(dst_write[1]));
 BUF_X1 output153 (.A(net153),
    .Z(dst_write[2]));
 BUF_X1 output154 (.A(net154),
    .Z(dst_write[3]));
 BUF_X1 output155 (.A(net155),
    .Z(src_read[0]));
 BUF_X1 output156 (.A(net156),
    .Z(src_read[1]));
 BUF_X1 output157 (.A(net157),
    .Z(src_read[2]));
 BUF_X1 output158 (.A(net158),
    .Z(src_read[3]));
 BUF_X1 output159 (.A(net159),
    .Z(src_rready[0]));
 BUF_X1 output160 (.A(net160),
    .Z(src_rready[1]));
 BUF_X1 output161 (.A(net161),
    .Z(src_rready[2]));
 BUF_X1 output162 (.A(net162),
    .Z(src_rready[3]));
 LOGIC0_X1 _3421__163 (.Z(net163));
 LOGIC0_X1 _3422__164 (.Z(net164));
 LOGIC0_X1 _3423__165 (.Z(net165));
 LOGIC0_X1 _3424__166 (.Z(net166));
 LOGIC0_X1 _3425__167 (.Z(net167));
 LOGIC0_X1 _3426__168 (.Z(net168));
 LOGIC0_X1 _3427__169 (.Z(net169));
 LOGIC0_X1 _3428__170 (.Z(net170));
 LOGIC0_X1 _3429__171 (.Z(net171));
 LOGIC0_X1 _3430__172 (.Z(net172));
 LOGIC0_X1 _3431__173 (.Z(net173));
 LOGIC0_X1 _3432__174 (.Z(net174));
 LOGIC0_X1 _3433__175 (.Z(net175));
 LOGIC0_X1 _3434__176 (.Z(net176));
 LOGIC0_X1 _3435__177 (.Z(net177));
 LOGIC0_X1 _3436__178 (.Z(net178));
 LOGIC0_X1 _3437__179 (.Z(net179));
 LOGIC0_X1 _3438__180 (.Z(net180));
 LOGIC0_X1 _3439__181 (.Z(net181));
 LOGIC0_X1 _3440__182 (.Z(net182));
 LOGIC0_X1 _3441__183 (.Z(net183));
 LOGIC0_X1 _3442__184 (.Z(net184));
 LOGIC0_X1 _3443__185 (.Z(net185));
 LOGIC0_X1 _3444__186 (.Z(net186));
 LOGIC0_X1 _3445__187 (.Z(net187));
 LOGIC0_X1 _3446__188 (.Z(net188));
 LOGIC0_X1 _3447__189 (.Z(net189));
 LOGIC0_X1 _3448__190 (.Z(net190));
 LOGIC0_X1 _3449__191 (.Z(net191));
 LOGIC0_X1 _3450__192 (.Z(net192));
 LOGIC0_X1 _3451__193 (.Z(net193));
 LOGIC0_X1 _3452__194 (.Z(net194));
 LOGIC0_X1 _3453__195 (.Z(net195));
 LOGIC0_X1 _3454__196 (.Z(net196));
 LOGIC0_X1 _3455__197 (.Z(net197));
 LOGIC0_X1 _3456__198 (.Z(net198));
 LOGIC0_X1 _3457__199 (.Z(net199));
 LOGIC0_X1 _3458__200 (.Z(net200));
 LOGIC0_X1 _3459__201 (.Z(net201));
 LOGIC0_X1 _3460__202 (.Z(net202));
 LOGIC0_X1 _3461__203 (.Z(net203));
 LOGIC0_X1 _3462__204 (.Z(net204));
 LOGIC0_X1 _3463__205 (.Z(net205));
 LOGIC0_X1 _3464__206 (.Z(net206));
 LOGIC0_X1 _3465__207 (.Z(net207));
 LOGIC0_X1 _3466__208 (.Z(net208));
 LOGIC0_X1 _3467__209 (.Z(net209));
 LOGIC0_X1 _3468__210 (.Z(net210));
 LOGIC0_X1 _3469__211 (.Z(net211));
 LOGIC0_X1 _3470__212 (.Z(net212));
 LOGIC0_X1 _3471__213 (.Z(net213));
 LOGIC0_X1 _3472__214 (.Z(net214));
 LOGIC0_X1 _3473__215 (.Z(net215));
 LOGIC0_X1 _3474__216 (.Z(net216));
 LOGIC0_X1 _3475__217 (.Z(net217));
 LOGIC0_X1 _3476__218 (.Z(net218));
 LOGIC0_X1 _3477__219 (.Z(net219));
 LOGIC0_X1 _3478__220 (.Z(net220));
 LOGIC0_X1 _3479__221 (.Z(net221));
 LOGIC0_X1 _3480__222 (.Z(net222));
 LOGIC0_X1 _3481__223 (.Z(net223));
 LOGIC0_X1 _3482__224 (.Z(net224));
 LOGIC0_X1 _3483__225 (.Z(net225));
 LOGIC0_X1 _3484__226 (.Z(net226));
 LOGIC0_X1 _3485__227 (.Z(net227));
 LOGIC0_X1 _3486__228 (.Z(net228));
 LOGIC0_X1 _3487__229 (.Z(net229));
 LOGIC0_X1 _3488__230 (.Z(net230));
 LOGIC0_X1 _3489__231 (.Z(net231));
 LOGIC0_X1 _3490__232 (.Z(net232));
 LOGIC0_X1 _3491__233 (.Z(net233));
 LOGIC0_X1 _3492__234 (.Z(net234));
 LOGIC0_X1 _3493__235 (.Z(net235));
 LOGIC0_X1 _3494__236 (.Z(net236));
 LOGIC0_X1 _3495__237 (.Z(net237));
 LOGIC0_X1 _3496__238 (.Z(net238));
 LOGIC0_X1 _3497__239 (.Z(net239));
 LOGIC0_X1 _3498__240 (.Z(net240));
 LOGIC0_X1 _3499__241 (.Z(net241));
 LOGIC0_X1 _3500__242 (.Z(net242));
 LOGIC0_X1 _3501__243 (.Z(net243));
 LOGIC0_X1 _3502__244 (.Z(net244));
 LOGIC0_X1 _3503__245 (.Z(net245));
 LOGIC0_X1 _3504__246 (.Z(net246));
 LOGIC0_X1 _3505__247 (.Z(net247));
 LOGIC0_X1 _3506__248 (.Z(net248));
 LOGIC0_X1 _3507__249 (.Z(net249));
 LOGIC0_X1 _3508__250 (.Z(net250));
 LOGIC0_X1 _3509__251 (.Z(net251));
 LOGIC0_X1 _3510__252 (.Z(net252));
 LOGIC0_X1 _3511__253 (.Z(net253));
 LOGIC0_X1 _3512__254 (.Z(net254));
 LOGIC0_X1 _3513__255 (.Z(net255));
 LOGIC0_X1 _3514__256 (.Z(net256));
 LOGIC0_X1 _3515__257 (.Z(net257));
 LOGIC0_X1 _3516__258 (.Z(net258));
 LOGIC0_X1 _3517__259 (.Z(net259));
 LOGIC0_X1 _3518__260 (.Z(net260));
 LOGIC0_X1 _3519__261 (.Z(net261));
 LOGIC0_X1 _3520__262 (.Z(net262));
 LOGIC0_X1 _3521__263 (.Z(net263));
 LOGIC0_X1 _3522__264 (.Z(net264));
 LOGIC0_X1 _3523__265 (.Z(net265));
 LOGIC0_X1 _3524__266 (.Z(net266));
 LOGIC0_X1 _3525__267 (.Z(net267));
 LOGIC0_X1 _3526__268 (.Z(net268));
 LOGIC0_X1 _3527__269 (.Z(net269));
 LOGIC0_X1 _3528__270 (.Z(net270));
 LOGIC0_X1 _3529__271 (.Z(net271));
 LOGIC0_X1 _3530__272 (.Z(net272));
 LOGIC0_X1 _3531__273 (.Z(net273));
 LOGIC0_X1 _3532__274 (.Z(net274));
 LOGIC0_X1 _3533__275 (.Z(net275));
 LOGIC0_X1 _3534__276 (.Z(net276));
 LOGIC0_X1 _3535__277 (.Z(net277));
 LOGIC0_X1 _3536__278 (.Z(net278));
 LOGIC0_X1 _3537__279 (.Z(net279));
 LOGIC0_X1 _3538__280 (.Z(net280));
 LOGIC0_X1 _3539__281 (.Z(net281));
 LOGIC0_X1 _3540__282 (.Z(net282));
 LOGIC0_X1 _3541__283 (.Z(net283));
 LOGIC0_X1 _3542__284 (.Z(net284));
 LOGIC0_X1 _3543__285 (.Z(net285));
 LOGIC0_X1 _3544__286 (.Z(net286));
 LOGIC0_X1 _3545__287 (.Z(net287));
 LOGIC0_X1 _3546__288 (.Z(net288));
 LOGIC0_X1 _3547__289 (.Z(net289));
 LOGIC0_X1 _3548__290 (.Z(net290));
 LOGIC0_X1 _3549__291 (.Z(net291));
 LOGIC0_X1 _3550__292 (.Z(net292));
 LOGIC0_X1 _3551__293 (.Z(net293));
 LOGIC0_X1 _3552__294 (.Z(net294));
 LOGIC0_X1 _3553__295 (.Z(net295));
 LOGIC0_X1 _3554__296 (.Z(net296));
 LOGIC0_X1 _3555__297 (.Z(net297));
 LOGIC0_X1 _3556__298 (.Z(net298));
 LOGIC0_X1 _3557__299 (.Z(net299));
 LOGIC0_X1 _3558__300 (.Z(net300));
 LOGIC0_X1 _3559__301 (.Z(net301));
 LOGIC0_X1 _3560__302 (.Z(net302));
 LOGIC0_X1 _3561__303 (.Z(net303));
 LOGIC0_X1 _3562__304 (.Z(net304));
 LOGIC0_X1 _3563__305 (.Z(net305));
 LOGIC0_X1 _3564__306 (.Z(net306));
 LOGIC0_X1 _3565__307 (.Z(net307));
 LOGIC0_X1 _3566__308 (.Z(net308));
 LOGIC0_X1 _3567__309 (.Z(net309));
 LOGIC0_X1 _3568__310 (.Z(net310));
 LOGIC0_X1 _3569__311 (.Z(net311));
 LOGIC0_X1 _3570__312 (.Z(net312));
 LOGIC0_X1 _3571__313 (.Z(net313));
 LOGIC0_X1 _3572__314 (.Z(net314));
 LOGIC0_X1 _3573__315 (.Z(net315));
 LOGIC0_X1 _3574__316 (.Z(net316));
 LOGIC0_X1 _3575__317 (.Z(net317));
 LOGIC0_X1 _3576__318 (.Z(net318));
 LOGIC0_X1 _3577__319 (.Z(net319));
 LOGIC0_X1 _3578__320 (.Z(net320));
 LOGIC0_X1 _3579__321 (.Z(net321));
 LOGIC0_X1 _3580__322 (.Z(net322));
 LOGIC0_X1 _3581__323 (.Z(net323));
 LOGIC0_X1 _3582__324 (.Z(net324));
 LOGIC0_X1 _3583__325 (.Z(net325));
 LOGIC0_X1 _3584__326 (.Z(net326));
 LOGIC0_X1 _3585__327 (.Z(net327));
 LOGIC0_X1 _3586__328 (.Z(net328));
 LOGIC0_X1 _3587__329 (.Z(net329));
 LOGIC0_X1 _3588__330 (.Z(net330));
 LOGIC0_X1 _3589__331 (.Z(net331));
 LOGIC0_X1 _3590__332 (.Z(net332));
 LOGIC0_X1 _3591__333 (.Z(net333));
 LOGIC0_X1 _3592__334 (.Z(net334));
 LOGIC0_X1 _3593__335 (.Z(net335));
 LOGIC0_X1 _3594__336 (.Z(net336));
 LOGIC0_X1 _3595__337 (.Z(net337));
 LOGIC0_X1 _3596__338 (.Z(net338));
 LOGIC0_X1 _3597__339 (.Z(net339));
 LOGIC0_X1 _3598__340 (.Z(net340));
 LOGIC0_X1 _3599__341 (.Z(net341));
 LOGIC0_X1 _3600__342 (.Z(net342));
 LOGIC0_X1 _3601__343 (.Z(net343));
 LOGIC0_X1 _3602__344 (.Z(net344));
 LOGIC0_X1 _3603__345 (.Z(net345));
 LOGIC0_X1 _3604__346 (.Z(net346));
 LOGIC0_X1 _3605__347 (.Z(net347));
 LOGIC0_X1 _3606__348 (.Z(net348));
 LOGIC0_X1 _3607__349 (.Z(net349));
 LOGIC0_X1 _3608__350 (.Z(net350));
 LOGIC0_X1 _3609__351 (.Z(net351));
 LOGIC0_X1 _3610__352 (.Z(net352));
 LOGIC0_X1 _3611__353 (.Z(net353));
 LOGIC0_X1 _3612__354 (.Z(net354));
 LOGIC0_X1 _3613__355 (.Z(net355));
 LOGIC0_X1 _3614__356 (.Z(net356));
 LOGIC0_X1 _3615__357 (.Z(net357));
 LOGIC0_X1 _3616__358 (.Z(net358));
 LOGIC0_X1 _3617__359 (.Z(net359));
 LOGIC0_X1 _3618__360 (.Z(net360));
 LOGIC0_X1 _3619__361 (.Z(net361));
 LOGIC0_X1 _3620__362 (.Z(net362));
 LOGIC0_X1 _3621__363 (.Z(net363));
 LOGIC0_X1 _3622__364 (.Z(net364));
 LOGIC0_X1 _3623__365 (.Z(net365));
 LOGIC0_X1 _3624__366 (.Z(net366));
 LOGIC0_X1 _3625__367 (.Z(net367));
 LOGIC0_X1 _3626__368 (.Z(net368));
 LOGIC0_X1 _3627__369 (.Z(net369));
 LOGIC0_X1 _3628__370 (.Z(net370));
 LOGIC0_X1 _3629__371 (.Z(net371));
 LOGIC0_X1 _3630__372 (.Z(net372));
 LOGIC0_X1 _3631__373 (.Z(net373));
 LOGIC0_X1 _3632__374 (.Z(net374));
 LOGIC0_X1 _3633__375 (.Z(net375));
 LOGIC0_X1 _3634__376 (.Z(net376));
 LOGIC0_X1 _3635__377 (.Z(net377));
 LOGIC0_X1 _3636__378 (.Z(net378));
 LOGIC0_X1 _3637__379 (.Z(net379));
 LOGIC0_X1 _3638__380 (.Z(net380));
 LOGIC0_X1 _3639__381 (.Z(net381));
 LOGIC0_X1 _3640__382 (.Z(net382));
 LOGIC0_X1 _3641__383 (.Z(net383));
 LOGIC0_X1 _3642__384 (.Z(net384));
 LOGIC0_X1 _3643__385 (.Z(net385));
 LOGIC0_X1 _3644__386 (.Z(net386));
 LOGIC0_X1 _3645__387 (.Z(net387));
 LOGIC0_X1 _3646__388 (.Z(net388));
 LOGIC0_X1 _3647__389 (.Z(net389));
 LOGIC0_X1 _3648__390 (.Z(net390));
 LOGIC0_X1 _3649__391 (.Z(net391));
 LOGIC0_X1 _3650__392 (.Z(net392));
 LOGIC0_X1 _3651__393 (.Z(net393));
 LOGIC0_X1 _3652__394 (.Z(net394));
 LOGIC0_X1 _3653__395 (.Z(net395));
 LOGIC0_X1 _3654__396 (.Z(net396));
 LOGIC0_X1 _3655__397 (.Z(net397));
 LOGIC0_X1 _3656__398 (.Z(net398));
 LOGIC0_X1 _3657__399 (.Z(net399));
 LOGIC0_X1 _3658__400 (.Z(net400));
 LOGIC0_X1 _3659__401 (.Z(net401));
 LOGIC0_X1 _3660__402 (.Z(net402));
 LOGIC0_X1 _3661__403 (.Z(net403));
 LOGIC0_X1 _3662__404 (.Z(net404));
 LOGIC0_X1 _3663__405 (.Z(net405));
 LOGIC0_X1 _3664__406 (.Z(net406));
 LOGIC0_X1 _3665__407 (.Z(net407));
 LOGIC0_X1 _3666__408 (.Z(net408));
 LOGIC0_X1 _3667__409 (.Z(net409));
 LOGIC0_X1 _3668__410 (.Z(net410));
 LOGIC0_X1 _3669__411 (.Z(net411));
 LOGIC0_X1 _3670__412 (.Z(net412));
 LOGIC0_X1 _3671__413 (.Z(net413));
 LOGIC0_X1 _3672__414 (.Z(net414));
 LOGIC0_X1 _3673__415 (.Z(net415));
 LOGIC0_X1 _3674__416 (.Z(net416));
 LOGIC0_X1 _3675__417 (.Z(net417));
 LOGIC0_X1 _3676__418 (.Z(net418));
 LOGIC0_X1 _3677__419 (.Z(net419));
 LOGIC0_X1 _3678__420 (.Z(net420));
 LOGIC0_X1 _3679__421 (.Z(net421));
 LOGIC0_X1 _3680__422 (.Z(net422));
 LOGIC0_X1 _3681__423 (.Z(net423));
 LOGIC0_X1 _3682__424 (.Z(net424));
 LOGIC0_X1 _3683__425 (.Z(net425));
 LOGIC0_X1 _3684__426 (.Z(net426));
 LOGIC0_X1 _3685__427 (.Z(net427));
 LOGIC0_X1 _3686__428 (.Z(net428));
 LOGIC0_X1 _3687__429 (.Z(net429));
 LOGIC0_X1 _3688__430 (.Z(net430));
 LOGIC0_X1 _3689__431 (.Z(net431));
 LOGIC0_X1 _3690__432 (.Z(net432));
 LOGIC0_X1 _3691__433 (.Z(net433));
 LOGIC0_X1 _3692__434 (.Z(net434));
 LOGIC0_X1 _3693__435 (.Z(net435));
 LOGIC0_X1 _3694__436 (.Z(net436));
 LOGIC0_X1 _3695__437 (.Z(net437));
 LOGIC0_X1 _3696__438 (.Z(net438));
 LOGIC0_X1 _3697__439 (.Z(net439));
 LOGIC0_X1 _3698__440 (.Z(net440));
 LOGIC0_X1 _3699__441 (.Z(net441));
 LOGIC0_X1 _3700__442 (.Z(net442));
 LOGIC0_X1 _3701__443 (.Z(net443));
 LOGIC0_X1 _3702__444 (.Z(net444));
 LOGIC0_X1 _3703__445 (.Z(net445));
 LOGIC0_X1 _3704__446 (.Z(net446));
 LOGIC0_X1 _3705__447 (.Z(net447));
 LOGIC0_X1 _3706__448 (.Z(net448));
 LOGIC0_X1 _3707__449 (.Z(net449));
 LOGIC0_X1 _3708__450 (.Z(net450));
 LOGIC0_X1 _3709__451 (.Z(net451));
 LOGIC0_X1 _3710__452 (.Z(net452));
 LOGIC0_X1 _3711__453 (.Z(net453));
 LOGIC0_X1 _3712__454 (.Z(net454));
 LOGIC0_X1 _3713__455 (.Z(net455));
 LOGIC0_X1 _3714__456 (.Z(net456));
 LOGIC0_X1 _3715__457 (.Z(net457));
 LOGIC0_X1 _3716__458 (.Z(net458));
 LOGIC0_X1 _3717__459 (.Z(net459));
 LOGIC0_X1 _3718__460 (.Z(net460));
 LOGIC0_X1 _3719__461 (.Z(net461));
 LOGIC0_X1 _3720__462 (.Z(net462));
 LOGIC0_X1 _3721__463 (.Z(net463));
 LOGIC0_X1 _3722__464 (.Z(net464));
 LOGIC0_X1 _3723__465 (.Z(net465));
 LOGIC0_X1 _3724__466 (.Z(net466));
 LOGIC0_X1 _3725__467 (.Z(net467));
 LOGIC0_X1 _3726__468 (.Z(net468));
 LOGIC0_X1 _3727__469 (.Z(net469));
 LOGIC0_X1 _3728__470 (.Z(net470));
 LOGIC0_X1 _3729__471 (.Z(net471));
 LOGIC0_X1 _3730__472 (.Z(net472));
 LOGIC0_X1 _3731__473 (.Z(net473));
 LOGIC0_X1 _3732__474 (.Z(net474));
 LOGIC0_X1 _3733__475 (.Z(net475));
 LOGIC0_X1 _3734__476 (.Z(net476));
 LOGIC0_X1 _3735__477 (.Z(net477));
 LOGIC0_X1 _3736__478 (.Z(net478));
 LOGIC0_X1 _3737__479 (.Z(net479));
 LOGIC0_X1 _3738__480 (.Z(net480));
 LOGIC0_X1 _3739__481 (.Z(net481));
 LOGIC0_X1 _3740__482 (.Z(net482));
 LOGIC0_X1 _3741__483 (.Z(net483));
 LOGIC0_X1 _3742__484 (.Z(net484));
 LOGIC0_X1 _3743__485 (.Z(net485));
 LOGIC0_X1 _3744__486 (.Z(net486));
 LOGIC0_X1 _3745__487 (.Z(net487));
 LOGIC0_X1 _3746__488 (.Z(net488));
 LOGIC0_X1 _3747__489 (.Z(net489));
 LOGIC0_X1 _3748__490 (.Z(net490));
 LOGIC0_X1 _3749__491 (.Z(net491));
 LOGIC0_X1 _3750__492 (.Z(net492));
 LOGIC0_X1 _3751__493 (.Z(net493));
 LOGIC0_X1 _3752__494 (.Z(net494));
 LOGIC0_X1 _3753__495 (.Z(net495));
 LOGIC0_X1 _3754__496 (.Z(net496));
 LOGIC0_X1 _3755__497 (.Z(net497));
 LOGIC0_X1 _3756__498 (.Z(net498));
 LOGIC0_X1 _3757__499 (.Z(net499));
 LOGIC0_X1 _3758__500 (.Z(net500));
 LOGIC0_X1 _3759__501 (.Z(net501));
 LOGIC0_X1 _3760__502 (.Z(net502));
 LOGIC0_X1 _3761__503 (.Z(net503));
 LOGIC0_X1 _3762__504 (.Z(net504));
 LOGIC0_X1 _3763__505 (.Z(net505));
 LOGIC0_X1 _3764__506 (.Z(net506));
 LOGIC0_X1 _3765__507 (.Z(net507));
 LOGIC0_X1 _3766__508 (.Z(net508));
 LOGIC0_X1 _3767__509 (.Z(net509));
 LOGIC0_X1 _3768__510 (.Z(net510));
 LOGIC0_X1 _3769__511 (.Z(net511));
 LOGIC0_X1 _3770__512 (.Z(net512));
 LOGIC0_X1 _3771__513 (.Z(net513));
 LOGIC0_X1 _3772__514 (.Z(net514));
 LOGIC0_X1 _3773__515 (.Z(net515));
 LOGIC0_X1 _3774__516 (.Z(net516));
 LOGIC0_X1 _3775__517 (.Z(net517));
 LOGIC0_X1 _3776__518 (.Z(net518));
 LOGIC0_X1 _3777__519 (.Z(net519));
 LOGIC0_X1 _3778__520 (.Z(net520));
 LOGIC0_X1 _3779__521 (.Z(net521));
 LOGIC0_X1 _3780__522 (.Z(net522));
 LOGIC0_X1 _3781__523 (.Z(net523));
 LOGIC0_X1 _3782__524 (.Z(net524));
 LOGIC0_X1 _3783__525 (.Z(net525));
 LOGIC0_X1 _3784__526 (.Z(net526));
 LOGIC0_X1 _3785__527 (.Z(net527));
 LOGIC0_X1 _3786__528 (.Z(net528));
 LOGIC0_X1 _3787__529 (.Z(net529));
 LOGIC0_X1 _3788__530 (.Z(net530));
 LOGIC0_X1 _3789__531 (.Z(net531));
 LOGIC0_X1 _3790__532 (.Z(net532));
 LOGIC0_X1 _3791__533 (.Z(net533));
 LOGIC0_X1 _3792__534 (.Z(net534));
 LOGIC0_X1 _3793__535 (.Z(net535));
 LOGIC0_X1 _3794__536 (.Z(net536));
 LOGIC0_X1 _3795__537 (.Z(net537));
 LOGIC0_X1 _3796__538 (.Z(net538));
 LOGIC0_X1 _3797__539 (.Z(net539));
 LOGIC0_X1 _3798__540 (.Z(net540));
 LOGIC0_X1 _3799__541 (.Z(net541));
 LOGIC0_X1 _3800__542 (.Z(net542));
 LOGIC0_X1 _3801__543 (.Z(net543));
 LOGIC0_X1 _3802__544 (.Z(net544));
 LOGIC0_X1 _3803__545 (.Z(net545));
 LOGIC0_X1 _3804__546 (.Z(net546));
 LOGIC0_X1 _3805__547 (.Z(net547));
 LOGIC0_X1 _3806__548 (.Z(net548));
 LOGIC0_X1 _3807__549 (.Z(net549));
 LOGIC0_X1 _3808__550 (.Z(net550));
 LOGIC0_X1 _3809__551 (.Z(net551));
 LOGIC0_X1 _3810__552 (.Z(net552));
 LOGIC0_X1 _3811__553 (.Z(net553));
 LOGIC0_X1 _3812__554 (.Z(net554));
 LOGIC0_X1 _3813__555 (.Z(net555));
 LOGIC0_X1 _3814__556 (.Z(net556));
 LOGIC0_X1 _3815__557 (.Z(net557));
 LOGIC0_X1 _3816__558 (.Z(net558));
 LOGIC0_X1 _3817__559 (.Z(net559));
 LOGIC0_X1 _3818__560 (.Z(net560));
 LOGIC0_X1 _3819__561 (.Z(net561));
 LOGIC0_X1 _3820__562 (.Z(net562));
 LOGIC0_X1 _3821__563 (.Z(net563));
 LOGIC0_X1 _3822__564 (.Z(net564));
 LOGIC0_X1 _3823__565 (.Z(net565));
 LOGIC0_X1 _3824__566 (.Z(net566));
 LOGIC0_X1 _3825__567 (.Z(net567));
 LOGIC0_X1 _3826__568 (.Z(net568));
 LOGIC0_X1 _3827__569 (.Z(net569));
 LOGIC0_X1 _3828__570 (.Z(net570));
 LOGIC0_X1 _3829__571 (.Z(net571));
 LOGIC0_X1 _3830__572 (.Z(net572));
 LOGIC0_X1 _3831__573 (.Z(net573));
 LOGIC0_X1 _3832__574 (.Z(net574));
 LOGIC0_X1 _3833__575 (.Z(net575));
 LOGIC0_X1 _3834__576 (.Z(net576));
 LOGIC0_X1 _3835__577 (.Z(net577));
 LOGIC0_X1 _3836__578 (.Z(net578));
 LOGIC0_X1 _3837__579 (.Z(net579));
 LOGIC0_X1 _3838__580 (.Z(net580));
 LOGIC0_X1 _3839__581 (.Z(net581));
 LOGIC0_X1 _3840__582 (.Z(net582));
 LOGIC0_X1 _3841__583 (.Z(net583));
 LOGIC0_X1 _3842__584 (.Z(net584));
 LOGIC0_X1 _3843__585 (.Z(net585));
 LOGIC0_X1 _3844__586 (.Z(net586));
 LOGIC0_X1 _3845__587 (.Z(net587));
 LOGIC0_X1 _3846__588 (.Z(net588));
 LOGIC0_X1 _3847__589 (.Z(net589));
 LOGIC0_X1 _3848__590 (.Z(net590));
 LOGIC0_X1 _3849__591 (.Z(net591));
 LOGIC0_X1 _3850__592 (.Z(net592));
 LOGIC0_X1 _3851__593 (.Z(net593));
 LOGIC0_X1 _3852__594 (.Z(net594));
 LOGIC0_X1 _3853__595 (.Z(net595));
 LOGIC0_X1 _3854__596 (.Z(net596));
 LOGIC0_X1 _3855__597 (.Z(net597));
 LOGIC0_X1 _3856__598 (.Z(net598));
 LOGIC0_X1 _3857__599 (.Z(net599));
 LOGIC0_X1 _3858__600 (.Z(net600));
 LOGIC0_X1 _3859__601 (.Z(net601));
 LOGIC0_X1 _3860__602 (.Z(net602));
 LOGIC0_X1 _3861__603 (.Z(net603));
 LOGIC0_X1 _3862__604 (.Z(net604));
 LOGIC0_X1 _3863__605 (.Z(net605));
 LOGIC0_X1 _3864__606 (.Z(net606));
 LOGIC0_X1 _3865__607 (.Z(net607));
 LOGIC0_X1 _3866__608 (.Z(net608));
 LOGIC0_X1 _3867__609 (.Z(net609));
 LOGIC0_X1 _3868__610 (.Z(net610));
 LOGIC0_X1 _3869__611 (.Z(net611));
 LOGIC0_X1 _3870__612 (.Z(net612));
 LOGIC0_X1 _3871__613 (.Z(net613));
 LOGIC0_X1 _3872__614 (.Z(net614));
 LOGIC0_X1 _3873__615 (.Z(net615));
 LOGIC0_X1 _3874__616 (.Z(net616));
 LOGIC0_X1 _3875__617 (.Z(net617));
 LOGIC0_X1 _3876__618 (.Z(net618));
 LOGIC0_X1 _3877__619 (.Z(net619));
 LOGIC0_X1 _3878__620 (.Z(net620));
 LOGIC0_X1 _3879__621 (.Z(net621));
 LOGIC0_X1 _3880__622 (.Z(net622));
 LOGIC0_X1 _3881__623 (.Z(net623));
 LOGIC0_X1 _3882__624 (.Z(net624));
 LOGIC0_X1 _3883__625 (.Z(net625));
 LOGIC0_X1 _3884__626 (.Z(net626));
 LOGIC0_X1 _3885__627 (.Z(net627));
 LOGIC0_X1 _3886__628 (.Z(net628));
 LOGIC0_X1 _3887__629 (.Z(net629));
 LOGIC0_X1 _3888__630 (.Z(net630));
 LOGIC0_X1 _3889__631 (.Z(net631));
 LOGIC0_X1 _3890__632 (.Z(net632));
 LOGIC0_X1 _3891__633 (.Z(net633));
 LOGIC0_X1 _3892__634 (.Z(net634));
 LOGIC0_X1 _3893__635 (.Z(net635));
 LOGIC0_X1 _3894__636 (.Z(net636));
 LOGIC0_X1 _3895__637 (.Z(net637));
 LOGIC0_X1 _3896__638 (.Z(net638));
 LOGIC0_X1 _3897__639 (.Z(net639));
 LOGIC0_X1 _3898__640 (.Z(net640));
 LOGIC0_X1 _3899__641 (.Z(net641));
 LOGIC0_X1 _3900__642 (.Z(net642));
 LOGIC0_X1 _3901__643 (.Z(net643));
 LOGIC0_X1 _3902__644 (.Z(net644));
 LOGIC0_X1 _3903__645 (.Z(net645));
 LOGIC0_X1 _3904__646 (.Z(net646));
 LOGIC0_X1 _3905__647 (.Z(net647));
 LOGIC0_X1 _3906__648 (.Z(net648));
 LOGIC0_X1 _3907__649 (.Z(net649));
 LOGIC0_X1 _3908__650 (.Z(net650));
 LOGIC0_X1 _3909__651 (.Z(net651));
 LOGIC0_X1 _3910__652 (.Z(net652));
 LOGIC0_X1 _3911__653 (.Z(net653));
 LOGIC0_X1 _3912__654 (.Z(net654));
 LOGIC0_X1 _3913__655 (.Z(net655));
 LOGIC0_X1 _3914__656 (.Z(net656));
 LOGIC0_X1 _3915__657 (.Z(net657));
 LOGIC0_X1 _3916__658 (.Z(net658));
 LOGIC0_X1 _3917__659 (.Z(net659));
 LOGIC0_X1 _3918__660 (.Z(net660));
 LOGIC0_X1 _3919__661 (.Z(net661));
 LOGIC0_X1 _3920__662 (.Z(net662));
 LOGIC0_X1 _3921__663 (.Z(net663));
 LOGIC0_X1 _3922__664 (.Z(net664));
 LOGIC0_X1 _3923__665 (.Z(net665));
 LOGIC0_X1 _3924__666 (.Z(net666));
 LOGIC0_X1 _3925__667 (.Z(net667));
 LOGIC0_X1 _3926__668 (.Z(net668));
 LOGIC0_X1 _3927__669 (.Z(net669));
 LOGIC0_X1 _3928__670 (.Z(net670));
 LOGIC0_X1 _3929__671 (.Z(net671));
 LOGIC0_X1 _3930__672 (.Z(net672));
 LOGIC0_X1 _3931__673 (.Z(net673));
 LOGIC0_X1 _3932__674 (.Z(net674));
 LOGIC0_X1 _3933__675 (.Z(net675));
 LOGIC0_X1 _3934__676 (.Z(net676));
 LOGIC0_X1 _3935__677 (.Z(net677));
 LOGIC0_X1 _3936__678 (.Z(net678));
 LOGIC0_X1 _3937__679 (.Z(net679));
 LOGIC0_X1 _3938__680 (.Z(net680));
 LOGIC0_X1 _3939__681 (.Z(net681));
 LOGIC0_X1 _3940__682 (.Z(net682));
 LOGIC0_X1 _3941__683 (.Z(net683));
 LOGIC0_X1 _3942__684 (.Z(net684));
 LOGIC0_X1 _3943__685 (.Z(net685));
 LOGIC0_X1 _3944__686 (.Z(net686));
 LOGIC0_X1 _3945__687 (.Z(net687));
 LOGIC0_X1 _3946__688 (.Z(net688));
 LOGIC0_X1 _3947__689 (.Z(net689));
 LOGIC0_X1 _3948__690 (.Z(net690));
 LOGIC0_X1 _3949__691 (.Z(net691));
 LOGIC0_X1 _3950__692 (.Z(net692));
 LOGIC0_X1 _3951__693 (.Z(net693));
 LOGIC0_X1 _3952__694 (.Z(net694));
 LOGIC0_X1 _3953__695 (.Z(net695));
 LOGIC0_X1 _3954__696 (.Z(net696));
 LOGIC0_X1 _3955__697 (.Z(net697));
 LOGIC0_X1 _3956__698 (.Z(net698));
 LOGIC0_X1 _3957__699 (.Z(net699));
 LOGIC0_X1 _3958__700 (.Z(net700));
 LOGIC0_X1 _3959__701 (.Z(net701));
 LOGIC0_X1 _3960__702 (.Z(net702));
 LOGIC0_X1 _3961__703 (.Z(net703));
 LOGIC0_X1 _3962__704 (.Z(net704));
 LOGIC0_X1 _3963__705 (.Z(net705));
 LOGIC0_X1 _3964__706 (.Z(net706));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X8 clkload0 (.A(clknet_4_0_0_clk));
 INV_X8 clkload1 (.A(clknet_4_1_0_clk));
 INV_X8 clkload2 (.A(clknet_4_2_0_clk));
 INV_X4 clkload3 (.A(clknet_4_3_0_clk));
 INV_X8 clkload4 (.A(clknet_4_4_0_clk));
 INV_X4 clkload5 (.A(clknet_4_5_0_clk));
 INV_X4 clkload6 (.A(clknet_4_6_0_clk));
 INV_X8 clkload7 (.A(clknet_4_8_0_clk));
 INV_X8 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_10_0_clk));
 INV_X8 clkload10 (.A(clknet_4_11_0_clk));
 INV_X8 clkload11 (.A(clknet_4_12_0_clk));
 INV_X8 clkload12 (.A(clknet_4_13_0_clk));
 INV_X8 clkload13 (.A(clknet_4_14_0_clk));
 INV_X4 clkload14 (.A(clknet_4_15_0_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X16 FILLER_0_632 ();
 FILLCELL_X8 FILLER_0_648 ();
 FILLCELL_X4 FILLER_0_656 ();
 FILLCELL_X4 FILLER_0_664 ();
 FILLCELL_X2 FILLER_0_668 ();
 FILLCELL_X1 FILLER_0_682 ();
 FILLCELL_X1 FILLER_0_687 ();
 FILLCELL_X4 FILLER_0_691 ();
 FILLCELL_X2 FILLER_0_695 ();
 FILLCELL_X8 FILLER_0_701 ();
 FILLCELL_X1 FILLER_0_716 ();
 FILLCELL_X1 FILLER_0_720 ();
 FILLCELL_X1 FILLER_0_728 ();
 FILLCELL_X4 FILLER_0_733 ();
 FILLCELL_X32 FILLER_0_740 ();
 FILLCELL_X16 FILLER_0_772 ();
 FILLCELL_X4 FILLER_0_788 ();
 FILLCELL_X1 FILLER_0_792 ();
 FILLCELL_X1 FILLER_0_797 ();
 FILLCELL_X1 FILLER_0_802 ();
 FILLCELL_X1 FILLER_0_815 ();
 FILLCELL_X1 FILLER_0_820 ();
 FILLCELL_X2 FILLER_0_824 ();
 FILLCELL_X2 FILLER_0_838 ();
 FILLCELL_X1 FILLER_0_843 ();
 FILLCELL_X1 FILLER_0_868 ();
 FILLCELL_X1 FILLER_0_878 ();
 FILLCELL_X2 FILLER_0_894 ();
 FILLCELL_X2 FILLER_0_947 ();
 FILLCELL_X1 FILLER_0_1024 ();
 FILLCELL_X1 FILLER_0_1028 ();
 FILLCELL_X1 FILLER_0_1032 ();
 FILLCELL_X1 FILLER_0_1036 ();
 FILLCELL_X1 FILLER_0_1040 ();
 FILLCELL_X1 FILLER_0_1044 ();
 FILLCELL_X1 FILLER_0_1051 ();
 FILLCELL_X1 FILLER_0_1055 ();
 FILLCELL_X1 FILLER_0_1071 ();
 FILLCELL_X1 FILLER_0_1075 ();
 FILLCELL_X1 FILLER_0_1082 ();
 FILLCELL_X1 FILLER_0_1089 ();
 FILLCELL_X1 FILLER_0_1096 ();
 FILLCELL_X2 FILLER_0_1103 ();
 FILLCELL_X2 FILLER_0_1108 ();
 FILLCELL_X2 FILLER_0_1116 ();
 FILLCELL_X1 FILLER_0_1118 ();
 FILLCELL_X1 FILLER_0_1134 ();
 FILLCELL_X16 FILLER_0_1150 ();
 FILLCELL_X4 FILLER_0_1166 ();
 FILLCELL_X2 FILLER_0_1170 ();
 FILLCELL_X2 FILLER_0_1181 ();
 FILLCELL_X2 FILLER_0_1192 ();
 FILLCELL_X1 FILLER_0_1194 ();
 FILLCELL_X2 FILLER_0_1216 ();
 FILLCELL_X2 FILLER_0_1227 ();
 FILLCELL_X2 FILLER_0_1259 ();
 FILLCELL_X1 FILLER_0_1261 ();
 FILLCELL_X1 FILLER_0_1278 ();
 FILLCELL_X1 FILLER_0_1282 ();
 FILLCELL_X1 FILLER_0_1289 ();
 FILLCELL_X2 FILLER_0_1293 ();
 FILLCELL_X1 FILLER_0_1304 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X16 FILLER_1_673 ();
 FILLCELL_X1 FILLER_1_689 ();
 FILLCELL_X16 FILLER_1_693 ();
 FILLCELL_X2 FILLER_1_709 ();
 FILLCELL_X8 FILLER_1_715 ();
 FILLCELL_X32 FILLER_1_727 ();
 FILLCELL_X32 FILLER_1_759 ();
 FILLCELL_X8 FILLER_1_791 ();
 FILLCELL_X4 FILLER_1_799 ();
 FILLCELL_X2 FILLER_1_803 ();
 FILLCELL_X4 FILLER_1_809 ();
 FILLCELL_X1 FILLER_1_818 ();
 FILLCELL_X4 FILLER_1_825 ();
 FILLCELL_X1 FILLER_1_831 ();
 FILLCELL_X4 FILLER_1_841 ();
 FILLCELL_X1 FILLER_1_845 ();
 FILLCELL_X2 FILLER_1_850 ();
 FILLCELL_X1 FILLER_1_852 ();
 FILLCELL_X1 FILLER_1_855 ();
 FILLCELL_X1 FILLER_1_858 ();
 FILLCELL_X2 FILLER_1_863 ();
 FILLCELL_X4 FILLER_1_867 ();
 FILLCELL_X2 FILLER_1_873 ();
 FILLCELL_X2 FILLER_1_877 ();
 FILLCELL_X2 FILLER_1_881 ();
 FILLCELL_X1 FILLER_1_887 ();
 FILLCELL_X1 FILLER_1_895 ();
 FILLCELL_X1 FILLER_1_898 ();
 FILLCELL_X1 FILLER_1_901 ();
 FILLCELL_X1 FILLER_1_904 ();
 FILLCELL_X1 FILLER_1_907 ();
 FILLCELL_X1 FILLER_1_910 ();
 FILLCELL_X1 FILLER_1_913 ();
 FILLCELL_X1 FILLER_1_916 ();
 FILLCELL_X1 FILLER_1_919 ();
 FILLCELL_X1 FILLER_1_922 ();
 FILLCELL_X1 FILLER_1_925 ();
 FILLCELL_X1 FILLER_1_928 ();
 FILLCELL_X1 FILLER_1_931 ();
 FILLCELL_X1 FILLER_1_934 ();
 FILLCELL_X1 FILLER_1_937 ();
 FILLCELL_X1 FILLER_1_940 ();
 FILLCELL_X1 FILLER_1_943 ();
 FILLCELL_X1 FILLER_1_946 ();
 FILLCELL_X1 FILLER_1_952 ();
 FILLCELL_X1 FILLER_1_957 ();
 FILLCELL_X2 FILLER_1_962 ();
 FILLCELL_X1 FILLER_1_966 ();
 FILLCELL_X1 FILLER_1_969 ();
 FILLCELL_X1 FILLER_1_972 ();
 FILLCELL_X1 FILLER_1_975 ();
 FILLCELL_X1 FILLER_1_978 ();
 FILLCELL_X1 FILLER_1_981 ();
 FILLCELL_X1 FILLER_1_984 ();
 FILLCELL_X2 FILLER_1_989 ();
 FILLCELL_X1 FILLER_1_993 ();
 FILLCELL_X1 FILLER_1_996 ();
 FILLCELL_X1 FILLER_1_999 ();
 FILLCELL_X1 FILLER_1_1002 ();
 FILLCELL_X1 FILLER_1_1005 ();
 FILLCELL_X1 FILLER_1_1008 ();
 FILLCELL_X1 FILLER_1_1011 ();
 FILLCELL_X1 FILLER_1_1014 ();
 FILLCELL_X1 FILLER_1_1017 ();
 FILLCELL_X1 FILLER_1_1020 ();
 FILLCELL_X1 FILLER_1_1032 ();
 FILLCELL_X2 FILLER_1_1035 ();
 FILLCELL_X2 FILLER_1_1039 ();
 FILLCELL_X2 FILLER_1_1043 ();
 FILLCELL_X1 FILLER_1_1045 ();
 FILLCELL_X2 FILLER_1_1059 ();
 FILLCELL_X1 FILLER_1_1061 ();
 FILLCELL_X1 FILLER_1_1064 ();
 FILLCELL_X1 FILLER_1_1067 ();
 FILLCELL_X2 FILLER_1_1070 ();
 FILLCELL_X1 FILLER_1_1074 ();
 FILLCELL_X2 FILLER_1_1088 ();
 FILLCELL_X1 FILLER_1_1092 ();
 FILLCELL_X2 FILLER_1_1095 ();
 FILLCELL_X2 FILLER_1_1099 ();
 FILLCELL_X2 FILLER_1_1103 ();
 FILLCELL_X1 FILLER_1_1107 ();
 FILLCELL_X1 FILLER_1_1110 ();
 FILLCELL_X2 FILLER_1_1118 ();
 FILLCELL_X1 FILLER_1_1126 ();
 FILLCELL_X1 FILLER_1_1134 ();
 FILLCELL_X1 FILLER_1_1137 ();
 FILLCELL_X1 FILLER_1_1140 ();
 FILLCELL_X1 FILLER_1_1143 ();
 FILLCELL_X1 FILLER_1_1146 ();
 FILLCELL_X16 FILLER_1_1149 ();
 FILLCELL_X4 FILLER_1_1165 ();
 FILLCELL_X2 FILLER_1_1169 ();
 FILLCELL_X1 FILLER_1_1171 ();
 FILLCELL_X1 FILLER_1_1174 ();
 FILLCELL_X1 FILLER_1_1177 ();
 FILLCELL_X2 FILLER_1_1180 ();
 FILLCELL_X1 FILLER_1_1182 ();
 FILLCELL_X1 FILLER_1_1189 ();
 FILLCELL_X1 FILLER_1_1197 ();
 FILLCELL_X2 FILLER_1_1200 ();
 FILLCELL_X1 FILLER_1_1202 ();
 FILLCELL_X1 FILLER_1_1213 ();
 FILLCELL_X1 FILLER_1_1223 ();
 FILLCELL_X1 FILLER_1_1231 ();
 FILLCELL_X1 FILLER_1_1234 ();
 FILLCELL_X1 FILLER_1_1237 ();
 FILLCELL_X1 FILLER_1_1240 ();
 FILLCELL_X1 FILLER_1_1243 ();
 FILLCELL_X1 FILLER_1_1246 ();
 FILLCELL_X1 FILLER_1_1249 ();
 FILLCELL_X1 FILLER_1_1252 ();
 FILLCELL_X1 FILLER_1_1255 ();
 FILLCELL_X4 FILLER_1_1258 ();
 FILLCELL_X1 FILLER_1_1262 ();
 FILLCELL_X1 FILLER_1_1266 ();
 FILLCELL_X1 FILLER_1_1271 ();
 FILLCELL_X2 FILLER_1_1274 ();
 FILLCELL_X1 FILLER_1_1278 ();
 FILLCELL_X2 FILLER_1_1281 ();
 FILLCELL_X1 FILLER_1_1283 ();
 FILLCELL_X1 FILLER_1_1288 ();
 FILLCELL_X1 FILLER_1_1294 ();
 FILLCELL_X1 FILLER_1_1297 ();
 FILLCELL_X2 FILLER_1_1302 ();
 FILLCELL_X1 FILLER_1_1304 ();
 FILLCELL_X1 FILLER_1_1307 ();
 FILLCELL_X2 FILLER_1_1310 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X2 FILLER_2_824 ();
 FILLCELL_X1 FILLER_2_826 ();
 FILLCELL_X8 FILLER_2_829 ();
 FILLCELL_X2 FILLER_2_837 ();
 FILLCELL_X1 FILLER_2_839 ();
 FILLCELL_X8 FILLER_2_842 ();
 FILLCELL_X2 FILLER_2_850 ();
 FILLCELL_X1 FILLER_2_852 ();
 FILLCELL_X16 FILLER_2_855 ();
 FILLCELL_X4 FILLER_2_873 ();
 FILLCELL_X8 FILLER_2_882 ();
 FILLCELL_X2 FILLER_2_890 ();
 FILLCELL_X32 FILLER_2_894 ();
 FILLCELL_X16 FILLER_2_926 ();
 FILLCELL_X4 FILLER_2_942 ();
 FILLCELL_X2 FILLER_2_946 ();
 FILLCELL_X32 FILLER_2_950 ();
 FILLCELL_X32 FILLER_2_982 ();
 FILLCELL_X16 FILLER_2_1014 ();
 FILLCELL_X1 FILLER_2_1030 ();
 FILLCELL_X16 FILLER_2_1036 ();
 FILLCELL_X8 FILLER_2_1052 ();
 FILLCELL_X16 FILLER_2_1062 ();
 FILLCELL_X8 FILLER_2_1078 ();
 FILLCELL_X1 FILLER_2_1086 ();
 FILLCELL_X8 FILLER_2_1092 ();
 FILLCELL_X4 FILLER_2_1100 ();
 FILLCELL_X2 FILLER_2_1104 ();
 FILLCELL_X1 FILLER_2_1109 ();
 FILLCELL_X16 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1130 ();
 FILLCELL_X32 FILLER_2_1162 ();
 FILLCELL_X32 FILLER_2_1194 ();
 FILLCELL_X32 FILLER_2_1228 ();
 FILLCELL_X2 FILLER_2_1260 ();
 FILLCELL_X16 FILLER_2_1272 ();
 FILLCELL_X4 FILLER_2_1288 ();
 FILLCELL_X1 FILLER_2_1304 ();
 FILLCELL_X1 FILLER_2_1307 ();
 FILLCELL_X1 FILLER_2_1311 ();
 FILLCELL_X1 FILLER_2_1324 ();
 FILLCELL_X1 FILLER_2_1327 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X8 FILLER_3_1296 ();
 FILLCELL_X1 FILLER_3_1304 ();
 FILLCELL_X2 FILLER_3_1307 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X2 FILLER_4_1304 ();
 FILLCELL_X1 FILLER_4_1306 ();
 FILLCELL_X1 FILLER_4_1314 ();
 FILLCELL_X1 FILLER_4_1318 ();
 FILLCELL_X2 FILLER_4_1326 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X16 FILLER_5_1296 ();
 FILLCELL_X1 FILLER_5_1327 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X4 FILLER_6_1304 ();
 FILLCELL_X2 FILLER_6_1308 ();
 FILLCELL_X1 FILLER_6_1310 ();
 FILLCELL_X2 FILLER_6_1326 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X16 FILLER_7_1296 ();
 FILLCELL_X4 FILLER_7_1312 ();
 FILLCELL_X2 FILLER_7_1316 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X8 FILLER_8_1304 ();
 FILLCELL_X2 FILLER_8_1312 ();
 FILLCELL_X1 FILLER_8_1327 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X16 FILLER_9_1296 ();
 FILLCELL_X2 FILLER_9_1312 ();
 FILLCELL_X1 FILLER_9_1314 ();
 FILLCELL_X1 FILLER_9_1325 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X4 FILLER_10_1304 ();
 FILLCELL_X1 FILLER_10_1308 ();
 FILLCELL_X2 FILLER_10_1316 ();
 FILLCELL_X1 FILLER_10_1318 ();
 FILLCELL_X1 FILLER_10_1322 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X16 FILLER_11_1296 ();
 FILLCELL_X1 FILLER_11_1314 ();
 FILLCELL_X1 FILLER_11_1321 ();
 FILLCELL_X1 FILLER_11_1327 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X4 FILLER_12_1304 ();
 FILLCELL_X2 FILLER_12_1308 ();
 FILLCELL_X1 FILLER_12_1310 ();
 FILLCELL_X1 FILLER_12_1313 ();
 FILLCELL_X1 FILLER_12_1317 ();
 FILLCELL_X1 FILLER_12_1320 ();
 FILLCELL_X1 FILLER_12_1323 ();
 FILLCELL_X1 FILLER_12_1327 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X8 FILLER_13_1296 ();
 FILLCELL_X4 FILLER_13_1304 ();
 FILLCELL_X2 FILLER_13_1308 ();
 FILLCELL_X1 FILLER_13_1310 ();
 FILLCELL_X1 FILLER_13_1316 ();
 FILLCELL_X1 FILLER_13_1327 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X8 FILLER_14_1304 ();
 FILLCELL_X4 FILLER_14_1312 ();
 FILLCELL_X2 FILLER_14_1321 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X8 FILLER_15_1296 ();
 FILLCELL_X4 FILLER_15_1304 ();
 FILLCELL_X2 FILLER_15_1308 ();
 FILLCELL_X1 FILLER_15_1310 ();
 FILLCELL_X1 FILLER_15_1316 ();
 FILLCELL_X1 FILLER_15_1327 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X8 FILLER_16_1304 ();
 FILLCELL_X2 FILLER_16_1312 ();
 FILLCELL_X2 FILLER_16_1319 ();
 FILLCELL_X1 FILLER_16_1323 ();
 FILLCELL_X1 FILLER_16_1327 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X16 FILLER_17_1296 ();
 FILLCELL_X2 FILLER_17_1312 ();
 FILLCELL_X1 FILLER_17_1321 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X8 FILLER_18_1304 ();
 FILLCELL_X4 FILLER_18_1312 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X8 FILLER_19_1296 ();
 FILLCELL_X4 FILLER_19_1304 ();
 FILLCELL_X2 FILLER_19_1308 ();
 FILLCELL_X1 FILLER_19_1310 ();
 FILLCELL_X1 FILLER_19_1316 ();
 FILLCELL_X1 FILLER_19_1324 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X8 FILLER_20_1304 ();
 FILLCELL_X4 FILLER_20_1312 ();
 FILLCELL_X2 FILLER_20_1321 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X16 FILLER_21_1296 ();
 FILLCELL_X2 FILLER_21_1312 ();
 FILLCELL_X4 FILLER_21_1316 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X4 FILLER_22_1304 ();
 FILLCELL_X2 FILLER_22_1308 ();
 FILLCELL_X1 FILLER_22_1310 ();
 FILLCELL_X2 FILLER_22_1321 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X8 FILLER_23_1296 ();
 FILLCELL_X4 FILLER_23_1304 ();
 FILLCELL_X2 FILLER_23_1308 ();
 FILLCELL_X1 FILLER_23_1310 ();
 FILLCELL_X1 FILLER_23_1316 ();
 FILLCELL_X1 FILLER_23_1327 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X8 FILLER_24_1304 ();
 FILLCELL_X2 FILLER_24_1312 ();
 FILLCELL_X2 FILLER_24_1319 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X16 FILLER_25_1296 ();
 FILLCELL_X1 FILLER_25_1312 ();
 FILLCELL_X1 FILLER_25_1315 ();
 FILLCELL_X1 FILLER_25_1324 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X8 FILLER_26_1304 ();
 FILLCELL_X4 FILLER_26_1312 ();
 FILLCELL_X1 FILLER_26_1323 ();
 FILLCELL_X1 FILLER_26_1327 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X8 FILLER_27_1296 ();
 FILLCELL_X4 FILLER_27_1304 ();
 FILLCELL_X2 FILLER_27_1308 ();
 FILLCELL_X1 FILLER_27_1310 ();
 FILLCELL_X1 FILLER_27_1316 ();
 FILLCELL_X1 FILLER_27_1327 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X8 FILLER_28_1304 ();
 FILLCELL_X4 FILLER_28_1312 ();
 FILLCELL_X1 FILLER_28_1316 ();
 FILLCELL_X1 FILLER_28_1319 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X16 FILLER_29_1296 ();
 FILLCELL_X2 FILLER_29_1312 ();
 FILLCELL_X1 FILLER_29_1321 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X8 FILLER_30_1304 ();
 FILLCELL_X2 FILLER_30_1312 ();
 FILLCELL_X2 FILLER_30_1324 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X16 FILLER_31_1296 ();
 FILLCELL_X2 FILLER_31_1312 ();
 FILLCELL_X1 FILLER_31_1314 ();
 FILLCELL_X2 FILLER_31_1320 ();
 FILLCELL_X1 FILLER_31_1322 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X4 FILLER_32_1304 ();
 FILLCELL_X2 FILLER_32_1308 ();
 FILLCELL_X1 FILLER_32_1310 ();
 FILLCELL_X2 FILLER_32_1326 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X16 FILLER_33_1296 ();
 FILLCELL_X1 FILLER_33_1319 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X4 FILLER_34_1304 ();
 FILLCELL_X2 FILLER_34_1308 ();
 FILLCELL_X1 FILLER_34_1310 ();
 FILLCELL_X4 FILLER_34_1316 ();
 FILLCELL_X1 FILLER_34_1320 ();
 FILLCELL_X1 FILLER_34_1323 ();
 FILLCELL_X1 FILLER_34_1327 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X8 FILLER_35_1296 ();
 FILLCELL_X4 FILLER_35_1304 ();
 FILLCELL_X2 FILLER_35_1308 ();
 FILLCELL_X1 FILLER_35_1310 ();
 FILLCELL_X1 FILLER_35_1316 ();
 FILLCELL_X1 FILLER_35_1327 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X8 FILLER_36_1304 ();
 FILLCELL_X2 FILLER_36_1312 ();
 FILLCELL_X1 FILLER_36_1316 ();
 FILLCELL_X1 FILLER_36_1324 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X16 FILLER_37_1296 ();
 FILLCELL_X4 FILLER_37_1312 ();
 FILLCELL_X1 FILLER_37_1316 ();
 FILLCELL_X1 FILLER_37_1320 ();
 FILLCELL_X1 FILLER_37_1323 ();
 FILLCELL_X1 FILLER_37_1327 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X4 FILLER_38_1304 ();
 FILLCELL_X2 FILLER_38_1308 ();
 FILLCELL_X1 FILLER_38_1310 ();
 FILLCELL_X1 FILLER_38_1313 ();
 FILLCELL_X1 FILLER_38_1317 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X8 FILLER_39_1296 ();
 FILLCELL_X4 FILLER_39_1304 ();
 FILLCELL_X2 FILLER_39_1308 ();
 FILLCELL_X1 FILLER_39_1310 ();
 FILLCELL_X1 FILLER_39_1316 ();
 FILLCELL_X1 FILLER_39_1327 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X4 FILLER_40_1304 ();
 FILLCELL_X2 FILLER_40_1308 ();
 FILLCELL_X1 FILLER_40_1310 ();
 FILLCELL_X1 FILLER_40_1313 ();
 FILLCELL_X1 FILLER_40_1324 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X16 FILLER_41_1296 ();
 FILLCELL_X2 FILLER_41_1312 ();
 FILLCELL_X4 FILLER_41_1316 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X8 FILLER_42_1304 ();
 FILLCELL_X4 FILLER_42_1312 ();
 FILLCELL_X1 FILLER_42_1323 ();
 FILLCELL_X1 FILLER_42_1327 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X8 FILLER_43_1296 ();
 FILLCELL_X4 FILLER_43_1304 ();
 FILLCELL_X2 FILLER_43_1308 ();
 FILLCELL_X1 FILLER_43_1310 ();
 FILLCELL_X1 FILLER_43_1316 ();
 FILLCELL_X1 FILLER_43_1327 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X8 FILLER_44_1304 ();
 FILLCELL_X2 FILLER_44_1312 ();
 FILLCELL_X1 FILLER_44_1316 ();
 FILLCELL_X1 FILLER_44_1320 ();
 FILLCELL_X2 FILLER_44_1326 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X8 FILLER_45_1296 ();
 FILLCELL_X4 FILLER_45_1304 ();
 FILLCELL_X2 FILLER_45_1308 ();
 FILLCELL_X1 FILLER_45_1310 ();
 FILLCELL_X1 FILLER_45_1323 ();
 FILLCELL_X1 FILLER_45_1327 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X4 FILLER_46_1304 ();
 FILLCELL_X2 FILLER_46_1308 ();
 FILLCELL_X1 FILLER_46_1310 ();
 FILLCELL_X2 FILLER_46_1316 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X8 FILLER_47_1296 ();
 FILLCELL_X4 FILLER_47_1304 ();
 FILLCELL_X2 FILLER_47_1308 ();
 FILLCELL_X1 FILLER_47_1310 ();
 FILLCELL_X4 FILLER_47_1316 ();
 FILLCELL_X2 FILLER_47_1320 ();
 FILLCELL_X1 FILLER_47_1327 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X8 FILLER_48_1304 ();
 FILLCELL_X4 FILLER_48_1312 ();
 FILLCELL_X1 FILLER_48_1318 ();
 FILLCELL_X1 FILLER_48_1327 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X8 FILLER_49_1296 ();
 FILLCELL_X4 FILLER_49_1304 ();
 FILLCELL_X2 FILLER_49_1308 ();
 FILLCELL_X1 FILLER_49_1310 ();
 FILLCELL_X1 FILLER_49_1313 ();
 FILLCELL_X1 FILLER_49_1317 ();
 FILLCELL_X1 FILLER_49_1321 ();
 FILLCELL_X1 FILLER_49_1324 ();
 FILLCELL_X32 FILLER_50_6 ();
 FILLCELL_X32 FILLER_50_38 ();
 FILLCELL_X32 FILLER_50_70 ();
 FILLCELL_X32 FILLER_50_102 ();
 FILLCELL_X32 FILLER_50_134 ();
 FILLCELL_X32 FILLER_50_166 ();
 FILLCELL_X32 FILLER_50_198 ();
 FILLCELL_X32 FILLER_50_230 ();
 FILLCELL_X32 FILLER_50_262 ();
 FILLCELL_X32 FILLER_50_294 ();
 FILLCELL_X32 FILLER_50_326 ();
 FILLCELL_X32 FILLER_50_358 ();
 FILLCELL_X32 FILLER_50_390 ();
 FILLCELL_X32 FILLER_50_422 ();
 FILLCELL_X32 FILLER_50_454 ();
 FILLCELL_X32 FILLER_50_486 ();
 FILLCELL_X32 FILLER_50_518 ();
 FILLCELL_X32 FILLER_50_550 ();
 FILLCELL_X32 FILLER_50_582 ();
 FILLCELL_X16 FILLER_50_614 ();
 FILLCELL_X1 FILLER_50_630 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X8 FILLER_50_1304 ();
 FILLCELL_X4 FILLER_50_1312 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X8 FILLER_51_705 ();
 FILLCELL_X1 FILLER_51_713 ();
 FILLCELL_X32 FILLER_51_734 ();
 FILLCELL_X32 FILLER_51_766 ();
 FILLCELL_X32 FILLER_51_798 ();
 FILLCELL_X32 FILLER_51_830 ();
 FILLCELL_X32 FILLER_51_862 ();
 FILLCELL_X32 FILLER_51_894 ();
 FILLCELL_X32 FILLER_51_926 ();
 FILLCELL_X32 FILLER_51_958 ();
 FILLCELL_X32 FILLER_51_990 ();
 FILLCELL_X32 FILLER_51_1022 ();
 FILLCELL_X32 FILLER_51_1054 ();
 FILLCELL_X32 FILLER_51_1086 ();
 FILLCELL_X32 FILLER_51_1118 ();
 FILLCELL_X32 FILLER_51_1150 ();
 FILLCELL_X32 FILLER_51_1182 ();
 FILLCELL_X32 FILLER_51_1214 ();
 FILLCELL_X16 FILLER_51_1246 ();
 FILLCELL_X1 FILLER_51_1262 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X8 FILLER_51_1296 ();
 FILLCELL_X4 FILLER_51_1304 ();
 FILLCELL_X2 FILLER_51_1308 ();
 FILLCELL_X1 FILLER_51_1310 ();
 FILLCELL_X1 FILLER_51_1318 ();
 FILLCELL_X1 FILLER_51_1327 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X16 FILLER_52_696 ();
 FILLCELL_X1 FILLER_52_716 ();
 FILLCELL_X2 FILLER_52_729 ();
 FILLCELL_X1 FILLER_52_731 ();
 FILLCELL_X32 FILLER_52_746 ();
 FILLCELL_X32 FILLER_52_778 ();
 FILLCELL_X32 FILLER_52_810 ();
 FILLCELL_X32 FILLER_52_842 ();
 FILLCELL_X32 FILLER_52_874 ();
 FILLCELL_X32 FILLER_52_906 ();
 FILLCELL_X32 FILLER_52_938 ();
 FILLCELL_X32 FILLER_52_970 ();
 FILLCELL_X32 FILLER_52_1002 ();
 FILLCELL_X32 FILLER_52_1034 ();
 FILLCELL_X32 FILLER_52_1066 ();
 FILLCELL_X32 FILLER_52_1098 ();
 FILLCELL_X32 FILLER_52_1130 ();
 FILLCELL_X32 FILLER_52_1162 ();
 FILLCELL_X32 FILLER_52_1194 ();
 FILLCELL_X32 FILLER_52_1226 ();
 FILLCELL_X32 FILLER_52_1258 ();
 FILLCELL_X16 FILLER_52_1290 ();
 FILLCELL_X8 FILLER_52_1306 ();
 FILLCELL_X2 FILLER_52_1319 ();
 FILLCELL_X2 FILLER_52_1326 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X16 FILLER_53_641 ();
 FILLCELL_X8 FILLER_53_657 ();
 FILLCELL_X4 FILLER_53_665 ();
 FILLCELL_X1 FILLER_53_669 ();
 FILLCELL_X16 FILLER_53_690 ();
 FILLCELL_X8 FILLER_53_706 ();
 FILLCELL_X32 FILLER_53_728 ();
 FILLCELL_X32 FILLER_53_760 ();
 FILLCELL_X32 FILLER_53_792 ();
 FILLCELL_X32 FILLER_53_824 ();
 FILLCELL_X32 FILLER_53_856 ();
 FILLCELL_X32 FILLER_53_888 ();
 FILLCELL_X32 FILLER_53_920 ();
 FILLCELL_X32 FILLER_53_952 ();
 FILLCELL_X32 FILLER_53_984 ();
 FILLCELL_X32 FILLER_53_1016 ();
 FILLCELL_X32 FILLER_53_1048 ();
 FILLCELL_X32 FILLER_53_1080 ();
 FILLCELL_X32 FILLER_53_1112 ();
 FILLCELL_X32 FILLER_53_1144 ();
 FILLCELL_X32 FILLER_53_1176 ();
 FILLCELL_X32 FILLER_53_1208 ();
 FILLCELL_X16 FILLER_53_1240 ();
 FILLCELL_X4 FILLER_53_1256 ();
 FILLCELL_X2 FILLER_53_1260 ();
 FILLCELL_X1 FILLER_53_1262 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X8 FILLER_53_1296 ();
 FILLCELL_X4 FILLER_53_1304 ();
 FILLCELL_X2 FILLER_53_1308 ();
 FILLCELL_X1 FILLER_53_1310 ();
 FILLCELL_X1 FILLER_53_1318 ();
 FILLCELL_X1 FILLER_53_1327 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X16 FILLER_54_632 ();
 FILLCELL_X8 FILLER_54_648 ();
 FILLCELL_X2 FILLER_54_656 ();
 FILLCELL_X1 FILLER_54_658 ();
 FILLCELL_X2 FILLER_54_677 ();
 FILLCELL_X1 FILLER_54_683 ();
 FILLCELL_X32 FILLER_54_688 ();
 FILLCELL_X32 FILLER_54_720 ();
 FILLCELL_X32 FILLER_54_752 ();
 FILLCELL_X32 FILLER_54_784 ();
 FILLCELL_X32 FILLER_54_816 ();
 FILLCELL_X32 FILLER_54_848 ();
 FILLCELL_X32 FILLER_54_880 ();
 FILLCELL_X32 FILLER_54_912 ();
 FILLCELL_X32 FILLER_54_944 ();
 FILLCELL_X32 FILLER_54_976 ();
 FILLCELL_X32 FILLER_54_1008 ();
 FILLCELL_X32 FILLER_54_1040 ();
 FILLCELL_X32 FILLER_54_1072 ();
 FILLCELL_X32 FILLER_54_1104 ();
 FILLCELL_X32 FILLER_54_1136 ();
 FILLCELL_X32 FILLER_54_1168 ();
 FILLCELL_X32 FILLER_54_1200 ();
 FILLCELL_X32 FILLER_54_1232 ();
 FILLCELL_X32 FILLER_54_1264 ();
 FILLCELL_X16 FILLER_54_1296 ();
 FILLCELL_X4 FILLER_54_1312 ();
 FILLCELL_X2 FILLER_54_1326 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X8 FILLER_55_641 ();
 FILLCELL_X2 FILLER_55_649 ();
 FILLCELL_X32 FILLER_55_685 ();
 FILLCELL_X32 FILLER_55_717 ();
 FILLCELL_X32 FILLER_55_749 ();
 FILLCELL_X32 FILLER_55_781 ();
 FILLCELL_X32 FILLER_55_813 ();
 FILLCELL_X32 FILLER_55_845 ();
 FILLCELL_X32 FILLER_55_877 ();
 FILLCELL_X32 FILLER_55_909 ();
 FILLCELL_X32 FILLER_55_941 ();
 FILLCELL_X32 FILLER_55_973 ();
 FILLCELL_X32 FILLER_55_1005 ();
 FILLCELL_X32 FILLER_55_1037 ();
 FILLCELL_X32 FILLER_55_1069 ();
 FILLCELL_X32 FILLER_55_1101 ();
 FILLCELL_X32 FILLER_55_1133 ();
 FILLCELL_X32 FILLER_55_1165 ();
 FILLCELL_X32 FILLER_55_1197 ();
 FILLCELL_X32 FILLER_55_1229 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X8 FILLER_55_1296 ();
 FILLCELL_X4 FILLER_55_1304 ();
 FILLCELL_X2 FILLER_55_1308 ();
 FILLCELL_X1 FILLER_55_1310 ();
 FILLCELL_X1 FILLER_55_1316 ();
 FILLCELL_X1 FILLER_55_1324 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X8 FILLER_56_696 ();
 FILLCELL_X4 FILLER_56_704 ();
 FILLCELL_X4 FILLER_56_722 ();
 FILLCELL_X32 FILLER_56_736 ();
 FILLCELL_X32 FILLER_56_768 ();
 FILLCELL_X32 FILLER_56_800 ();
 FILLCELL_X32 FILLER_56_832 ();
 FILLCELL_X32 FILLER_56_864 ();
 FILLCELL_X32 FILLER_56_896 ();
 FILLCELL_X32 FILLER_56_928 ();
 FILLCELL_X32 FILLER_56_960 ();
 FILLCELL_X32 FILLER_56_992 ();
 FILLCELL_X32 FILLER_56_1024 ();
 FILLCELL_X32 FILLER_56_1056 ();
 FILLCELL_X32 FILLER_56_1088 ();
 FILLCELL_X32 FILLER_56_1120 ();
 FILLCELL_X32 FILLER_56_1152 ();
 FILLCELL_X32 FILLER_56_1184 ();
 FILLCELL_X32 FILLER_56_1216 ();
 FILLCELL_X32 FILLER_56_1248 ();
 FILLCELL_X32 FILLER_56_1280 ();
 FILLCELL_X2 FILLER_56_1312 ();
 FILLCELL_X2 FILLER_56_1319 ();
 FILLCELL_X1 FILLER_56_1323 ();
 FILLCELL_X1 FILLER_56_1327 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X16 FILLER_57_641 ();
 FILLCELL_X4 FILLER_57_657 ();
 FILLCELL_X2 FILLER_57_661 ();
 FILLCELL_X1 FILLER_57_663 ();
 FILLCELL_X4 FILLER_57_691 ();
 FILLCELL_X2 FILLER_57_695 ();
 FILLCELL_X1 FILLER_57_713 ();
 FILLCELL_X32 FILLER_57_728 ();
 FILLCELL_X32 FILLER_57_760 ();
 FILLCELL_X32 FILLER_57_792 ();
 FILLCELL_X32 FILLER_57_824 ();
 FILLCELL_X32 FILLER_57_856 ();
 FILLCELL_X32 FILLER_57_888 ();
 FILLCELL_X32 FILLER_57_920 ();
 FILLCELL_X32 FILLER_57_952 ();
 FILLCELL_X32 FILLER_57_984 ();
 FILLCELL_X32 FILLER_57_1016 ();
 FILLCELL_X32 FILLER_57_1048 ();
 FILLCELL_X32 FILLER_57_1080 ();
 FILLCELL_X32 FILLER_57_1112 ();
 FILLCELL_X32 FILLER_57_1144 ();
 FILLCELL_X32 FILLER_57_1176 ();
 FILLCELL_X32 FILLER_57_1208 ();
 FILLCELL_X16 FILLER_57_1240 ();
 FILLCELL_X4 FILLER_57_1256 ();
 FILLCELL_X2 FILLER_57_1260 ();
 FILLCELL_X1 FILLER_57_1262 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X8 FILLER_57_1296 ();
 FILLCELL_X4 FILLER_57_1304 ();
 FILLCELL_X2 FILLER_57_1308 ();
 FILLCELL_X1 FILLER_57_1310 ();
 FILLCELL_X1 FILLER_57_1318 ();
 FILLCELL_X1 FILLER_57_1324 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X8 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_90 ();
 FILLCELL_X32 FILLER_58_122 ();
 FILLCELL_X32 FILLER_58_154 ();
 FILLCELL_X32 FILLER_58_186 ();
 FILLCELL_X32 FILLER_58_218 ();
 FILLCELL_X32 FILLER_58_250 ();
 FILLCELL_X32 FILLER_58_282 ();
 FILLCELL_X32 FILLER_58_314 ();
 FILLCELL_X32 FILLER_58_346 ();
 FILLCELL_X32 FILLER_58_378 ();
 FILLCELL_X32 FILLER_58_410 ();
 FILLCELL_X32 FILLER_58_442 ();
 FILLCELL_X32 FILLER_58_474 ();
 FILLCELL_X32 FILLER_58_506 ();
 FILLCELL_X32 FILLER_58_538 ();
 FILLCELL_X32 FILLER_58_570 ();
 FILLCELL_X16 FILLER_58_602 ();
 FILLCELL_X8 FILLER_58_618 ();
 FILLCELL_X4 FILLER_58_626 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X1 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_674 ();
 FILLCELL_X8 FILLER_58_706 ();
 FILLCELL_X4 FILLER_58_714 ();
 FILLCELL_X8 FILLER_58_728 ();
 FILLCELL_X4 FILLER_58_736 ();
 FILLCELL_X2 FILLER_58_740 ();
 FILLCELL_X1 FILLER_58_742 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X4 FILLER_58_1304 ();
 FILLCELL_X2 FILLER_58_1308 ();
 FILLCELL_X1 FILLER_58_1310 ();
 FILLCELL_X4 FILLER_58_1313 ();
 FILLCELL_X1 FILLER_58_1317 ();
 FILLCELL_X1 FILLER_58_1323 ();
 FILLCELL_X1 FILLER_58_1327 ();
 FILLCELL_X32 FILLER_59_6 ();
 FILLCELL_X16 FILLER_59_38 ();
 FILLCELL_X8 FILLER_59_54 ();
 FILLCELL_X1 FILLER_59_62 ();
 FILLCELL_X16 FILLER_59_83 ();
 FILLCELL_X1 FILLER_59_99 ();
 FILLCELL_X16 FILLER_59_117 ();
 FILLCELL_X4 FILLER_59_133 ();
 FILLCELL_X2 FILLER_59_137 ();
 FILLCELL_X32 FILLER_59_156 ();
 FILLCELL_X32 FILLER_59_188 ();
 FILLCELL_X32 FILLER_59_220 ();
 FILLCELL_X32 FILLER_59_252 ();
 FILLCELL_X32 FILLER_59_284 ();
 FILLCELL_X32 FILLER_59_316 ();
 FILLCELL_X32 FILLER_59_348 ();
 FILLCELL_X32 FILLER_59_380 ();
 FILLCELL_X32 FILLER_59_412 ();
 FILLCELL_X32 FILLER_59_444 ();
 FILLCELL_X32 FILLER_59_476 ();
 FILLCELL_X32 FILLER_59_508 ();
 FILLCELL_X32 FILLER_59_540 ();
 FILLCELL_X32 FILLER_59_572 ();
 FILLCELL_X16 FILLER_59_604 ();
 FILLCELL_X4 FILLER_59_620 ();
 FILLCELL_X2 FILLER_59_624 ();
 FILLCELL_X1 FILLER_59_626 ();
 FILLCELL_X32 FILLER_59_652 ();
 FILLCELL_X32 FILLER_59_684 ();
 FILLCELL_X16 FILLER_59_716 ();
 FILLCELL_X1 FILLER_59_732 ();
 FILLCELL_X4 FILLER_59_749 ();
 FILLCELL_X2 FILLER_59_753 ();
 FILLCELL_X1 FILLER_59_755 ();
 FILLCELL_X32 FILLER_59_760 ();
 FILLCELL_X32 FILLER_59_792 ();
 FILLCELL_X32 FILLER_59_824 ();
 FILLCELL_X32 FILLER_59_856 ();
 FILLCELL_X32 FILLER_59_888 ();
 FILLCELL_X32 FILLER_59_920 ();
 FILLCELL_X32 FILLER_59_952 ();
 FILLCELL_X32 FILLER_59_984 ();
 FILLCELL_X32 FILLER_59_1016 ();
 FILLCELL_X32 FILLER_59_1048 ();
 FILLCELL_X32 FILLER_59_1080 ();
 FILLCELL_X32 FILLER_59_1112 ();
 FILLCELL_X32 FILLER_59_1144 ();
 FILLCELL_X32 FILLER_59_1176 ();
 FILLCELL_X32 FILLER_59_1208 ();
 FILLCELL_X16 FILLER_59_1240 ();
 FILLCELL_X4 FILLER_59_1256 ();
 FILLCELL_X2 FILLER_59_1260 ();
 FILLCELL_X1 FILLER_59_1262 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X16 FILLER_59_1296 ();
 FILLCELL_X2 FILLER_59_1312 ();
 FILLCELL_X2 FILLER_59_1319 ();
 FILLCELL_X1 FILLER_59_1321 ();
 FILLCELL_X1 FILLER_59_1324 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X8 FILLER_60_65 ();
 FILLCELL_X4 FILLER_60_73 ();
 FILLCELL_X1 FILLER_60_77 ();
 FILLCELL_X16 FILLER_60_85 ();
 FILLCELL_X4 FILLER_60_101 ();
 FILLCELL_X1 FILLER_60_105 ();
 FILLCELL_X2 FILLER_60_113 ();
 FILLCELL_X1 FILLER_60_115 ();
 FILLCELL_X32 FILLER_60_139 ();
 FILLCELL_X32 FILLER_60_171 ();
 FILLCELL_X32 FILLER_60_203 ();
 FILLCELL_X32 FILLER_60_235 ();
 FILLCELL_X32 FILLER_60_267 ();
 FILLCELL_X32 FILLER_60_299 ();
 FILLCELL_X32 FILLER_60_331 ();
 FILLCELL_X32 FILLER_60_363 ();
 FILLCELL_X32 FILLER_60_395 ();
 FILLCELL_X32 FILLER_60_427 ();
 FILLCELL_X32 FILLER_60_459 ();
 FILLCELL_X32 FILLER_60_491 ();
 FILLCELL_X32 FILLER_60_523 ();
 FILLCELL_X32 FILLER_60_555 ();
 FILLCELL_X32 FILLER_60_587 ();
 FILLCELL_X8 FILLER_60_619 ();
 FILLCELL_X4 FILLER_60_627 ();
 FILLCELL_X8 FILLER_60_632 ();
 FILLCELL_X2 FILLER_60_640 ();
 FILLCELL_X1 FILLER_60_642 ();
 FILLCELL_X8 FILLER_60_651 ();
 FILLCELL_X4 FILLER_60_659 ();
 FILLCELL_X1 FILLER_60_663 ();
 FILLCELL_X16 FILLER_60_681 ();
 FILLCELL_X8 FILLER_60_697 ();
 FILLCELL_X1 FILLER_60_705 ();
 FILLCELL_X8 FILLER_60_710 ();
 FILLCELL_X1 FILLER_60_718 ();
 FILLCELL_X8 FILLER_60_725 ();
 FILLCELL_X4 FILLER_60_733 ();
 FILLCELL_X2 FILLER_60_737 ();
 FILLCELL_X1 FILLER_60_739 ();
 FILLCELL_X1 FILLER_60_750 ();
 FILLCELL_X32 FILLER_60_777 ();
 FILLCELL_X32 FILLER_60_809 ();
 FILLCELL_X32 FILLER_60_841 ();
 FILLCELL_X32 FILLER_60_873 ();
 FILLCELL_X32 FILLER_60_905 ();
 FILLCELL_X32 FILLER_60_937 ();
 FILLCELL_X32 FILLER_60_969 ();
 FILLCELL_X32 FILLER_60_1001 ();
 FILLCELL_X32 FILLER_60_1033 ();
 FILLCELL_X32 FILLER_60_1065 ();
 FILLCELL_X32 FILLER_60_1097 ();
 FILLCELL_X32 FILLER_60_1129 ();
 FILLCELL_X32 FILLER_60_1161 ();
 FILLCELL_X32 FILLER_60_1193 ();
 FILLCELL_X32 FILLER_60_1225 ();
 FILLCELL_X32 FILLER_60_1257 ();
 FILLCELL_X16 FILLER_60_1289 ();
 FILLCELL_X4 FILLER_60_1305 ();
 FILLCELL_X2 FILLER_60_1309 ();
 FILLCELL_X1 FILLER_60_1321 ();
 FILLCELL_X1 FILLER_60_1324 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X4 FILLER_61_65 ();
 FILLCELL_X2 FILLER_61_69 ();
 FILLCELL_X2 FILLER_61_77 ();
 FILLCELL_X8 FILLER_61_89 ();
 FILLCELL_X16 FILLER_61_110 ();
 FILLCELL_X4 FILLER_61_126 ();
 FILLCELL_X2 FILLER_61_130 ();
 FILLCELL_X4 FILLER_61_139 ();
 FILLCELL_X32 FILLER_61_147 ();
 FILLCELL_X32 FILLER_61_179 ();
 FILLCELL_X32 FILLER_61_211 ();
 FILLCELL_X32 FILLER_61_243 ();
 FILLCELL_X32 FILLER_61_275 ();
 FILLCELL_X32 FILLER_61_307 ();
 FILLCELL_X32 FILLER_61_339 ();
 FILLCELL_X32 FILLER_61_371 ();
 FILLCELL_X32 FILLER_61_403 ();
 FILLCELL_X32 FILLER_61_435 ();
 FILLCELL_X32 FILLER_61_467 ();
 FILLCELL_X32 FILLER_61_499 ();
 FILLCELL_X32 FILLER_61_531 ();
 FILLCELL_X32 FILLER_61_563 ();
 FILLCELL_X32 FILLER_61_595 ();
 FILLCELL_X16 FILLER_61_627 ();
 FILLCELL_X2 FILLER_61_643 ();
 FILLCELL_X4 FILLER_61_651 ();
 FILLCELL_X2 FILLER_61_655 ();
 FILLCELL_X1 FILLER_61_657 ();
 FILLCELL_X2 FILLER_61_663 ();
 FILLCELL_X8 FILLER_61_686 ();
 FILLCELL_X1 FILLER_61_694 ();
 FILLCELL_X32 FILLER_61_716 ();
 FILLCELL_X32 FILLER_61_757 ();
 FILLCELL_X32 FILLER_61_789 ();
 FILLCELL_X32 FILLER_61_821 ();
 FILLCELL_X32 FILLER_61_853 ();
 FILLCELL_X32 FILLER_61_885 ();
 FILLCELL_X32 FILLER_61_917 ();
 FILLCELL_X32 FILLER_61_949 ();
 FILLCELL_X32 FILLER_61_981 ();
 FILLCELL_X32 FILLER_61_1013 ();
 FILLCELL_X32 FILLER_61_1045 ();
 FILLCELL_X32 FILLER_61_1077 ();
 FILLCELL_X32 FILLER_61_1109 ();
 FILLCELL_X32 FILLER_61_1141 ();
 FILLCELL_X32 FILLER_61_1173 ();
 FILLCELL_X32 FILLER_61_1205 ();
 FILLCELL_X16 FILLER_61_1237 ();
 FILLCELL_X8 FILLER_61_1253 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X8 FILLER_61_1296 ();
 FILLCELL_X4 FILLER_61_1304 ();
 FILLCELL_X2 FILLER_61_1308 ();
 FILLCELL_X1 FILLER_61_1310 ();
 FILLCELL_X1 FILLER_61_1313 ();
 FILLCELL_X1 FILLER_61_1317 ();
 FILLCELL_X1 FILLER_61_1323 ();
 FILLCELL_X1 FILLER_61_1327 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X1 FILLER_62_33 ();
 FILLCELL_X16 FILLER_62_54 ();
 FILLCELL_X2 FILLER_62_70 ();
 FILLCELL_X8 FILLER_62_85 ();
 FILLCELL_X1 FILLER_62_93 ();
 FILLCELL_X2 FILLER_62_112 ();
 FILLCELL_X4 FILLER_62_117 ();
 FILLCELL_X4 FILLER_62_131 ();
 FILLCELL_X2 FILLER_62_169 ();
 FILLCELL_X2 FILLER_62_173 ();
 FILLCELL_X1 FILLER_62_175 ();
 FILLCELL_X32 FILLER_62_180 ();
 FILLCELL_X32 FILLER_62_212 ();
 FILLCELL_X32 FILLER_62_244 ();
 FILLCELL_X32 FILLER_62_276 ();
 FILLCELL_X32 FILLER_62_308 ();
 FILLCELL_X32 FILLER_62_340 ();
 FILLCELL_X32 FILLER_62_372 ();
 FILLCELL_X32 FILLER_62_404 ();
 FILLCELL_X32 FILLER_62_436 ();
 FILLCELL_X32 FILLER_62_468 ();
 FILLCELL_X32 FILLER_62_500 ();
 FILLCELL_X32 FILLER_62_532 ();
 FILLCELL_X32 FILLER_62_564 ();
 FILLCELL_X32 FILLER_62_596 ();
 FILLCELL_X2 FILLER_62_628 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X8 FILLER_62_664 ();
 FILLCELL_X16 FILLER_62_674 ();
 FILLCELL_X8 FILLER_62_690 ();
 FILLCELL_X4 FILLER_62_698 ();
 FILLCELL_X2 FILLER_62_702 ();
 FILLCELL_X4 FILLER_62_711 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X8 FILLER_62_1304 ();
 FILLCELL_X4 FILLER_62_1312 ();
 FILLCELL_X2 FILLER_63_1 ();
 FILLCELL_X4 FILLER_63_6 ();
 FILLCELL_X2 FILLER_63_10 ();
 FILLCELL_X8 FILLER_63_15 ();
 FILLCELL_X4 FILLER_63_23 ();
 FILLCELL_X2 FILLER_63_27 ();
 FILLCELL_X1 FILLER_63_29 ();
 FILLCELL_X4 FILLER_63_47 ();
 FILLCELL_X2 FILLER_63_51 ();
 FILLCELL_X16 FILLER_63_63 ();
 FILLCELL_X8 FILLER_63_79 ();
 FILLCELL_X2 FILLER_63_87 ();
 FILLCELL_X2 FILLER_63_107 ();
 FILLCELL_X1 FILLER_63_109 ();
 FILLCELL_X16 FILLER_63_119 ();
 FILLCELL_X2 FILLER_63_146 ();
 FILLCELL_X4 FILLER_63_154 ();
 FILLCELL_X4 FILLER_63_168 ();
 FILLCELL_X1 FILLER_63_172 ();
 FILLCELL_X32 FILLER_63_182 ();
 FILLCELL_X32 FILLER_63_214 ();
 FILLCELL_X32 FILLER_63_246 ();
 FILLCELL_X32 FILLER_63_278 ();
 FILLCELL_X32 FILLER_63_310 ();
 FILLCELL_X32 FILLER_63_342 ();
 FILLCELL_X32 FILLER_63_374 ();
 FILLCELL_X32 FILLER_63_406 ();
 FILLCELL_X32 FILLER_63_438 ();
 FILLCELL_X32 FILLER_63_470 ();
 FILLCELL_X32 FILLER_63_502 ();
 FILLCELL_X32 FILLER_63_534 ();
 FILLCELL_X32 FILLER_63_566 ();
 FILLCELL_X32 FILLER_63_598 ();
 FILLCELL_X8 FILLER_63_630 ();
 FILLCELL_X4 FILLER_63_638 ();
 FILLCELL_X1 FILLER_63_642 ();
 FILLCELL_X2 FILLER_63_649 ();
 FILLCELL_X1 FILLER_63_651 ();
 FILLCELL_X16 FILLER_63_679 ();
 FILLCELL_X8 FILLER_63_695 ();
 FILLCELL_X2 FILLER_63_703 ();
 FILLCELL_X1 FILLER_63_705 ();
 FILLCELL_X8 FILLER_63_709 ();
 FILLCELL_X2 FILLER_63_717 ();
 FILLCELL_X4 FILLER_63_722 ();
 FILLCELL_X2 FILLER_63_726 ();
 FILLCELL_X1 FILLER_63_743 ();
 FILLCELL_X32 FILLER_63_750 ();
 FILLCELL_X32 FILLER_63_782 ();
 FILLCELL_X32 FILLER_63_814 ();
 FILLCELL_X32 FILLER_63_846 ();
 FILLCELL_X32 FILLER_63_878 ();
 FILLCELL_X32 FILLER_63_910 ();
 FILLCELL_X32 FILLER_63_942 ();
 FILLCELL_X32 FILLER_63_974 ();
 FILLCELL_X32 FILLER_63_1006 ();
 FILLCELL_X32 FILLER_63_1038 ();
 FILLCELL_X32 FILLER_63_1070 ();
 FILLCELL_X32 FILLER_63_1102 ();
 FILLCELL_X32 FILLER_63_1134 ();
 FILLCELL_X32 FILLER_63_1166 ();
 FILLCELL_X32 FILLER_63_1198 ();
 FILLCELL_X32 FILLER_63_1230 ();
 FILLCELL_X1 FILLER_63_1262 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X16 FILLER_63_1296 ();
 FILLCELL_X2 FILLER_63_1312 ();
 FILLCELL_X1 FILLER_63_1314 ();
 FILLCELL_X1 FILLER_63_1317 ();
 FILLCELL_X1 FILLER_63_1323 ();
 FILLCELL_X1 FILLER_63_1327 ();
 FILLCELL_X8 FILLER_64_4 ();
 FILLCELL_X2 FILLER_64_25 ();
 FILLCELL_X4 FILLER_64_45 ();
 FILLCELL_X2 FILLER_64_49 ();
 FILLCELL_X16 FILLER_64_55 ();
 FILLCELL_X4 FILLER_64_71 ();
 FILLCELL_X8 FILLER_64_81 ();
 FILLCELL_X4 FILLER_64_106 ();
 FILLCELL_X2 FILLER_64_122 ();
 FILLCELL_X16 FILLER_64_146 ();
 FILLCELL_X4 FILLER_64_162 ();
 FILLCELL_X2 FILLER_64_166 ();
 FILLCELL_X1 FILLER_64_180 ();
 FILLCELL_X2 FILLER_64_185 ();
 FILLCELL_X32 FILLER_64_191 ();
 FILLCELL_X32 FILLER_64_223 ();
 FILLCELL_X32 FILLER_64_255 ();
 FILLCELL_X32 FILLER_64_287 ();
 FILLCELL_X32 FILLER_64_319 ();
 FILLCELL_X32 FILLER_64_351 ();
 FILLCELL_X32 FILLER_64_383 ();
 FILLCELL_X32 FILLER_64_415 ();
 FILLCELL_X32 FILLER_64_447 ();
 FILLCELL_X32 FILLER_64_479 ();
 FILLCELL_X32 FILLER_64_511 ();
 FILLCELL_X32 FILLER_64_543 ();
 FILLCELL_X32 FILLER_64_575 ();
 FILLCELL_X16 FILLER_64_607 ();
 FILLCELL_X8 FILLER_64_623 ();
 FILLCELL_X4 FILLER_64_632 ();
 FILLCELL_X2 FILLER_64_636 ();
 FILLCELL_X8 FILLER_64_652 ();
 FILLCELL_X4 FILLER_64_660 ();
 FILLCELL_X1 FILLER_64_674 ();
 FILLCELL_X32 FILLER_64_680 ();
 FILLCELL_X2 FILLER_64_712 ();
 FILLCELL_X1 FILLER_64_714 ();
 FILLCELL_X2 FILLER_64_742 ();
 FILLCELL_X1 FILLER_64_744 ();
 FILLCELL_X32 FILLER_64_750 ();
 FILLCELL_X32 FILLER_64_782 ();
 FILLCELL_X32 FILLER_64_814 ();
 FILLCELL_X32 FILLER_64_846 ();
 FILLCELL_X32 FILLER_64_878 ();
 FILLCELL_X32 FILLER_64_910 ();
 FILLCELL_X32 FILLER_64_942 ();
 FILLCELL_X32 FILLER_64_974 ();
 FILLCELL_X32 FILLER_64_1006 ();
 FILLCELL_X32 FILLER_64_1038 ();
 FILLCELL_X32 FILLER_64_1070 ();
 FILLCELL_X32 FILLER_64_1102 ();
 FILLCELL_X32 FILLER_64_1134 ();
 FILLCELL_X32 FILLER_64_1166 ();
 FILLCELL_X32 FILLER_64_1198 ();
 FILLCELL_X32 FILLER_64_1230 ();
 FILLCELL_X32 FILLER_64_1262 ();
 FILLCELL_X16 FILLER_64_1294 ();
 FILLCELL_X1 FILLER_64_1310 ();
 FILLCELL_X2 FILLER_64_1326 ();
 FILLCELL_X1 FILLER_65_7 ();
 FILLCELL_X4 FILLER_65_11 ();
 FILLCELL_X1 FILLER_65_19 ();
 FILLCELL_X4 FILLER_65_34 ();
 FILLCELL_X2 FILLER_65_38 ();
 FILLCELL_X1 FILLER_65_40 ();
 FILLCELL_X16 FILLER_65_48 ();
 FILLCELL_X4 FILLER_65_64 ();
 FILLCELL_X1 FILLER_65_68 ();
 FILLCELL_X16 FILLER_65_90 ();
 FILLCELL_X2 FILLER_65_106 ();
 FILLCELL_X32 FILLER_65_118 ();
 FILLCELL_X16 FILLER_65_150 ();
 FILLCELL_X8 FILLER_65_166 ();
 FILLCELL_X2 FILLER_65_174 ();
 FILLCELL_X1 FILLER_65_176 ();
 FILLCELL_X32 FILLER_65_194 ();
 FILLCELL_X32 FILLER_65_226 ();
 FILLCELL_X32 FILLER_65_258 ();
 FILLCELL_X32 FILLER_65_290 ();
 FILLCELL_X32 FILLER_65_322 ();
 FILLCELL_X32 FILLER_65_354 ();
 FILLCELL_X32 FILLER_65_386 ();
 FILLCELL_X32 FILLER_65_418 ();
 FILLCELL_X32 FILLER_65_450 ();
 FILLCELL_X32 FILLER_65_482 ();
 FILLCELL_X32 FILLER_65_514 ();
 FILLCELL_X32 FILLER_65_546 ();
 FILLCELL_X32 FILLER_65_578 ();
 FILLCELL_X8 FILLER_65_610 ();
 FILLCELL_X2 FILLER_65_618 ();
 FILLCELL_X1 FILLER_65_620 ();
 FILLCELL_X16 FILLER_65_647 ();
 FILLCELL_X4 FILLER_65_663 ();
 FILLCELL_X2 FILLER_65_667 ();
 FILLCELL_X2 FILLER_65_672 ();
 FILLCELL_X32 FILLER_65_679 ();
 FILLCELL_X2 FILLER_65_711 ();
 FILLCELL_X4 FILLER_65_740 ();
 FILLCELL_X1 FILLER_65_744 ();
 FILLCELL_X32 FILLER_65_762 ();
 FILLCELL_X32 FILLER_65_794 ();
 FILLCELL_X32 FILLER_65_826 ();
 FILLCELL_X32 FILLER_65_858 ();
 FILLCELL_X32 FILLER_65_890 ();
 FILLCELL_X32 FILLER_65_922 ();
 FILLCELL_X32 FILLER_65_954 ();
 FILLCELL_X32 FILLER_65_986 ();
 FILLCELL_X32 FILLER_65_1018 ();
 FILLCELL_X32 FILLER_65_1050 ();
 FILLCELL_X32 FILLER_65_1082 ();
 FILLCELL_X32 FILLER_65_1114 ();
 FILLCELL_X32 FILLER_65_1146 ();
 FILLCELL_X32 FILLER_65_1178 ();
 FILLCELL_X32 FILLER_65_1210 ();
 FILLCELL_X16 FILLER_65_1242 ();
 FILLCELL_X4 FILLER_65_1258 ();
 FILLCELL_X1 FILLER_65_1262 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X8 FILLER_65_1296 ();
 FILLCELL_X4 FILLER_65_1304 ();
 FILLCELL_X2 FILLER_65_1308 ();
 FILLCELL_X1 FILLER_65_1310 ();
 FILLCELL_X1 FILLER_65_1316 ();
 FILLCELL_X1 FILLER_65_1327 ();
 FILLCELL_X2 FILLER_66_4 ();
 FILLCELL_X1 FILLER_66_6 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X16 FILLER_66_65 ();
 FILLCELL_X1 FILLER_66_81 ();
 FILLCELL_X32 FILLER_66_89 ();
 FILLCELL_X32 FILLER_66_121 ();
 FILLCELL_X32 FILLER_66_153 ();
 FILLCELL_X32 FILLER_66_185 ();
 FILLCELL_X32 FILLER_66_217 ();
 FILLCELL_X32 FILLER_66_249 ();
 FILLCELL_X32 FILLER_66_281 ();
 FILLCELL_X32 FILLER_66_313 ();
 FILLCELL_X32 FILLER_66_345 ();
 FILLCELL_X32 FILLER_66_377 ();
 FILLCELL_X32 FILLER_66_409 ();
 FILLCELL_X32 FILLER_66_441 ();
 FILLCELL_X32 FILLER_66_473 ();
 FILLCELL_X32 FILLER_66_505 ();
 FILLCELL_X32 FILLER_66_537 ();
 FILLCELL_X32 FILLER_66_569 ();
 FILLCELL_X16 FILLER_66_601 ();
 FILLCELL_X8 FILLER_66_617 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X4 FILLER_66_632 ();
 FILLCELL_X1 FILLER_66_636 ();
 FILLCELL_X32 FILLER_66_641 ();
 FILLCELL_X32 FILLER_66_673 ();
 FILLCELL_X8 FILLER_66_705 ();
 FILLCELL_X2 FILLER_66_713 ();
 FILLCELL_X1 FILLER_66_715 ();
 FILLCELL_X4 FILLER_66_730 ();
 FILLCELL_X2 FILLER_66_734 ();
 FILLCELL_X32 FILLER_66_741 ();
 FILLCELL_X32 FILLER_66_773 ();
 FILLCELL_X32 FILLER_66_805 ();
 FILLCELL_X32 FILLER_66_837 ();
 FILLCELL_X32 FILLER_66_869 ();
 FILLCELL_X32 FILLER_66_901 ();
 FILLCELL_X32 FILLER_66_933 ();
 FILLCELL_X32 FILLER_66_965 ();
 FILLCELL_X32 FILLER_66_997 ();
 FILLCELL_X32 FILLER_66_1029 ();
 FILLCELL_X32 FILLER_66_1061 ();
 FILLCELL_X32 FILLER_66_1093 ();
 FILLCELL_X32 FILLER_66_1125 ();
 FILLCELL_X32 FILLER_66_1157 ();
 FILLCELL_X32 FILLER_66_1189 ();
 FILLCELL_X32 FILLER_66_1221 ();
 FILLCELL_X32 FILLER_66_1253 ();
 FILLCELL_X16 FILLER_66_1285 ();
 FILLCELL_X8 FILLER_66_1301 ();
 FILLCELL_X2 FILLER_66_1309 ();
 FILLCELL_X4 FILLER_66_1313 ();
 FILLCELL_X1 FILLER_66_1320 ();
 FILLCELL_X8 FILLER_67_1 ();
 FILLCELL_X4 FILLER_67_9 ();
 FILLCELL_X2 FILLER_67_13 ();
 FILLCELL_X32 FILLER_67_25 ();
 FILLCELL_X16 FILLER_67_57 ();
 FILLCELL_X4 FILLER_67_73 ();
 FILLCELL_X1 FILLER_67_77 ();
 FILLCELL_X1 FILLER_67_91 ();
 FILLCELL_X16 FILLER_67_110 ();
 FILLCELL_X8 FILLER_67_126 ();
 FILLCELL_X4 FILLER_67_134 ();
 FILLCELL_X1 FILLER_67_155 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X16 FILLER_67_609 ();
 FILLCELL_X8 FILLER_67_625 ();
 FILLCELL_X2 FILLER_67_633 ();
 FILLCELL_X1 FILLER_67_635 ();
 FILLCELL_X32 FILLER_67_642 ();
 FILLCELL_X32 FILLER_67_674 ();
 FILLCELL_X4 FILLER_67_706 ();
 FILLCELL_X2 FILLER_67_710 ();
 FILLCELL_X16 FILLER_67_721 ();
 FILLCELL_X8 FILLER_67_737 ();
 FILLCELL_X16 FILLER_67_761 ();
 FILLCELL_X8 FILLER_67_777 ();
 FILLCELL_X4 FILLER_67_785 ();
 FILLCELL_X1 FILLER_67_789 ();
 FILLCELL_X32 FILLER_67_811 ();
 FILLCELL_X32 FILLER_67_843 ();
 FILLCELL_X32 FILLER_67_875 ();
 FILLCELL_X32 FILLER_67_907 ();
 FILLCELL_X32 FILLER_67_939 ();
 FILLCELL_X32 FILLER_67_971 ();
 FILLCELL_X32 FILLER_67_1003 ();
 FILLCELL_X32 FILLER_67_1035 ();
 FILLCELL_X32 FILLER_67_1067 ();
 FILLCELL_X32 FILLER_67_1099 ();
 FILLCELL_X32 FILLER_67_1131 ();
 FILLCELL_X32 FILLER_67_1163 ();
 FILLCELL_X32 FILLER_67_1195 ();
 FILLCELL_X32 FILLER_67_1227 ();
 FILLCELL_X4 FILLER_67_1259 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X8 FILLER_67_1296 ();
 FILLCELL_X4 FILLER_67_1304 ();
 FILLCELL_X2 FILLER_67_1308 ();
 FILLCELL_X1 FILLER_67_1310 ();
 FILLCELL_X2 FILLER_67_1313 ();
 FILLCELL_X1 FILLER_67_1315 ();
 FILLCELL_X1 FILLER_67_1321 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X4 FILLER_68_129 ();
 FILLCELL_X2 FILLER_68_133 ();
 FILLCELL_X4 FILLER_68_142 ();
 FILLCELL_X1 FILLER_68_146 ();
 FILLCELL_X32 FILLER_68_151 ();
 FILLCELL_X32 FILLER_68_183 ();
 FILLCELL_X32 FILLER_68_215 ();
 FILLCELL_X32 FILLER_68_247 ();
 FILLCELL_X32 FILLER_68_279 ();
 FILLCELL_X32 FILLER_68_311 ();
 FILLCELL_X32 FILLER_68_343 ();
 FILLCELL_X32 FILLER_68_375 ();
 FILLCELL_X32 FILLER_68_407 ();
 FILLCELL_X32 FILLER_68_439 ();
 FILLCELL_X32 FILLER_68_471 ();
 FILLCELL_X32 FILLER_68_503 ();
 FILLCELL_X32 FILLER_68_535 ();
 FILLCELL_X32 FILLER_68_567 ();
 FILLCELL_X32 FILLER_68_599 ();
 FILLCELL_X8 FILLER_68_653 ();
 FILLCELL_X4 FILLER_68_661 ();
 FILLCELL_X2 FILLER_68_665 ();
 FILLCELL_X2 FILLER_68_669 ();
 FILLCELL_X16 FILLER_68_676 ();
 FILLCELL_X4 FILLER_68_692 ();
 FILLCELL_X2 FILLER_68_696 ();
 FILLCELL_X1 FILLER_68_719 ();
 FILLCELL_X16 FILLER_68_724 ();
 FILLCELL_X8 FILLER_68_740 ();
 FILLCELL_X1 FILLER_68_748 ();
 FILLCELL_X16 FILLER_68_772 ();
 FILLCELL_X1 FILLER_68_788 ();
 FILLCELL_X1 FILLER_68_793 ();
 FILLCELL_X32 FILLER_68_807 ();
 FILLCELL_X32 FILLER_68_839 ();
 FILLCELL_X32 FILLER_68_871 ();
 FILLCELL_X32 FILLER_68_903 ();
 FILLCELL_X32 FILLER_68_935 ();
 FILLCELL_X32 FILLER_68_967 ();
 FILLCELL_X32 FILLER_68_999 ();
 FILLCELL_X32 FILLER_68_1031 ();
 FILLCELL_X32 FILLER_68_1063 ();
 FILLCELL_X32 FILLER_68_1095 ();
 FILLCELL_X32 FILLER_68_1127 ();
 FILLCELL_X32 FILLER_68_1159 ();
 FILLCELL_X32 FILLER_68_1191 ();
 FILLCELL_X32 FILLER_68_1223 ();
 FILLCELL_X32 FILLER_68_1255 ();
 FILLCELL_X16 FILLER_68_1287 ();
 FILLCELL_X8 FILLER_68_1303 ();
 FILLCELL_X4 FILLER_68_1311 ();
 FILLCELL_X1 FILLER_68_1315 ();
 FILLCELL_X2 FILLER_68_1321 ();
 FILLCELL_X4 FILLER_69_1 ();
 FILLCELL_X1 FILLER_69_5 ();
 FILLCELL_X4 FILLER_69_12 ();
 FILLCELL_X1 FILLER_69_16 ();
 FILLCELL_X32 FILLER_69_20 ();
 FILLCELL_X1 FILLER_69_52 ();
 FILLCELL_X16 FILLER_69_63 ();
 FILLCELL_X8 FILLER_69_79 ();
 FILLCELL_X2 FILLER_69_87 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X2 FILLER_69_129 ();
 FILLCELL_X1 FILLER_69_131 ();
 FILLCELL_X4 FILLER_69_136 ();
 FILLCELL_X16 FILLER_69_143 ();
 FILLCELL_X8 FILLER_69_159 ();
 FILLCELL_X32 FILLER_69_184 ();
 FILLCELL_X32 FILLER_69_216 ();
 FILLCELL_X32 FILLER_69_248 ();
 FILLCELL_X32 FILLER_69_280 ();
 FILLCELL_X32 FILLER_69_312 ();
 FILLCELL_X32 FILLER_69_344 ();
 FILLCELL_X32 FILLER_69_376 ();
 FILLCELL_X32 FILLER_69_408 ();
 FILLCELL_X32 FILLER_69_440 ();
 FILLCELL_X32 FILLER_69_472 ();
 FILLCELL_X32 FILLER_69_504 ();
 FILLCELL_X32 FILLER_69_536 ();
 FILLCELL_X32 FILLER_69_568 ();
 FILLCELL_X8 FILLER_69_600 ();
 FILLCELL_X2 FILLER_69_608 ();
 FILLCELL_X2 FILLER_69_638 ();
 FILLCELL_X2 FILLER_69_644 ();
 FILLCELL_X4 FILLER_69_648 ();
 FILLCELL_X32 FILLER_69_677 ();
 FILLCELL_X4 FILLER_69_709 ();
 FILLCELL_X4 FILLER_69_717 ();
 FILLCELL_X2 FILLER_69_721 ();
 FILLCELL_X4 FILLER_69_733 ();
 FILLCELL_X8 FILLER_69_752 ();
 FILLCELL_X4 FILLER_69_760 ();
 FILLCELL_X1 FILLER_69_764 ();
 FILLCELL_X16 FILLER_69_769 ();
 FILLCELL_X4 FILLER_69_785 ();
 FILLCELL_X2 FILLER_69_789 ();
 FILLCELL_X1 FILLER_69_794 ();
 FILLCELL_X32 FILLER_69_824 ();
 FILLCELL_X32 FILLER_69_856 ();
 FILLCELL_X32 FILLER_69_888 ();
 FILLCELL_X32 FILLER_69_920 ();
 FILLCELL_X32 FILLER_69_952 ();
 FILLCELL_X32 FILLER_69_984 ();
 FILLCELL_X32 FILLER_69_1016 ();
 FILLCELL_X32 FILLER_69_1048 ();
 FILLCELL_X32 FILLER_69_1080 ();
 FILLCELL_X32 FILLER_69_1112 ();
 FILLCELL_X32 FILLER_69_1144 ();
 FILLCELL_X32 FILLER_69_1176 ();
 FILLCELL_X32 FILLER_69_1208 ();
 FILLCELL_X16 FILLER_69_1240 ();
 FILLCELL_X4 FILLER_69_1256 ();
 FILLCELL_X2 FILLER_69_1260 ();
 FILLCELL_X1 FILLER_69_1262 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X8 FILLER_69_1296 ();
 FILLCELL_X4 FILLER_69_1304 ();
 FILLCELL_X2 FILLER_69_1308 ();
 FILLCELL_X1 FILLER_69_1310 ();
 FILLCELL_X1 FILLER_69_1316 ();
 FILLCELL_X1 FILLER_69_1327 ();
 FILLCELL_X2 FILLER_70_1 ();
 FILLCELL_X1 FILLER_70_3 ();
 FILLCELL_X2 FILLER_70_7 ();
 FILLCELL_X1 FILLER_70_9 ();
 FILLCELL_X4 FILLER_70_40 ();
 FILLCELL_X4 FILLER_70_61 ();
 FILLCELL_X2 FILLER_70_65 ();
 FILLCELL_X16 FILLER_70_77 ();
 FILLCELL_X1 FILLER_70_93 ();
 FILLCELL_X8 FILLER_70_120 ();
 FILLCELL_X1 FILLER_70_128 ();
 FILLCELL_X2 FILLER_70_153 ();
 FILLCELL_X1 FILLER_70_155 ();
 FILLCELL_X4 FILLER_70_172 ();
 FILLCELL_X1 FILLER_70_176 ();
 FILLCELL_X32 FILLER_70_203 ();
 FILLCELL_X32 FILLER_70_235 ();
 FILLCELL_X32 FILLER_70_267 ();
 FILLCELL_X32 FILLER_70_299 ();
 FILLCELL_X32 FILLER_70_331 ();
 FILLCELL_X32 FILLER_70_363 ();
 FILLCELL_X32 FILLER_70_395 ();
 FILLCELL_X32 FILLER_70_427 ();
 FILLCELL_X32 FILLER_70_459 ();
 FILLCELL_X32 FILLER_70_491 ();
 FILLCELL_X32 FILLER_70_523 ();
 FILLCELL_X32 FILLER_70_555 ();
 FILLCELL_X16 FILLER_70_587 ();
 FILLCELL_X2 FILLER_70_603 ();
 FILLCELL_X1 FILLER_70_605 ();
 FILLCELL_X2 FILLER_70_610 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X16 FILLER_70_632 ();
 FILLCELL_X8 FILLER_70_648 ();
 FILLCELL_X2 FILLER_70_656 ();
 FILLCELL_X1 FILLER_70_658 ();
 FILLCELL_X32 FILLER_70_678 ();
 FILLCELL_X16 FILLER_70_710 ();
 FILLCELL_X8 FILLER_70_726 ();
 FILLCELL_X4 FILLER_70_734 ();
 FILLCELL_X8 FILLER_70_751 ();
 FILLCELL_X4 FILLER_70_759 ();
 FILLCELL_X1 FILLER_70_763 ();
 FILLCELL_X32 FILLER_70_775 ();
 FILLCELL_X8 FILLER_70_807 ();
 FILLCELL_X1 FILLER_70_815 ();
 FILLCELL_X32 FILLER_70_820 ();
 FILLCELL_X32 FILLER_70_852 ();
 FILLCELL_X32 FILLER_70_884 ();
 FILLCELL_X32 FILLER_70_916 ();
 FILLCELL_X32 FILLER_70_948 ();
 FILLCELL_X32 FILLER_70_980 ();
 FILLCELL_X32 FILLER_70_1012 ();
 FILLCELL_X32 FILLER_70_1044 ();
 FILLCELL_X32 FILLER_70_1076 ();
 FILLCELL_X32 FILLER_70_1108 ();
 FILLCELL_X32 FILLER_70_1140 ();
 FILLCELL_X32 FILLER_70_1172 ();
 FILLCELL_X32 FILLER_70_1204 ();
 FILLCELL_X32 FILLER_70_1236 ();
 FILLCELL_X32 FILLER_70_1268 ();
 FILLCELL_X16 FILLER_70_1300 ();
 FILLCELL_X2 FILLER_70_1326 ();
 FILLCELL_X2 FILLER_71_4 ();
 FILLCELL_X1 FILLER_71_6 ();
 FILLCELL_X8 FILLER_71_24 ();
 FILLCELL_X2 FILLER_71_57 ();
 FILLCELL_X8 FILLER_71_69 ();
 FILLCELL_X4 FILLER_71_77 ();
 FILLCELL_X2 FILLER_71_81 ();
 FILLCELL_X1 FILLER_71_83 ();
 FILLCELL_X2 FILLER_71_104 ();
 FILLCELL_X1 FILLER_71_106 ();
 FILLCELL_X8 FILLER_71_122 ();
 FILLCELL_X2 FILLER_71_130 ();
 FILLCELL_X1 FILLER_71_132 ();
 FILLCELL_X1 FILLER_71_142 ();
 FILLCELL_X8 FILLER_71_148 ();
 FILLCELL_X4 FILLER_71_156 ();
 FILLCELL_X1 FILLER_71_160 ();
 FILLCELL_X4 FILLER_71_172 ();
 FILLCELL_X2 FILLER_71_176 ();
 FILLCELL_X4 FILLER_71_183 ();
 FILLCELL_X2 FILLER_71_187 ();
 FILLCELL_X1 FILLER_71_189 ();
 FILLCELL_X32 FILLER_71_207 ();
 FILLCELL_X32 FILLER_71_239 ();
 FILLCELL_X32 FILLER_71_271 ();
 FILLCELL_X32 FILLER_71_303 ();
 FILLCELL_X32 FILLER_71_335 ();
 FILLCELL_X32 FILLER_71_367 ();
 FILLCELL_X32 FILLER_71_399 ();
 FILLCELL_X32 FILLER_71_431 ();
 FILLCELL_X32 FILLER_71_463 ();
 FILLCELL_X32 FILLER_71_495 ();
 FILLCELL_X32 FILLER_71_527 ();
 FILLCELL_X32 FILLER_71_559 ();
 FILLCELL_X8 FILLER_71_591 ();
 FILLCELL_X1 FILLER_71_599 ();
 FILLCELL_X16 FILLER_71_628 ();
 FILLCELL_X4 FILLER_71_644 ();
 FILLCELL_X2 FILLER_71_648 ();
 FILLCELL_X1 FILLER_71_650 ();
 FILLCELL_X32 FILLER_71_664 ();
 FILLCELL_X4 FILLER_71_696 ();
 FILLCELL_X2 FILLER_71_700 ();
 FILLCELL_X32 FILLER_71_712 ();
 FILLCELL_X2 FILLER_71_749 ();
 FILLCELL_X1 FILLER_71_751 ();
 FILLCELL_X16 FILLER_71_773 ();
 FILLCELL_X8 FILLER_71_789 ();
 FILLCELL_X4 FILLER_71_797 ();
 FILLCELL_X2 FILLER_71_801 ();
 FILLCELL_X1 FILLER_71_803 ();
 FILLCELL_X32 FILLER_71_821 ();
 FILLCELL_X32 FILLER_71_853 ();
 FILLCELL_X32 FILLER_71_885 ();
 FILLCELL_X32 FILLER_71_917 ();
 FILLCELL_X32 FILLER_71_949 ();
 FILLCELL_X32 FILLER_71_981 ();
 FILLCELL_X32 FILLER_71_1013 ();
 FILLCELL_X32 FILLER_71_1045 ();
 FILLCELL_X32 FILLER_71_1077 ();
 FILLCELL_X32 FILLER_71_1109 ();
 FILLCELL_X32 FILLER_71_1141 ();
 FILLCELL_X32 FILLER_71_1173 ();
 FILLCELL_X32 FILLER_71_1205 ();
 FILLCELL_X16 FILLER_71_1237 ();
 FILLCELL_X8 FILLER_71_1253 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X16 FILLER_71_1296 ();
 FILLCELL_X1 FILLER_71_1312 ();
 FILLCELL_X2 FILLER_72_5 ();
 FILLCELL_X1 FILLER_72_7 ();
 FILLCELL_X4 FILLER_72_50 ();
 FILLCELL_X1 FILLER_72_54 ();
 FILLCELL_X32 FILLER_72_59 ();
 FILLCELL_X2 FILLER_72_91 ();
 FILLCELL_X1 FILLER_72_93 ();
 FILLCELL_X32 FILLER_72_98 ();
 FILLCELL_X8 FILLER_72_130 ();
 FILLCELL_X4 FILLER_72_138 ();
 FILLCELL_X2 FILLER_72_142 ();
 FILLCELL_X32 FILLER_72_166 ();
 FILLCELL_X32 FILLER_72_198 ();
 FILLCELL_X32 FILLER_72_230 ();
 FILLCELL_X32 FILLER_72_262 ();
 FILLCELL_X32 FILLER_72_294 ();
 FILLCELL_X32 FILLER_72_326 ();
 FILLCELL_X32 FILLER_72_358 ();
 FILLCELL_X32 FILLER_72_390 ();
 FILLCELL_X32 FILLER_72_422 ();
 FILLCELL_X32 FILLER_72_454 ();
 FILLCELL_X32 FILLER_72_486 ();
 FILLCELL_X32 FILLER_72_518 ();
 FILLCELL_X32 FILLER_72_550 ();
 FILLCELL_X16 FILLER_72_582 ();
 FILLCELL_X1 FILLER_72_598 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X16 FILLER_72_632 ();
 FILLCELL_X8 FILLER_72_648 ();
 FILLCELL_X1 FILLER_72_656 ();
 FILLCELL_X16 FILLER_72_665 ();
 FILLCELL_X1 FILLER_72_681 ();
 FILLCELL_X16 FILLER_72_684 ();
 FILLCELL_X8 FILLER_72_700 ();
 FILLCELL_X8 FILLER_72_722 ();
 FILLCELL_X16 FILLER_72_735 ();
 FILLCELL_X8 FILLER_72_751 ();
 FILLCELL_X1 FILLER_72_766 ();
 FILLCELL_X4 FILLER_72_773 ();
 FILLCELL_X1 FILLER_72_777 ();
 FILLCELL_X4 FILLER_72_784 ();
 FILLCELL_X1 FILLER_72_788 ();
 FILLCELL_X4 FILLER_72_799 ();
 FILLCELL_X32 FILLER_72_812 ();
 FILLCELL_X32 FILLER_72_844 ();
 FILLCELL_X32 FILLER_72_876 ();
 FILLCELL_X32 FILLER_72_908 ();
 FILLCELL_X32 FILLER_72_940 ();
 FILLCELL_X32 FILLER_72_972 ();
 FILLCELL_X32 FILLER_72_1004 ();
 FILLCELL_X32 FILLER_72_1036 ();
 FILLCELL_X32 FILLER_72_1068 ();
 FILLCELL_X32 FILLER_72_1100 ();
 FILLCELL_X32 FILLER_72_1132 ();
 FILLCELL_X32 FILLER_72_1164 ();
 FILLCELL_X32 FILLER_72_1196 ();
 FILLCELL_X32 FILLER_72_1228 ();
 FILLCELL_X32 FILLER_72_1260 ();
 FILLCELL_X16 FILLER_72_1292 ();
 FILLCELL_X8 FILLER_72_1308 ();
 FILLCELL_X1 FILLER_73_9 ();
 FILLCELL_X16 FILLER_73_24 ();
 FILLCELL_X1 FILLER_73_40 ();
 FILLCELL_X32 FILLER_73_49 ();
 FILLCELL_X32 FILLER_73_81 ();
 FILLCELL_X32 FILLER_73_113 ();
 FILLCELL_X2 FILLER_73_145 ();
 FILLCELL_X1 FILLER_73_147 ();
 FILLCELL_X1 FILLER_73_157 ();
 FILLCELL_X1 FILLER_73_165 ();
 FILLCELL_X1 FILLER_73_176 ();
 FILLCELL_X2 FILLER_73_185 ();
 FILLCELL_X32 FILLER_73_204 ();
 FILLCELL_X32 FILLER_73_236 ();
 FILLCELL_X32 FILLER_73_268 ();
 FILLCELL_X32 FILLER_73_300 ();
 FILLCELL_X32 FILLER_73_332 ();
 FILLCELL_X32 FILLER_73_364 ();
 FILLCELL_X32 FILLER_73_396 ();
 FILLCELL_X32 FILLER_73_428 ();
 FILLCELL_X32 FILLER_73_460 ();
 FILLCELL_X32 FILLER_73_492 ();
 FILLCELL_X32 FILLER_73_524 ();
 FILLCELL_X32 FILLER_73_556 ();
 FILLCELL_X32 FILLER_73_588 ();
 FILLCELL_X2 FILLER_73_620 ();
 FILLCELL_X1 FILLER_73_622 ();
 FILLCELL_X4 FILLER_73_629 ();
 FILLCELL_X2 FILLER_73_650 ();
 FILLCELL_X1 FILLER_73_656 ();
 FILLCELL_X2 FILLER_73_661 ();
 FILLCELL_X2 FILLER_73_677 ();
 FILLCELL_X1 FILLER_73_679 ();
 FILLCELL_X16 FILLER_73_684 ();
 FILLCELL_X1 FILLER_73_700 ();
 FILLCELL_X2 FILLER_73_722 ();
 FILLCELL_X1 FILLER_73_724 ();
 FILLCELL_X1 FILLER_73_733 ();
 FILLCELL_X32 FILLER_73_738 ();
 FILLCELL_X16 FILLER_73_770 ();
 FILLCELL_X8 FILLER_73_786 ();
 FILLCELL_X1 FILLER_73_794 ();
 FILLCELL_X32 FILLER_73_806 ();
 FILLCELL_X32 FILLER_73_838 ();
 FILLCELL_X32 FILLER_73_870 ();
 FILLCELL_X32 FILLER_73_902 ();
 FILLCELL_X32 FILLER_73_934 ();
 FILLCELL_X32 FILLER_73_966 ();
 FILLCELL_X32 FILLER_73_998 ();
 FILLCELL_X32 FILLER_73_1030 ();
 FILLCELL_X32 FILLER_73_1062 ();
 FILLCELL_X32 FILLER_73_1094 ();
 FILLCELL_X32 FILLER_73_1126 ();
 FILLCELL_X32 FILLER_73_1158 ();
 FILLCELL_X32 FILLER_73_1190 ();
 FILLCELL_X32 FILLER_73_1222 ();
 FILLCELL_X8 FILLER_73_1254 ();
 FILLCELL_X1 FILLER_73_1262 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X16 FILLER_73_1296 ();
 FILLCELL_X2 FILLER_73_1312 ();
 FILLCELL_X1 FILLER_73_1324 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X8 FILLER_74_97 ();
 FILLCELL_X4 FILLER_74_105 ();
 FILLCELL_X2 FILLER_74_109 ();
 FILLCELL_X1 FILLER_74_111 ();
 FILLCELL_X16 FILLER_74_128 ();
 FILLCELL_X8 FILLER_74_144 ();
 FILLCELL_X2 FILLER_74_152 ();
 FILLCELL_X1 FILLER_74_154 ();
 FILLCELL_X2 FILLER_74_160 ();
 FILLCELL_X8 FILLER_74_173 ();
 FILLCELL_X1 FILLER_74_181 ();
 FILLCELL_X1 FILLER_74_186 ();
 FILLCELL_X1 FILLER_74_199 ();
 FILLCELL_X16 FILLER_74_234 ();
 FILLCELL_X4 FILLER_74_250 ();
 FILLCELL_X2 FILLER_74_254 ();
 FILLCELL_X1 FILLER_74_256 ();
 FILLCELL_X32 FILLER_74_270 ();
 FILLCELL_X32 FILLER_74_302 ();
 FILLCELL_X32 FILLER_74_334 ();
 FILLCELL_X32 FILLER_74_366 ();
 FILLCELL_X32 FILLER_74_398 ();
 FILLCELL_X32 FILLER_74_430 ();
 FILLCELL_X32 FILLER_74_462 ();
 FILLCELL_X32 FILLER_74_494 ();
 FILLCELL_X32 FILLER_74_526 ();
 FILLCELL_X32 FILLER_74_558 ();
 FILLCELL_X32 FILLER_74_590 ();
 FILLCELL_X8 FILLER_74_622 ();
 FILLCELL_X1 FILLER_74_630 ();
 FILLCELL_X4 FILLER_74_638 ();
 FILLCELL_X2 FILLER_74_642 ();
 FILLCELL_X1 FILLER_74_644 ();
 FILLCELL_X16 FILLER_74_662 ();
 FILLCELL_X1 FILLER_74_678 ();
 FILLCELL_X4 FILLER_74_707 ();
 FILLCELL_X2 FILLER_74_735 ();
 FILLCELL_X32 FILLER_74_747 ();
 FILLCELL_X16 FILLER_74_779 ();
 FILLCELL_X1 FILLER_74_795 ();
 FILLCELL_X32 FILLER_74_799 ();
 FILLCELL_X32 FILLER_74_831 ();
 FILLCELL_X32 FILLER_74_863 ();
 FILLCELL_X32 FILLER_74_895 ();
 FILLCELL_X32 FILLER_74_927 ();
 FILLCELL_X32 FILLER_74_959 ();
 FILLCELL_X32 FILLER_74_991 ();
 FILLCELL_X32 FILLER_74_1023 ();
 FILLCELL_X32 FILLER_74_1055 ();
 FILLCELL_X32 FILLER_74_1087 ();
 FILLCELL_X32 FILLER_74_1119 ();
 FILLCELL_X32 FILLER_74_1151 ();
 FILLCELL_X32 FILLER_74_1183 ();
 FILLCELL_X32 FILLER_74_1215 ();
 FILLCELL_X32 FILLER_74_1247 ();
 FILLCELL_X32 FILLER_74_1279 ();
 FILLCELL_X2 FILLER_74_1311 ();
 FILLCELL_X1 FILLER_74_1313 ();
 FILLCELL_X2 FILLER_74_1319 ();
 FILLCELL_X1 FILLER_74_1323 ();
 FILLCELL_X1 FILLER_74_1327 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X8 FILLER_75_65 ();
 FILLCELL_X4 FILLER_75_73 ();
 FILLCELL_X1 FILLER_75_77 ();
 FILLCELL_X2 FILLER_75_81 ();
 FILLCELL_X4 FILLER_75_102 ();
 FILLCELL_X1 FILLER_75_106 ();
 FILLCELL_X2 FILLER_75_116 ();
 FILLCELL_X1 FILLER_75_118 ();
 FILLCELL_X1 FILLER_75_128 ();
 FILLCELL_X8 FILLER_75_148 ();
 FILLCELL_X4 FILLER_75_156 ();
 FILLCELL_X2 FILLER_75_160 ();
 FILLCELL_X1 FILLER_75_162 ();
 FILLCELL_X1 FILLER_75_167 ();
 FILLCELL_X32 FILLER_75_180 ();
 FILLCELL_X32 FILLER_75_212 ();
 FILLCELL_X32 FILLER_75_244 ();
 FILLCELL_X32 FILLER_75_276 ();
 FILLCELL_X32 FILLER_75_308 ();
 FILLCELL_X32 FILLER_75_340 ();
 FILLCELL_X32 FILLER_75_372 ();
 FILLCELL_X32 FILLER_75_404 ();
 FILLCELL_X32 FILLER_75_436 ();
 FILLCELL_X32 FILLER_75_468 ();
 FILLCELL_X32 FILLER_75_500 ();
 FILLCELL_X32 FILLER_75_532 ();
 FILLCELL_X32 FILLER_75_564 ();
 FILLCELL_X32 FILLER_75_596 ();
 FILLCELL_X1 FILLER_75_628 ();
 FILLCELL_X32 FILLER_75_646 ();
 FILLCELL_X32 FILLER_75_678 ();
 FILLCELL_X16 FILLER_75_710 ();
 FILLCELL_X8 FILLER_75_726 ();
 FILLCELL_X4 FILLER_75_734 ();
 FILLCELL_X2 FILLER_75_738 ();
 FILLCELL_X16 FILLER_75_767 ();
 FILLCELL_X8 FILLER_75_783 ();
 FILLCELL_X4 FILLER_75_791 ();
 FILLCELL_X32 FILLER_75_809 ();
 FILLCELL_X32 FILLER_75_841 ();
 FILLCELL_X32 FILLER_75_873 ();
 FILLCELL_X32 FILLER_75_905 ();
 FILLCELL_X32 FILLER_75_937 ();
 FILLCELL_X32 FILLER_75_969 ();
 FILLCELL_X32 FILLER_75_1001 ();
 FILLCELL_X32 FILLER_75_1033 ();
 FILLCELL_X32 FILLER_75_1065 ();
 FILLCELL_X32 FILLER_75_1097 ();
 FILLCELL_X32 FILLER_75_1129 ();
 FILLCELL_X32 FILLER_75_1161 ();
 FILLCELL_X32 FILLER_75_1193 ();
 FILLCELL_X32 FILLER_75_1225 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X8 FILLER_75_1296 ();
 FILLCELL_X4 FILLER_75_1304 ();
 FILLCELL_X2 FILLER_75_1308 ();
 FILLCELL_X1 FILLER_75_1310 ();
 FILLCELL_X1 FILLER_75_1318 ();
 FILLCELL_X1 FILLER_75_1327 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X8 FILLER_76_65 ();
 FILLCELL_X2 FILLER_76_87 ();
 FILLCELL_X1 FILLER_76_89 ();
 FILLCELL_X32 FILLER_76_93 ();
 FILLCELL_X32 FILLER_76_125 ();
 FILLCELL_X4 FILLER_76_157 ();
 FILLCELL_X2 FILLER_76_161 ();
 FILLCELL_X1 FILLER_76_173 ();
 FILLCELL_X32 FILLER_76_179 ();
 FILLCELL_X32 FILLER_76_211 ();
 FILLCELL_X32 FILLER_76_243 ();
 FILLCELL_X32 FILLER_76_275 ();
 FILLCELL_X32 FILLER_76_307 ();
 FILLCELL_X32 FILLER_76_339 ();
 FILLCELL_X32 FILLER_76_371 ();
 FILLCELL_X32 FILLER_76_403 ();
 FILLCELL_X32 FILLER_76_435 ();
 FILLCELL_X32 FILLER_76_467 ();
 FILLCELL_X32 FILLER_76_499 ();
 FILLCELL_X32 FILLER_76_531 ();
 FILLCELL_X32 FILLER_76_563 ();
 FILLCELL_X32 FILLER_76_595 ();
 FILLCELL_X4 FILLER_76_627 ();
 FILLCELL_X16 FILLER_76_632 ();
 FILLCELL_X8 FILLER_76_648 ();
 FILLCELL_X4 FILLER_76_656 ();
 FILLCELL_X2 FILLER_76_660 ();
 FILLCELL_X32 FILLER_76_669 ();
 FILLCELL_X4 FILLER_76_701 ();
 FILLCELL_X2 FILLER_76_705 ();
 FILLCELL_X1 FILLER_76_707 ();
 FILLCELL_X32 FILLER_76_713 ();
 FILLCELL_X32 FILLER_76_747 ();
 FILLCELL_X16 FILLER_76_779 ();
 FILLCELL_X1 FILLER_76_795 ();
 FILLCELL_X32 FILLER_76_821 ();
 FILLCELL_X32 FILLER_76_853 ();
 FILLCELL_X32 FILLER_76_885 ();
 FILLCELL_X32 FILLER_76_917 ();
 FILLCELL_X32 FILLER_76_949 ();
 FILLCELL_X32 FILLER_76_981 ();
 FILLCELL_X32 FILLER_76_1013 ();
 FILLCELL_X32 FILLER_76_1045 ();
 FILLCELL_X32 FILLER_76_1077 ();
 FILLCELL_X32 FILLER_76_1109 ();
 FILLCELL_X32 FILLER_76_1141 ();
 FILLCELL_X32 FILLER_76_1173 ();
 FILLCELL_X32 FILLER_76_1205 ();
 FILLCELL_X32 FILLER_76_1237 ();
 FILLCELL_X32 FILLER_76_1269 ();
 FILLCELL_X8 FILLER_76_1301 ();
 FILLCELL_X2 FILLER_76_1309 ();
 FILLCELL_X1 FILLER_76_1313 ();
 FILLCELL_X1 FILLER_76_1319 ();
 FILLCELL_X8 FILLER_77_1 ();
 FILLCELL_X4 FILLER_77_9 ();
 FILLCELL_X2 FILLER_77_13 ();
 FILLCELL_X1 FILLER_77_15 ();
 FILLCELL_X1 FILLER_77_40 ();
 FILLCELL_X8 FILLER_77_54 ();
 FILLCELL_X2 FILLER_77_62 ();
 FILLCELL_X1 FILLER_77_64 ();
 FILLCELL_X1 FILLER_77_73 ();
 FILLCELL_X8 FILLER_77_98 ();
 FILLCELL_X1 FILLER_77_106 ();
 FILLCELL_X4 FILLER_77_117 ();
 FILLCELL_X4 FILLER_77_131 ();
 FILLCELL_X16 FILLER_77_139 ();
 FILLCELL_X4 FILLER_77_155 ();
 FILLCELL_X2 FILLER_77_159 ();
 FILLCELL_X1 FILLER_77_161 ();
 FILLCELL_X8 FILLER_77_167 ();
 FILLCELL_X4 FILLER_77_175 ();
 FILLCELL_X2 FILLER_77_179 ();
 FILLCELL_X1 FILLER_77_181 ();
 FILLCELL_X2 FILLER_77_186 ();
 FILLCELL_X4 FILLER_77_194 ();
 FILLCELL_X2 FILLER_77_198 ();
 FILLCELL_X2 FILLER_77_202 ();
 FILLCELL_X32 FILLER_77_229 ();
 FILLCELL_X32 FILLER_77_261 ();
 FILLCELL_X32 FILLER_77_293 ();
 FILLCELL_X32 FILLER_77_325 ();
 FILLCELL_X32 FILLER_77_357 ();
 FILLCELL_X32 FILLER_77_389 ();
 FILLCELL_X32 FILLER_77_421 ();
 FILLCELL_X32 FILLER_77_453 ();
 FILLCELL_X32 FILLER_77_485 ();
 FILLCELL_X32 FILLER_77_517 ();
 FILLCELL_X32 FILLER_77_549 ();
 FILLCELL_X32 FILLER_77_581 ();
 FILLCELL_X32 FILLER_77_613 ();
 FILLCELL_X4 FILLER_77_645 ();
 FILLCELL_X2 FILLER_77_649 ();
 FILLCELL_X1 FILLER_77_656 ();
 FILLCELL_X16 FILLER_77_660 ();
 FILLCELL_X4 FILLER_77_676 ();
 FILLCELL_X2 FILLER_77_680 ();
 FILLCELL_X1 FILLER_77_682 ();
 FILLCELL_X8 FILLER_77_688 ();
 FILLCELL_X2 FILLER_77_696 ();
 FILLCELL_X32 FILLER_77_703 ();
 FILLCELL_X32 FILLER_77_735 ();
 FILLCELL_X16 FILLER_77_767 ();
 FILLCELL_X8 FILLER_77_783 ();
 FILLCELL_X1 FILLER_77_814 ();
 FILLCELL_X2 FILLER_77_819 ();
 FILLCELL_X32 FILLER_77_825 ();
 FILLCELL_X32 FILLER_77_857 ();
 FILLCELL_X32 FILLER_77_889 ();
 FILLCELL_X32 FILLER_77_921 ();
 FILLCELL_X32 FILLER_77_953 ();
 FILLCELL_X32 FILLER_77_985 ();
 FILLCELL_X32 FILLER_77_1017 ();
 FILLCELL_X32 FILLER_77_1049 ();
 FILLCELL_X32 FILLER_77_1081 ();
 FILLCELL_X32 FILLER_77_1113 ();
 FILLCELL_X32 FILLER_77_1145 ();
 FILLCELL_X32 FILLER_77_1177 ();
 FILLCELL_X32 FILLER_77_1209 ();
 FILLCELL_X16 FILLER_77_1241 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X16 FILLER_77_1296 ();
 FILLCELL_X2 FILLER_77_1312 ();
 FILLCELL_X4 FILLER_77_1324 ();
 FILLCELL_X8 FILLER_78_1 ();
 FILLCELL_X2 FILLER_78_9 ();
 FILLCELL_X4 FILLER_78_20 ();
 FILLCELL_X2 FILLER_78_24 ();
 FILLCELL_X16 FILLER_78_30 ();
 FILLCELL_X4 FILLER_78_46 ();
 FILLCELL_X2 FILLER_78_67 ();
 FILLCELL_X1 FILLER_78_69 ();
 FILLCELL_X16 FILLER_78_78 ();
 FILLCELL_X8 FILLER_78_94 ();
 FILLCELL_X4 FILLER_78_102 ();
 FILLCELL_X1 FILLER_78_106 ();
 FILLCELL_X1 FILLER_78_112 ();
 FILLCELL_X1 FILLER_78_139 ();
 FILLCELL_X16 FILLER_78_143 ();
 FILLCELL_X2 FILLER_78_159 ();
 FILLCELL_X1 FILLER_78_161 ();
 FILLCELL_X4 FILLER_78_181 ();
 FILLCELL_X2 FILLER_78_185 ();
 FILLCELL_X1 FILLER_78_187 ();
 FILLCELL_X32 FILLER_78_216 ();
 FILLCELL_X16 FILLER_78_248 ();
 FILLCELL_X8 FILLER_78_264 ();
 FILLCELL_X2 FILLER_78_272 ();
 FILLCELL_X1 FILLER_78_274 ();
 FILLCELL_X32 FILLER_78_282 ();
 FILLCELL_X32 FILLER_78_314 ();
 FILLCELL_X32 FILLER_78_346 ();
 FILLCELL_X32 FILLER_78_378 ();
 FILLCELL_X32 FILLER_78_410 ();
 FILLCELL_X32 FILLER_78_442 ();
 FILLCELL_X32 FILLER_78_474 ();
 FILLCELL_X32 FILLER_78_506 ();
 FILLCELL_X32 FILLER_78_538 ();
 FILLCELL_X32 FILLER_78_570 ();
 FILLCELL_X16 FILLER_78_602 ();
 FILLCELL_X8 FILLER_78_618 ();
 FILLCELL_X4 FILLER_78_626 ();
 FILLCELL_X1 FILLER_78_630 ();
 FILLCELL_X4 FILLER_78_632 ();
 FILLCELL_X2 FILLER_78_636 ();
 FILLCELL_X8 FILLER_78_641 ();
 FILLCELL_X2 FILLER_78_649 ();
 FILLCELL_X1 FILLER_78_651 ();
 FILLCELL_X2 FILLER_78_661 ();
 FILLCELL_X1 FILLER_78_663 ();
 FILLCELL_X16 FILLER_78_668 ();
 FILLCELL_X4 FILLER_78_684 ();
 FILLCELL_X2 FILLER_78_688 ();
 FILLCELL_X4 FILLER_78_715 ();
 FILLCELL_X1 FILLER_78_719 ();
 FILLCELL_X4 FILLER_78_722 ();
 FILLCELL_X2 FILLER_78_726 ();
 FILLCELL_X1 FILLER_78_728 ();
 FILLCELL_X4 FILLER_78_733 ();
 FILLCELL_X2 FILLER_78_737 ();
 FILLCELL_X1 FILLER_78_739 ();
 FILLCELL_X8 FILLER_78_748 ();
 FILLCELL_X8 FILLER_78_780 ();
 FILLCELL_X1 FILLER_78_788 ();
 FILLCELL_X2 FILLER_78_804 ();
 FILLCELL_X1 FILLER_78_806 ();
 FILLCELL_X32 FILLER_78_826 ();
 FILLCELL_X32 FILLER_78_858 ();
 FILLCELL_X32 FILLER_78_890 ();
 FILLCELL_X32 FILLER_78_922 ();
 FILLCELL_X32 FILLER_78_954 ();
 FILLCELL_X32 FILLER_78_986 ();
 FILLCELL_X32 FILLER_78_1018 ();
 FILLCELL_X32 FILLER_78_1050 ();
 FILLCELL_X32 FILLER_78_1082 ();
 FILLCELL_X32 FILLER_78_1114 ();
 FILLCELL_X32 FILLER_78_1146 ();
 FILLCELL_X32 FILLER_78_1178 ();
 FILLCELL_X32 FILLER_78_1210 ();
 FILLCELL_X32 FILLER_78_1242 ();
 FILLCELL_X32 FILLER_78_1274 ();
 FILLCELL_X8 FILLER_78_1306 ();
 FILLCELL_X4 FILLER_78_1316 ();
 FILLCELL_X1 FILLER_79_1 ();
 FILLCELL_X4 FILLER_79_5 ();
 FILLCELL_X2 FILLER_79_9 ();
 FILLCELL_X1 FILLER_79_11 ();
 FILLCELL_X2 FILLER_79_25 ();
 FILLCELL_X1 FILLER_79_30 ();
 FILLCELL_X16 FILLER_79_41 ();
 FILLCELL_X8 FILLER_79_57 ();
 FILLCELL_X2 FILLER_79_65 ();
 FILLCELL_X4 FILLER_79_73 ();
 FILLCELL_X8 FILLER_79_79 ();
 FILLCELL_X2 FILLER_79_87 ();
 FILLCELL_X4 FILLER_79_104 ();
 FILLCELL_X8 FILLER_79_126 ();
 FILLCELL_X4 FILLER_79_134 ();
 FILLCELL_X2 FILLER_79_138 ();
 FILLCELL_X1 FILLER_79_140 ();
 FILLCELL_X16 FILLER_79_165 ();
 FILLCELL_X8 FILLER_79_181 ();
 FILLCELL_X4 FILLER_79_189 ();
 FILLCELL_X1 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_204 ();
 FILLCELL_X32 FILLER_79_236 ();
 FILLCELL_X32 FILLER_79_268 ();
 FILLCELL_X32 FILLER_79_300 ();
 FILLCELL_X32 FILLER_79_332 ();
 FILLCELL_X32 FILLER_79_364 ();
 FILLCELL_X32 FILLER_79_396 ();
 FILLCELL_X32 FILLER_79_428 ();
 FILLCELL_X32 FILLER_79_460 ();
 FILLCELL_X32 FILLER_79_492 ();
 FILLCELL_X32 FILLER_79_524 ();
 FILLCELL_X32 FILLER_79_556 ();
 FILLCELL_X32 FILLER_79_588 ();
 FILLCELL_X8 FILLER_79_620 ();
 FILLCELL_X4 FILLER_79_628 ();
 FILLCELL_X2 FILLER_79_632 ();
 FILLCELL_X16 FILLER_79_637 ();
 FILLCELL_X1 FILLER_79_660 ();
 FILLCELL_X2 FILLER_79_664 ();
 FILLCELL_X2 FILLER_79_669 ();
 FILLCELL_X4 FILLER_79_676 ();
 FILLCELL_X1 FILLER_79_680 ();
 FILLCELL_X2 FILLER_79_690 ();
 FILLCELL_X1 FILLER_79_692 ();
 FILLCELL_X1 FILLER_79_697 ();
 FILLCELL_X1 FILLER_79_726 ();
 FILLCELL_X1 FILLER_79_731 ();
 FILLCELL_X1 FILLER_79_736 ();
 FILLCELL_X4 FILLER_79_740 ();
 FILLCELL_X1 FILLER_79_744 ();
 FILLCELL_X4 FILLER_79_749 ();
 FILLCELL_X16 FILLER_79_764 ();
 FILLCELL_X8 FILLER_79_780 ();
 FILLCELL_X4 FILLER_79_788 ();
 FILLCELL_X2 FILLER_79_792 ();
 FILLCELL_X1 FILLER_79_794 ();
 FILLCELL_X32 FILLER_79_804 ();
 FILLCELL_X32 FILLER_79_836 ();
 FILLCELL_X32 FILLER_79_868 ();
 FILLCELL_X32 FILLER_79_900 ();
 FILLCELL_X32 FILLER_79_932 ();
 FILLCELL_X32 FILLER_79_964 ();
 FILLCELL_X32 FILLER_79_996 ();
 FILLCELL_X32 FILLER_79_1028 ();
 FILLCELL_X32 FILLER_79_1060 ();
 FILLCELL_X32 FILLER_79_1092 ();
 FILLCELL_X32 FILLER_79_1124 ();
 FILLCELL_X32 FILLER_79_1156 ();
 FILLCELL_X32 FILLER_79_1188 ();
 FILLCELL_X32 FILLER_79_1220 ();
 FILLCELL_X8 FILLER_79_1252 ();
 FILLCELL_X2 FILLER_79_1260 ();
 FILLCELL_X1 FILLER_79_1262 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X8 FILLER_79_1296 ();
 FILLCELL_X4 FILLER_79_1304 ();
 FILLCELL_X2 FILLER_79_1308 ();
 FILLCELL_X1 FILLER_79_1310 ();
 FILLCELL_X1 FILLER_79_1316 ();
 FILLCELL_X1 FILLER_79_1324 ();
 FILLCELL_X16 FILLER_80_1 ();
 FILLCELL_X2 FILLER_80_17 ();
 FILLCELL_X1 FILLER_80_31 ();
 FILLCELL_X32 FILLER_80_36 ();
 FILLCELL_X4 FILLER_80_68 ();
 FILLCELL_X2 FILLER_80_72 ();
 FILLCELL_X4 FILLER_80_89 ();
 FILLCELL_X32 FILLER_80_102 ();
 FILLCELL_X32 FILLER_80_134 ();
 FILLCELL_X32 FILLER_80_166 ();
 FILLCELL_X32 FILLER_80_198 ();
 FILLCELL_X32 FILLER_80_230 ();
 FILLCELL_X32 FILLER_80_262 ();
 FILLCELL_X32 FILLER_80_294 ();
 FILLCELL_X32 FILLER_80_326 ();
 FILLCELL_X32 FILLER_80_358 ();
 FILLCELL_X32 FILLER_80_390 ();
 FILLCELL_X32 FILLER_80_422 ();
 FILLCELL_X32 FILLER_80_454 ();
 FILLCELL_X32 FILLER_80_486 ();
 FILLCELL_X32 FILLER_80_518 ();
 FILLCELL_X32 FILLER_80_550 ();
 FILLCELL_X16 FILLER_80_582 ();
 FILLCELL_X2 FILLER_80_598 ();
 FILLCELL_X1 FILLER_80_600 ();
 FILLCELL_X1 FILLER_80_625 ();
 FILLCELL_X8 FILLER_80_632 ();
 FILLCELL_X4 FILLER_80_640 ();
 FILLCELL_X2 FILLER_80_659 ();
 FILLCELL_X4 FILLER_80_665 ();
 FILLCELL_X1 FILLER_80_669 ();
 FILLCELL_X8 FILLER_80_676 ();
 FILLCELL_X2 FILLER_80_684 ();
 FILLCELL_X1 FILLER_80_686 ();
 FILLCELL_X16 FILLER_80_701 ();
 FILLCELL_X8 FILLER_80_717 ();
 FILLCELL_X1 FILLER_80_725 ();
 FILLCELL_X32 FILLER_80_731 ();
 FILLCELL_X32 FILLER_80_763 ();
 FILLCELL_X32 FILLER_80_795 ();
 FILLCELL_X32 FILLER_80_827 ();
 FILLCELL_X32 FILLER_80_859 ();
 FILLCELL_X32 FILLER_80_891 ();
 FILLCELL_X32 FILLER_80_923 ();
 FILLCELL_X32 FILLER_80_955 ();
 FILLCELL_X32 FILLER_80_987 ();
 FILLCELL_X32 FILLER_80_1019 ();
 FILLCELL_X32 FILLER_80_1051 ();
 FILLCELL_X32 FILLER_80_1083 ();
 FILLCELL_X32 FILLER_80_1115 ();
 FILLCELL_X32 FILLER_80_1147 ();
 FILLCELL_X32 FILLER_80_1179 ();
 FILLCELL_X32 FILLER_80_1211 ();
 FILLCELL_X32 FILLER_80_1243 ();
 FILLCELL_X32 FILLER_80_1275 ();
 FILLCELL_X4 FILLER_80_1307 ();
 FILLCELL_X2 FILLER_80_1311 ();
 FILLCELL_X1 FILLER_80_1313 ();
 FILLCELL_X2 FILLER_80_1316 ();
 FILLCELL_X1 FILLER_80_1318 ();
 FILLCELL_X1 FILLER_80_1324 ();
 FILLCELL_X2 FILLER_81_1 ();
 FILLCELL_X1 FILLER_81_3 ();
 FILLCELL_X8 FILLER_81_7 ();
 FILLCELL_X4 FILLER_81_15 ();
 FILLCELL_X32 FILLER_81_29 ();
 FILLCELL_X1 FILLER_81_78 ();
 FILLCELL_X32 FILLER_81_83 ();
 FILLCELL_X16 FILLER_81_115 ();
 FILLCELL_X8 FILLER_81_131 ();
 FILLCELL_X4 FILLER_81_139 ();
 FILLCELL_X32 FILLER_81_160 ();
 FILLCELL_X8 FILLER_81_192 ();
 FILLCELL_X1 FILLER_81_200 ();
 FILLCELL_X32 FILLER_81_210 ();
 FILLCELL_X32 FILLER_81_242 ();
 FILLCELL_X32 FILLER_81_274 ();
 FILLCELL_X32 FILLER_81_306 ();
 FILLCELL_X32 FILLER_81_338 ();
 FILLCELL_X32 FILLER_81_370 ();
 FILLCELL_X32 FILLER_81_402 ();
 FILLCELL_X32 FILLER_81_434 ();
 FILLCELL_X32 FILLER_81_466 ();
 FILLCELL_X32 FILLER_81_498 ();
 FILLCELL_X32 FILLER_81_530 ();
 FILLCELL_X32 FILLER_81_562 ();
 FILLCELL_X16 FILLER_81_594 ();
 FILLCELL_X8 FILLER_81_610 ();
 FILLCELL_X1 FILLER_81_618 ();
 FILLCELL_X8 FILLER_81_625 ();
 FILLCELL_X2 FILLER_81_633 ();
 FILLCELL_X1 FILLER_81_635 ();
 FILLCELL_X4 FILLER_81_649 ();
 FILLCELL_X1 FILLER_81_653 ();
 FILLCELL_X8 FILLER_81_673 ();
 FILLCELL_X1 FILLER_81_681 ();
 FILLCELL_X2 FILLER_81_687 ();
 FILLCELL_X2 FILLER_81_691 ();
 FILLCELL_X1 FILLER_81_693 ();
 FILLCELL_X16 FILLER_81_700 ();
 FILLCELL_X4 FILLER_81_716 ();
 FILLCELL_X2 FILLER_81_720 ();
 FILLCELL_X32 FILLER_81_747 ();
 FILLCELL_X1 FILLER_81_779 ();
 FILLCELL_X8 FILLER_81_799 ();
 FILLCELL_X4 FILLER_81_807 ();
 FILLCELL_X32 FILLER_81_820 ();
 FILLCELL_X32 FILLER_81_852 ();
 FILLCELL_X32 FILLER_81_884 ();
 FILLCELL_X32 FILLER_81_916 ();
 FILLCELL_X32 FILLER_81_948 ();
 FILLCELL_X32 FILLER_81_980 ();
 FILLCELL_X32 FILLER_81_1012 ();
 FILLCELL_X32 FILLER_81_1044 ();
 FILLCELL_X32 FILLER_81_1076 ();
 FILLCELL_X32 FILLER_81_1108 ();
 FILLCELL_X32 FILLER_81_1140 ();
 FILLCELL_X32 FILLER_81_1172 ();
 FILLCELL_X32 FILLER_81_1204 ();
 FILLCELL_X16 FILLER_81_1236 ();
 FILLCELL_X8 FILLER_81_1252 ();
 FILLCELL_X2 FILLER_81_1260 ();
 FILLCELL_X1 FILLER_81_1262 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X8 FILLER_81_1296 ();
 FILLCELL_X4 FILLER_81_1304 ();
 FILLCELL_X2 FILLER_81_1308 ();
 FILLCELL_X1 FILLER_81_1310 ();
 FILLCELL_X1 FILLER_81_1321 ();
 FILLCELL_X1 FILLER_81_1327 ();
 FILLCELL_X4 FILLER_82_1 ();
 FILLCELL_X8 FILLER_82_8 ();
 FILLCELL_X4 FILLER_82_16 ();
 FILLCELL_X2 FILLER_82_20 ();
 FILLCELL_X8 FILLER_82_26 ();
 FILLCELL_X2 FILLER_82_34 ();
 FILLCELL_X16 FILLER_82_41 ();
 FILLCELL_X4 FILLER_82_57 ();
 FILLCELL_X2 FILLER_82_61 ();
 FILLCELL_X32 FILLER_82_67 ();
 FILLCELL_X32 FILLER_82_99 ();
 FILLCELL_X8 FILLER_82_131 ();
 FILLCELL_X2 FILLER_82_139 ();
 FILLCELL_X4 FILLER_82_148 ();
 FILLCELL_X1 FILLER_82_152 ();
 FILLCELL_X2 FILLER_82_167 ();
 FILLCELL_X1 FILLER_82_169 ();
 FILLCELL_X4 FILLER_82_180 ();
 FILLCELL_X2 FILLER_82_184 ();
 FILLCELL_X2 FILLER_82_190 ();
 FILLCELL_X1 FILLER_82_192 ();
 FILLCELL_X32 FILLER_82_216 ();
 FILLCELL_X32 FILLER_82_248 ();
 FILLCELL_X32 FILLER_82_280 ();
 FILLCELL_X32 FILLER_82_312 ();
 FILLCELL_X32 FILLER_82_344 ();
 FILLCELL_X32 FILLER_82_376 ();
 FILLCELL_X32 FILLER_82_408 ();
 FILLCELL_X32 FILLER_82_440 ();
 FILLCELL_X32 FILLER_82_472 ();
 FILLCELL_X32 FILLER_82_504 ();
 FILLCELL_X32 FILLER_82_536 ();
 FILLCELL_X32 FILLER_82_568 ();
 FILLCELL_X8 FILLER_82_600 ();
 FILLCELL_X2 FILLER_82_608 ();
 FILLCELL_X1 FILLER_82_610 ();
 FILLCELL_X2 FILLER_82_628 ();
 FILLCELL_X1 FILLER_82_630 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X8 FILLER_82_664 ();
 FILLCELL_X4 FILLER_82_672 ();
 FILLCELL_X2 FILLER_82_676 ();
 FILLCELL_X1 FILLER_82_678 ();
 FILLCELL_X2 FILLER_82_682 ();
 FILLCELL_X1 FILLER_82_684 ();
 FILLCELL_X16 FILLER_82_695 ();
 FILLCELL_X4 FILLER_82_711 ();
 FILLCELL_X2 FILLER_82_721 ();
 FILLCELL_X8 FILLER_82_748 ();
 FILLCELL_X2 FILLER_82_756 ();
 FILLCELL_X4 FILLER_82_762 ();
 FILLCELL_X1 FILLER_82_766 ();
 FILLCELL_X2 FILLER_82_771 ();
 FILLCELL_X1 FILLER_82_782 ();
 FILLCELL_X1 FILLER_82_792 ();
 FILLCELL_X1 FILLER_82_800 ();
 FILLCELL_X1 FILLER_82_806 ();
 FILLCELL_X8 FILLER_82_815 ();
 FILLCELL_X32 FILLER_82_827 ();
 FILLCELL_X32 FILLER_82_859 ();
 FILLCELL_X32 FILLER_82_891 ();
 FILLCELL_X32 FILLER_82_923 ();
 FILLCELL_X32 FILLER_82_955 ();
 FILLCELL_X32 FILLER_82_987 ();
 FILLCELL_X32 FILLER_82_1019 ();
 FILLCELL_X32 FILLER_82_1051 ();
 FILLCELL_X32 FILLER_82_1083 ();
 FILLCELL_X32 FILLER_82_1115 ();
 FILLCELL_X32 FILLER_82_1147 ();
 FILLCELL_X32 FILLER_82_1179 ();
 FILLCELL_X32 FILLER_82_1211 ();
 FILLCELL_X32 FILLER_82_1243 ();
 FILLCELL_X32 FILLER_82_1275 ();
 FILLCELL_X4 FILLER_82_1307 ();
 FILLCELL_X4 FILLER_82_1316 ();
 FILLCELL_X2 FILLER_82_1320 ();
 FILLCELL_X1 FILLER_82_1322 ();
 FILLCELL_X1 FILLER_83_7 ();
 FILLCELL_X8 FILLER_83_30 ();
 FILLCELL_X8 FILLER_83_40 ();
 FILLCELL_X1 FILLER_83_48 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X16 FILLER_83_161 ();
 FILLCELL_X2 FILLER_83_177 ();
 FILLCELL_X4 FILLER_83_187 ();
 FILLCELL_X2 FILLER_83_197 ();
 FILLCELL_X2 FILLER_83_208 ();
 FILLCELL_X1 FILLER_83_210 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X8 FILLER_83_609 ();
 FILLCELL_X1 FILLER_83_617 ();
 FILLCELL_X2 FILLER_83_622 ();
 FILLCELL_X32 FILLER_83_630 ();
 FILLCELL_X16 FILLER_83_662 ();
 FILLCELL_X2 FILLER_83_678 ();
 FILLCELL_X32 FILLER_83_684 ();
 FILLCELL_X8 FILLER_83_716 ();
 FILLCELL_X4 FILLER_83_724 ();
 FILLCELL_X2 FILLER_83_741 ();
 FILLCELL_X8 FILLER_83_748 ();
 FILLCELL_X4 FILLER_83_756 ();
 FILLCELL_X16 FILLER_83_781 ();
 FILLCELL_X4 FILLER_83_797 ();
 FILLCELL_X32 FILLER_83_831 ();
 FILLCELL_X32 FILLER_83_863 ();
 FILLCELL_X32 FILLER_83_895 ();
 FILLCELL_X32 FILLER_83_927 ();
 FILLCELL_X32 FILLER_83_959 ();
 FILLCELL_X32 FILLER_83_991 ();
 FILLCELL_X32 FILLER_83_1023 ();
 FILLCELL_X32 FILLER_83_1055 ();
 FILLCELL_X32 FILLER_83_1087 ();
 FILLCELL_X32 FILLER_83_1119 ();
 FILLCELL_X32 FILLER_83_1151 ();
 FILLCELL_X32 FILLER_83_1183 ();
 FILLCELL_X32 FILLER_83_1215 ();
 FILLCELL_X16 FILLER_83_1247 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X8 FILLER_83_1296 ();
 FILLCELL_X4 FILLER_83_1304 ();
 FILLCELL_X2 FILLER_83_1308 ();
 FILLCELL_X1 FILLER_83_1310 ();
 FILLCELL_X1 FILLER_83_1316 ();
 FILLCELL_X1 FILLER_83_1327 ();
 FILLCELL_X8 FILLER_84_1 ();
 FILLCELL_X2 FILLER_84_9 ();
 FILLCELL_X1 FILLER_84_11 ();
 FILLCELL_X2 FILLER_84_20 ();
 FILLCELL_X2 FILLER_84_50 ();
 FILLCELL_X1 FILLER_84_52 ();
 FILLCELL_X32 FILLER_84_61 ();
 FILLCELL_X1 FILLER_84_93 ();
 FILLCELL_X1 FILLER_84_98 ();
 FILLCELL_X32 FILLER_84_132 ();
 FILLCELL_X16 FILLER_84_164 ();
 FILLCELL_X4 FILLER_84_180 ();
 FILLCELL_X1 FILLER_84_184 ();
 FILLCELL_X1 FILLER_84_223 ();
 FILLCELL_X2 FILLER_84_230 ();
 FILLCELL_X32 FILLER_84_240 ();
 FILLCELL_X32 FILLER_84_272 ();
 FILLCELL_X16 FILLER_84_304 ();
 FILLCELL_X8 FILLER_84_320 ();
 FILLCELL_X2 FILLER_84_328 ();
 FILLCELL_X32 FILLER_84_337 ();
 FILLCELL_X32 FILLER_84_369 ();
 FILLCELL_X32 FILLER_84_401 ();
 FILLCELL_X32 FILLER_84_433 ();
 FILLCELL_X32 FILLER_84_465 ();
 FILLCELL_X32 FILLER_84_497 ();
 FILLCELL_X32 FILLER_84_529 ();
 FILLCELL_X8 FILLER_84_561 ();
 FILLCELL_X2 FILLER_84_569 ();
 FILLCELL_X1 FILLER_84_571 ();
 FILLCELL_X16 FILLER_84_576 ();
 FILLCELL_X4 FILLER_84_592 ();
 FILLCELL_X2 FILLER_84_596 ();
 FILLCELL_X1 FILLER_84_598 ();
 FILLCELL_X8 FILLER_84_619 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X2 FILLER_84_664 ();
 FILLCELL_X16 FILLER_84_687 ();
 FILLCELL_X4 FILLER_84_703 ();
 FILLCELL_X2 FILLER_84_707 ();
 FILLCELL_X32 FILLER_84_723 ();
 FILLCELL_X32 FILLER_84_755 ();
 FILLCELL_X32 FILLER_84_787 ();
 FILLCELL_X32 FILLER_84_819 ();
 FILLCELL_X32 FILLER_84_851 ();
 FILLCELL_X32 FILLER_84_883 ();
 FILLCELL_X32 FILLER_84_915 ();
 FILLCELL_X32 FILLER_84_947 ();
 FILLCELL_X32 FILLER_84_979 ();
 FILLCELL_X32 FILLER_84_1011 ();
 FILLCELL_X32 FILLER_84_1043 ();
 FILLCELL_X32 FILLER_84_1075 ();
 FILLCELL_X32 FILLER_84_1107 ();
 FILLCELL_X32 FILLER_84_1139 ();
 FILLCELL_X32 FILLER_84_1171 ();
 FILLCELL_X32 FILLER_84_1203 ();
 FILLCELL_X32 FILLER_84_1235 ();
 FILLCELL_X32 FILLER_84_1267 ();
 FILLCELL_X16 FILLER_84_1299 ();
 FILLCELL_X2 FILLER_84_1315 ();
 FILLCELL_X1 FILLER_84_1317 ();
 FILLCELL_X8 FILLER_85_1 ();
 FILLCELL_X4 FILLER_85_9 ();
 FILLCELL_X2 FILLER_85_13 ();
 FILLCELL_X1 FILLER_85_15 ();
 FILLCELL_X1 FILLER_85_19 ();
 FILLCELL_X2 FILLER_85_23 ();
 FILLCELL_X8 FILLER_85_39 ();
 FILLCELL_X4 FILLER_85_47 ();
 FILLCELL_X4 FILLER_85_65 ();
 FILLCELL_X2 FILLER_85_69 ();
 FILLCELL_X1 FILLER_85_71 ();
 FILLCELL_X8 FILLER_85_74 ();
 FILLCELL_X1 FILLER_85_107 ();
 FILLCELL_X2 FILLER_85_134 ();
 FILLCELL_X2 FILLER_85_140 ();
 FILLCELL_X16 FILLER_85_151 ();
 FILLCELL_X4 FILLER_85_167 ();
 FILLCELL_X2 FILLER_85_171 ();
 FILLCELL_X32 FILLER_85_177 ();
 FILLCELL_X8 FILLER_85_209 ();
 FILLCELL_X4 FILLER_85_217 ();
 FILLCELL_X1 FILLER_85_221 ();
 FILLCELL_X4 FILLER_85_226 ();
 FILLCELL_X2 FILLER_85_230 ();
 FILLCELL_X32 FILLER_85_253 ();
 FILLCELL_X32 FILLER_85_285 ();
 FILLCELL_X32 FILLER_85_317 ();
 FILLCELL_X32 FILLER_85_349 ();
 FILLCELL_X32 FILLER_85_381 ();
 FILLCELL_X32 FILLER_85_413 ();
 FILLCELL_X32 FILLER_85_445 ();
 FILLCELL_X32 FILLER_85_477 ();
 FILLCELL_X32 FILLER_85_509 ();
 FILLCELL_X32 FILLER_85_541 ();
 FILLCELL_X16 FILLER_85_573 ();
 FILLCELL_X8 FILLER_85_589 ();
 FILLCELL_X2 FILLER_85_597 ();
 FILLCELL_X2 FILLER_85_603 ();
 FILLCELL_X4 FILLER_85_622 ();
 FILLCELL_X2 FILLER_85_626 ();
 FILLCELL_X1 FILLER_85_628 ();
 FILLCELL_X16 FILLER_85_652 ();
 FILLCELL_X8 FILLER_85_668 ();
 FILLCELL_X4 FILLER_85_676 ();
 FILLCELL_X1 FILLER_85_680 ();
 FILLCELL_X16 FILLER_85_683 ();
 FILLCELL_X8 FILLER_85_699 ();
 FILLCELL_X4 FILLER_85_707 ();
 FILLCELL_X2 FILLER_85_711 ();
 FILLCELL_X1 FILLER_85_713 ();
 FILLCELL_X32 FILLER_85_738 ();
 FILLCELL_X16 FILLER_85_770 ();
 FILLCELL_X4 FILLER_85_786 ();
 FILLCELL_X1 FILLER_85_790 ();
 FILLCELL_X4 FILLER_85_796 ();
 FILLCELL_X2 FILLER_85_800 ();
 FILLCELL_X32 FILLER_85_806 ();
 FILLCELL_X32 FILLER_85_838 ();
 FILLCELL_X32 FILLER_85_870 ();
 FILLCELL_X32 FILLER_85_902 ();
 FILLCELL_X32 FILLER_85_934 ();
 FILLCELL_X32 FILLER_85_966 ();
 FILLCELL_X32 FILLER_85_998 ();
 FILLCELL_X32 FILLER_85_1030 ();
 FILLCELL_X32 FILLER_85_1062 ();
 FILLCELL_X32 FILLER_85_1094 ();
 FILLCELL_X32 FILLER_85_1126 ();
 FILLCELL_X32 FILLER_85_1158 ();
 FILLCELL_X32 FILLER_85_1190 ();
 FILLCELL_X32 FILLER_85_1222 ();
 FILLCELL_X8 FILLER_85_1254 ();
 FILLCELL_X1 FILLER_85_1262 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X8 FILLER_85_1296 ();
 FILLCELL_X4 FILLER_85_1304 ();
 FILLCELL_X2 FILLER_85_1308 ();
 FILLCELL_X1 FILLER_85_1310 ();
 FILLCELL_X1 FILLER_85_1316 ();
 FILLCELL_X1 FILLER_85_1327 ();
 FILLCELL_X4 FILLER_86_1 ();
 FILLCELL_X2 FILLER_86_5 ();
 FILLCELL_X4 FILLER_86_13 ();
 FILLCELL_X8 FILLER_86_26 ();
 FILLCELL_X2 FILLER_86_34 ();
 FILLCELL_X1 FILLER_86_36 ();
 FILLCELL_X32 FILLER_86_62 ();
 FILLCELL_X8 FILLER_86_94 ();
 FILLCELL_X4 FILLER_86_102 ();
 FILLCELL_X2 FILLER_86_106 ();
 FILLCELL_X1 FILLER_86_108 ();
 FILLCELL_X1 FILLER_86_124 ();
 FILLCELL_X8 FILLER_86_132 ();
 FILLCELL_X2 FILLER_86_140 ();
 FILLCELL_X1 FILLER_86_142 ();
 FILLCELL_X16 FILLER_86_151 ();
 FILLCELL_X16 FILLER_86_180 ();
 FILLCELL_X32 FILLER_86_201 ();
 FILLCELL_X32 FILLER_86_233 ();
 FILLCELL_X32 FILLER_86_265 ();
 FILLCELL_X32 FILLER_86_297 ();
 FILLCELL_X32 FILLER_86_329 ();
 FILLCELL_X32 FILLER_86_361 ();
 FILLCELL_X32 FILLER_86_393 ();
 FILLCELL_X32 FILLER_86_425 ();
 FILLCELL_X32 FILLER_86_457 ();
 FILLCELL_X32 FILLER_86_489 ();
 FILLCELL_X32 FILLER_86_521 ();
 FILLCELL_X32 FILLER_86_553 ();
 FILLCELL_X4 FILLER_86_585 ();
 FILLCELL_X2 FILLER_86_610 ();
 FILLCELL_X1 FILLER_86_612 ();
 FILLCELL_X16 FILLER_86_615 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X8 FILLER_86_664 ();
 FILLCELL_X2 FILLER_86_672 ();
 FILLCELL_X1 FILLER_86_674 ();
 FILLCELL_X32 FILLER_86_706 ();
 FILLCELL_X4 FILLER_86_738 ();
 FILLCELL_X2 FILLER_86_742 ();
 FILLCELL_X1 FILLER_86_744 ();
 FILLCELL_X16 FILLER_86_765 ();
 FILLCELL_X8 FILLER_86_781 ();
 FILLCELL_X4 FILLER_86_789 ();
 FILLCELL_X2 FILLER_86_793 ();
 FILLCELL_X2 FILLER_86_799 ();
 FILLCELL_X32 FILLER_86_805 ();
 FILLCELL_X32 FILLER_86_837 ();
 FILLCELL_X32 FILLER_86_869 ();
 FILLCELL_X32 FILLER_86_901 ();
 FILLCELL_X32 FILLER_86_933 ();
 FILLCELL_X32 FILLER_86_965 ();
 FILLCELL_X32 FILLER_86_997 ();
 FILLCELL_X32 FILLER_86_1029 ();
 FILLCELL_X32 FILLER_86_1061 ();
 FILLCELL_X32 FILLER_86_1093 ();
 FILLCELL_X32 FILLER_86_1125 ();
 FILLCELL_X32 FILLER_86_1157 ();
 FILLCELL_X32 FILLER_86_1189 ();
 FILLCELL_X32 FILLER_86_1221 ();
 FILLCELL_X32 FILLER_86_1253 ();
 FILLCELL_X16 FILLER_86_1285 ();
 FILLCELL_X8 FILLER_86_1301 ();
 FILLCELL_X4 FILLER_86_1309 ();
 FILLCELL_X1 FILLER_86_1313 ();
 FILLCELL_X2 FILLER_86_1319 ();
 FILLCELL_X2 FILLER_86_1326 ();
 FILLCELL_X2 FILLER_87_1 ();
 FILLCELL_X1 FILLER_87_3 ();
 FILLCELL_X4 FILLER_87_7 ();
 FILLCELL_X16 FILLER_87_14 ();
 FILLCELL_X2 FILLER_87_30 ();
 FILLCELL_X16 FILLER_87_35 ();
 FILLCELL_X16 FILLER_87_61 ();
 FILLCELL_X8 FILLER_87_77 ();
 FILLCELL_X4 FILLER_87_85 ();
 FILLCELL_X2 FILLER_87_89 ();
 FILLCELL_X1 FILLER_87_91 ();
 FILLCELL_X16 FILLER_87_95 ();
 FILLCELL_X2 FILLER_87_111 ();
 FILLCELL_X8 FILLER_87_126 ();
 FILLCELL_X2 FILLER_87_134 ();
 FILLCELL_X1 FILLER_87_136 ();
 FILLCELL_X2 FILLER_87_142 ();
 FILLCELL_X2 FILLER_87_166 ();
 FILLCELL_X1 FILLER_87_168 ();
 FILLCELL_X4 FILLER_87_191 ();
 FILLCELL_X1 FILLER_87_195 ();
 FILLCELL_X8 FILLER_87_205 ();
 FILLCELL_X4 FILLER_87_213 ();
 FILLCELL_X2 FILLER_87_217 ();
 FILLCELL_X8 FILLER_87_225 ();
 FILLCELL_X4 FILLER_87_233 ();
 FILLCELL_X1 FILLER_87_237 ();
 FILLCELL_X32 FILLER_87_240 ();
 FILLCELL_X32 FILLER_87_272 ();
 FILLCELL_X32 FILLER_87_304 ();
 FILLCELL_X32 FILLER_87_336 ();
 FILLCELL_X32 FILLER_87_368 ();
 FILLCELL_X32 FILLER_87_400 ();
 FILLCELL_X32 FILLER_87_432 ();
 FILLCELL_X32 FILLER_87_464 ();
 FILLCELL_X32 FILLER_87_496 ();
 FILLCELL_X32 FILLER_87_528 ();
 FILLCELL_X4 FILLER_87_560 ();
 FILLCELL_X1 FILLER_87_564 ();
 FILLCELL_X32 FILLER_87_569 ();
 FILLCELL_X16 FILLER_87_601 ();
 FILLCELL_X8 FILLER_87_617 ();
 FILLCELL_X16 FILLER_87_630 ();
 FILLCELL_X8 FILLER_87_646 ();
 FILLCELL_X4 FILLER_87_654 ();
 FILLCELL_X8 FILLER_87_665 ();
 FILLCELL_X1 FILLER_87_673 ();
 FILLCELL_X2 FILLER_87_678 ();
 FILLCELL_X4 FILLER_87_684 ();
 FILLCELL_X2 FILLER_87_697 ();
 FILLCELL_X1 FILLER_87_699 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X8 FILLER_87_737 ();
 FILLCELL_X4 FILLER_87_754 ();
 FILLCELL_X2 FILLER_87_758 ();
 FILLCELL_X4 FILLER_87_781 ();
 FILLCELL_X2 FILLER_87_785 ();
 FILLCELL_X32 FILLER_87_806 ();
 FILLCELL_X32 FILLER_87_838 ();
 FILLCELL_X32 FILLER_87_870 ();
 FILLCELL_X32 FILLER_87_902 ();
 FILLCELL_X32 FILLER_87_934 ();
 FILLCELL_X32 FILLER_87_966 ();
 FILLCELL_X32 FILLER_87_998 ();
 FILLCELL_X32 FILLER_87_1030 ();
 FILLCELL_X32 FILLER_87_1062 ();
 FILLCELL_X32 FILLER_87_1094 ();
 FILLCELL_X32 FILLER_87_1126 ();
 FILLCELL_X32 FILLER_87_1158 ();
 FILLCELL_X32 FILLER_87_1190 ();
 FILLCELL_X32 FILLER_87_1222 ();
 FILLCELL_X8 FILLER_87_1254 ();
 FILLCELL_X1 FILLER_87_1262 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X8 FILLER_87_1296 ();
 FILLCELL_X4 FILLER_87_1304 ();
 FILLCELL_X2 FILLER_87_1308 ();
 FILLCELL_X1 FILLER_87_1310 ();
 FILLCELL_X1 FILLER_87_1316 ();
 FILLCELL_X1 FILLER_87_1327 ();
 FILLCELL_X8 FILLER_88_1 ();
 FILLCELL_X2 FILLER_88_9 ();
 FILLCELL_X1 FILLER_88_11 ();
 FILLCELL_X2 FILLER_88_25 ();
 FILLCELL_X1 FILLER_88_27 ();
 FILLCELL_X32 FILLER_88_31 ();
 FILLCELL_X32 FILLER_88_63 ();
 FILLCELL_X32 FILLER_88_95 ();
 FILLCELL_X16 FILLER_88_127 ();
 FILLCELL_X4 FILLER_88_143 ();
 FILLCELL_X1 FILLER_88_147 ();
 FILLCELL_X32 FILLER_88_153 ();
 FILLCELL_X4 FILLER_88_185 ();
 FILLCELL_X1 FILLER_88_189 ();
 FILLCELL_X16 FILLER_88_217 ();
 FILLCELL_X32 FILLER_88_239 ();
 FILLCELL_X32 FILLER_88_271 ();
 FILLCELL_X32 FILLER_88_303 ();
 FILLCELL_X32 FILLER_88_335 ();
 FILLCELL_X32 FILLER_88_367 ();
 FILLCELL_X32 FILLER_88_399 ();
 FILLCELL_X32 FILLER_88_431 ();
 FILLCELL_X32 FILLER_88_463 ();
 FILLCELL_X32 FILLER_88_495 ();
 FILLCELL_X32 FILLER_88_527 ();
 FILLCELL_X32 FILLER_88_559 ();
 FILLCELL_X16 FILLER_88_591 ();
 FILLCELL_X4 FILLER_88_607 ();
 FILLCELL_X8 FILLER_88_632 ();
 FILLCELL_X1 FILLER_88_640 ();
 FILLCELL_X8 FILLER_88_658 ();
 FILLCELL_X4 FILLER_88_666 ();
 FILLCELL_X1 FILLER_88_670 ();
 FILLCELL_X2 FILLER_88_688 ();
 FILLCELL_X16 FILLER_88_698 ();
 FILLCELL_X8 FILLER_88_714 ();
 FILLCELL_X1 FILLER_88_722 ();
 FILLCELL_X8 FILLER_88_726 ();
 FILLCELL_X4 FILLER_88_734 ();
 FILLCELL_X4 FILLER_88_755 ();
 FILLCELL_X2 FILLER_88_759 ();
 FILLCELL_X16 FILLER_88_770 ();
 FILLCELL_X8 FILLER_88_786 ();
 FILLCELL_X2 FILLER_88_794 ();
 FILLCELL_X32 FILLER_88_800 ();
 FILLCELL_X32 FILLER_88_832 ();
 FILLCELL_X32 FILLER_88_864 ();
 FILLCELL_X32 FILLER_88_896 ();
 FILLCELL_X32 FILLER_88_928 ();
 FILLCELL_X32 FILLER_88_960 ();
 FILLCELL_X32 FILLER_88_992 ();
 FILLCELL_X32 FILLER_88_1024 ();
 FILLCELL_X32 FILLER_88_1056 ();
 FILLCELL_X32 FILLER_88_1088 ();
 FILLCELL_X32 FILLER_88_1120 ();
 FILLCELL_X32 FILLER_88_1152 ();
 FILLCELL_X32 FILLER_88_1184 ();
 FILLCELL_X32 FILLER_88_1216 ();
 FILLCELL_X32 FILLER_88_1248 ();
 FILLCELL_X32 FILLER_88_1280 ();
 FILLCELL_X4 FILLER_88_1312 ();
 FILLCELL_X1 FILLER_89_1 ();
 FILLCELL_X2 FILLER_89_5 ();
 FILLCELL_X1 FILLER_89_7 ();
 FILLCELL_X4 FILLER_89_26 ();
 FILLCELL_X2 FILLER_89_30 ();
 FILLCELL_X32 FILLER_89_35 ();
 FILLCELL_X8 FILLER_89_67 ();
 FILLCELL_X4 FILLER_89_75 ();
 FILLCELL_X2 FILLER_89_79 ();
 FILLCELL_X1 FILLER_89_81 ();
 FILLCELL_X2 FILLER_89_91 ();
 FILLCELL_X1 FILLER_89_93 ();
 FILLCELL_X1 FILLER_89_98 ();
 FILLCELL_X16 FILLER_89_103 ();
 FILLCELL_X4 FILLER_89_119 ();
 FILLCELL_X2 FILLER_89_123 ();
 FILLCELL_X1 FILLER_89_125 ();
 FILLCELL_X4 FILLER_89_130 ();
 FILLCELL_X1 FILLER_89_134 ();
 FILLCELL_X32 FILLER_89_145 ();
 FILLCELL_X2 FILLER_89_177 ();
 FILLCELL_X16 FILLER_89_200 ();
 FILLCELL_X2 FILLER_89_216 ();
 FILLCELL_X1 FILLER_89_229 ();
 FILLCELL_X32 FILLER_89_253 ();
 FILLCELL_X32 FILLER_89_285 ();
 FILLCELL_X32 FILLER_89_317 ();
 FILLCELL_X32 FILLER_89_349 ();
 FILLCELL_X32 FILLER_89_381 ();
 FILLCELL_X32 FILLER_89_413 ();
 FILLCELL_X32 FILLER_89_445 ();
 FILLCELL_X32 FILLER_89_477 ();
 FILLCELL_X32 FILLER_89_509 ();
 FILLCELL_X32 FILLER_89_541 ();
 FILLCELL_X32 FILLER_89_573 ();
 FILLCELL_X4 FILLER_89_605 ();
 FILLCELL_X1 FILLER_89_609 ();
 FILLCELL_X1 FILLER_89_618 ();
 FILLCELL_X32 FILLER_89_626 ();
 FILLCELL_X16 FILLER_89_658 ();
 FILLCELL_X4 FILLER_89_674 ();
 FILLCELL_X1 FILLER_89_678 ();
 FILLCELL_X16 FILLER_89_700 ();
 FILLCELL_X8 FILLER_89_716 ();
 FILLCELL_X8 FILLER_89_733 ();
 FILLCELL_X1 FILLER_89_745 ();
 FILLCELL_X16 FILLER_89_755 ();
 FILLCELL_X8 FILLER_89_771 ();
 FILLCELL_X2 FILLER_89_779 ();
 FILLCELL_X1 FILLER_89_781 ();
 FILLCELL_X32 FILLER_89_802 ();
 FILLCELL_X32 FILLER_89_834 ();
 FILLCELL_X32 FILLER_89_866 ();
 FILLCELL_X32 FILLER_89_898 ();
 FILLCELL_X32 FILLER_89_930 ();
 FILLCELL_X32 FILLER_89_962 ();
 FILLCELL_X32 FILLER_89_994 ();
 FILLCELL_X32 FILLER_89_1026 ();
 FILLCELL_X32 FILLER_89_1058 ();
 FILLCELL_X32 FILLER_89_1090 ();
 FILLCELL_X32 FILLER_89_1122 ();
 FILLCELL_X32 FILLER_89_1154 ();
 FILLCELL_X32 FILLER_89_1186 ();
 FILLCELL_X32 FILLER_89_1218 ();
 FILLCELL_X8 FILLER_89_1250 ();
 FILLCELL_X4 FILLER_89_1258 ();
 FILLCELL_X1 FILLER_89_1262 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X16 FILLER_89_1296 ();
 FILLCELL_X2 FILLER_89_1312 ();
 FILLCELL_X1 FILLER_89_1321 ();
 FILLCELL_X2 FILLER_90_1 ();
 FILLCELL_X2 FILLER_90_30 ();
 FILLCELL_X1 FILLER_90_32 ();
 FILLCELL_X8 FILLER_90_43 ();
 FILLCELL_X4 FILLER_90_51 ();
 FILLCELL_X2 FILLER_90_55 ();
 FILLCELL_X1 FILLER_90_61 ();
 FILLCELL_X2 FILLER_90_70 ();
 FILLCELL_X1 FILLER_90_88 ();
 FILLCELL_X4 FILLER_90_92 ();
 FILLCELL_X2 FILLER_90_96 ();
 FILLCELL_X1 FILLER_90_98 ();
 FILLCELL_X16 FILLER_90_104 ();
 FILLCELL_X2 FILLER_90_120 ();
 FILLCELL_X1 FILLER_90_122 ();
 FILLCELL_X2 FILLER_90_130 ();
 FILLCELL_X1 FILLER_90_144 ();
 FILLCELL_X32 FILLER_90_156 ();
 FILLCELL_X16 FILLER_90_188 ();
 FILLCELL_X4 FILLER_90_204 ();
 FILLCELL_X1 FILLER_90_214 ();
 FILLCELL_X32 FILLER_90_263 ();
 FILLCELL_X32 FILLER_90_295 ();
 FILLCELL_X32 FILLER_90_327 ();
 FILLCELL_X32 FILLER_90_359 ();
 FILLCELL_X32 FILLER_90_391 ();
 FILLCELL_X32 FILLER_90_423 ();
 FILLCELL_X32 FILLER_90_455 ();
 FILLCELL_X32 FILLER_90_487 ();
 FILLCELL_X32 FILLER_90_519 ();
 FILLCELL_X32 FILLER_90_551 ();
 FILLCELL_X8 FILLER_90_583 ();
 FILLCELL_X2 FILLER_90_591 ();
 FILLCELL_X4 FILLER_90_610 ();
 FILLCELL_X1 FILLER_90_614 ();
 FILLCELL_X8 FILLER_90_622 ();
 FILLCELL_X1 FILLER_90_630 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X8 FILLER_90_696 ();
 FILLCELL_X1 FILLER_90_736 ();
 FILLCELL_X4 FILLER_90_758 ();
 FILLCELL_X2 FILLER_90_762 ();
 FILLCELL_X16 FILLER_90_768 ();
 FILLCELL_X8 FILLER_90_784 ();
 FILLCELL_X4 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_816 ();
 FILLCELL_X32 FILLER_90_848 ();
 FILLCELL_X32 FILLER_90_880 ();
 FILLCELL_X32 FILLER_90_912 ();
 FILLCELL_X32 FILLER_90_944 ();
 FILLCELL_X32 FILLER_90_976 ();
 FILLCELL_X32 FILLER_90_1008 ();
 FILLCELL_X32 FILLER_90_1040 ();
 FILLCELL_X32 FILLER_90_1072 ();
 FILLCELL_X32 FILLER_90_1104 ();
 FILLCELL_X32 FILLER_90_1136 ();
 FILLCELL_X32 FILLER_90_1168 ();
 FILLCELL_X32 FILLER_90_1200 ();
 FILLCELL_X32 FILLER_90_1232 ();
 FILLCELL_X32 FILLER_90_1264 ();
 FILLCELL_X8 FILLER_90_1296 ();
 FILLCELL_X4 FILLER_90_1304 ();
 FILLCELL_X2 FILLER_90_1308 ();
 FILLCELL_X1 FILLER_90_1310 ();
 FILLCELL_X2 FILLER_90_1313 ();
 FILLCELL_X1 FILLER_90_1315 ();
 FILLCELL_X2 FILLER_90_1318 ();
 FILLCELL_X1 FILLER_90_1320 ();
 FILLCELL_X1 FILLER_90_1327 ();
 FILLCELL_X16 FILLER_91_1 ();
 FILLCELL_X1 FILLER_91_17 ();
 FILLCELL_X16 FILLER_91_28 ();
 FILLCELL_X4 FILLER_91_44 ();
 FILLCELL_X2 FILLER_91_67 ();
 FILLCELL_X1 FILLER_91_69 ();
 FILLCELL_X2 FILLER_91_74 ();
 FILLCELL_X16 FILLER_91_94 ();
 FILLCELL_X8 FILLER_91_110 ();
 FILLCELL_X2 FILLER_91_118 ();
 FILLCELL_X1 FILLER_91_130 ();
 FILLCELL_X16 FILLER_91_141 ();
 FILLCELL_X16 FILLER_91_182 ();
 FILLCELL_X8 FILLER_91_198 ();
 FILLCELL_X32 FILLER_91_223 ();
 FILLCELL_X4 FILLER_91_255 ();
 FILLCELL_X1 FILLER_91_259 ();
 FILLCELL_X4 FILLER_91_268 ();
 FILLCELL_X2 FILLER_91_272 ();
 FILLCELL_X32 FILLER_91_293 ();
 FILLCELL_X32 FILLER_91_325 ();
 FILLCELL_X32 FILLER_91_357 ();
 FILLCELL_X32 FILLER_91_389 ();
 FILLCELL_X32 FILLER_91_421 ();
 FILLCELL_X32 FILLER_91_453 ();
 FILLCELL_X32 FILLER_91_485 ();
 FILLCELL_X32 FILLER_91_517 ();
 FILLCELL_X32 FILLER_91_549 ();
 FILLCELL_X16 FILLER_91_581 ();
 FILLCELL_X8 FILLER_91_600 ();
 FILLCELL_X4 FILLER_91_608 ();
 FILLCELL_X1 FILLER_91_612 ();
 FILLCELL_X32 FILLER_91_620 ();
 FILLCELL_X32 FILLER_91_652 ();
 FILLCELL_X32 FILLER_91_684 ();
 FILLCELL_X8 FILLER_91_720 ();
 FILLCELL_X4 FILLER_91_728 ();
 FILLCELL_X2 FILLER_91_732 ();
 FILLCELL_X8 FILLER_91_738 ();
 FILLCELL_X4 FILLER_91_746 ();
 FILLCELL_X2 FILLER_91_750 ();
 FILLCELL_X1 FILLER_91_752 ();
 FILLCELL_X32 FILLER_91_757 ();
 FILLCELL_X4 FILLER_91_789 ();
 FILLCELL_X2 FILLER_91_793 ();
 FILLCELL_X1 FILLER_91_795 ();
 FILLCELL_X32 FILLER_91_810 ();
 FILLCELL_X32 FILLER_91_842 ();
 FILLCELL_X32 FILLER_91_874 ();
 FILLCELL_X32 FILLER_91_906 ();
 FILLCELL_X32 FILLER_91_938 ();
 FILLCELL_X32 FILLER_91_970 ();
 FILLCELL_X32 FILLER_91_1002 ();
 FILLCELL_X32 FILLER_91_1034 ();
 FILLCELL_X32 FILLER_91_1066 ();
 FILLCELL_X32 FILLER_91_1098 ();
 FILLCELL_X32 FILLER_91_1130 ();
 FILLCELL_X32 FILLER_91_1162 ();
 FILLCELL_X32 FILLER_91_1194 ();
 FILLCELL_X32 FILLER_91_1226 ();
 FILLCELL_X4 FILLER_91_1258 ();
 FILLCELL_X1 FILLER_91_1262 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X8 FILLER_91_1296 ();
 FILLCELL_X4 FILLER_91_1304 ();
 FILLCELL_X2 FILLER_91_1308 ();
 FILLCELL_X1 FILLER_91_1310 ();
 FILLCELL_X2 FILLER_91_1316 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X16 FILLER_92_33 ();
 FILLCELL_X8 FILLER_92_49 ();
 FILLCELL_X4 FILLER_92_57 ();
 FILLCELL_X2 FILLER_92_61 ();
 FILLCELL_X2 FILLER_92_67 ();
 FILLCELL_X4 FILLER_92_78 ();
 FILLCELL_X2 FILLER_92_92 ();
 FILLCELL_X16 FILLER_92_106 ();
 FILLCELL_X8 FILLER_92_122 ();
 FILLCELL_X32 FILLER_92_150 ();
 FILLCELL_X32 FILLER_92_182 ();
 FILLCELL_X32 FILLER_92_214 ();
 FILLCELL_X8 FILLER_92_246 ();
 FILLCELL_X4 FILLER_92_254 ();
 FILLCELL_X2 FILLER_92_258 ();
 FILLCELL_X32 FILLER_92_286 ();
 FILLCELL_X32 FILLER_92_318 ();
 FILLCELL_X32 FILLER_92_350 ();
 FILLCELL_X32 FILLER_92_382 ();
 FILLCELL_X32 FILLER_92_414 ();
 FILLCELL_X32 FILLER_92_446 ();
 FILLCELL_X32 FILLER_92_478 ();
 FILLCELL_X32 FILLER_92_510 ();
 FILLCELL_X32 FILLER_92_542 ();
 FILLCELL_X32 FILLER_92_574 ();
 FILLCELL_X8 FILLER_92_606 ();
 FILLCELL_X2 FILLER_92_614 ();
 FILLCELL_X1 FILLER_92_616 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X2 FILLER_92_728 ();
 FILLCELL_X1 FILLER_92_730 ();
 FILLCELL_X32 FILLER_92_767 ();
 FILLCELL_X32 FILLER_92_799 ();
 FILLCELL_X32 FILLER_92_831 ();
 FILLCELL_X32 FILLER_92_863 ();
 FILLCELL_X32 FILLER_92_895 ();
 FILLCELL_X32 FILLER_92_927 ();
 FILLCELL_X32 FILLER_92_959 ();
 FILLCELL_X32 FILLER_92_991 ();
 FILLCELL_X32 FILLER_92_1023 ();
 FILLCELL_X32 FILLER_92_1055 ();
 FILLCELL_X32 FILLER_92_1087 ();
 FILLCELL_X32 FILLER_92_1119 ();
 FILLCELL_X32 FILLER_92_1151 ();
 FILLCELL_X32 FILLER_92_1183 ();
 FILLCELL_X32 FILLER_92_1215 ();
 FILLCELL_X32 FILLER_92_1247 ();
 FILLCELL_X32 FILLER_92_1279 ();
 FILLCELL_X4 FILLER_92_1311 ();
 FILLCELL_X1 FILLER_92_1315 ();
 FILLCELL_X2 FILLER_92_1326 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X16 FILLER_93_33 ();
 FILLCELL_X8 FILLER_93_49 ();
 FILLCELL_X2 FILLER_93_57 ();
 FILLCELL_X8 FILLER_93_82 ();
 FILLCELL_X2 FILLER_93_90 ();
 FILLCELL_X8 FILLER_93_95 ();
 FILLCELL_X16 FILLER_93_110 ();
 FILLCELL_X8 FILLER_93_126 ();
 FILLCELL_X1 FILLER_93_134 ();
 FILLCELL_X1 FILLER_93_139 ();
 FILLCELL_X4 FILLER_93_145 ();
 FILLCELL_X32 FILLER_93_153 ();
 FILLCELL_X32 FILLER_93_185 ();
 FILLCELL_X32 FILLER_93_217 ();
 FILLCELL_X32 FILLER_93_249 ();
 FILLCELL_X32 FILLER_93_281 ();
 FILLCELL_X32 FILLER_93_313 ();
 FILLCELL_X32 FILLER_93_345 ();
 FILLCELL_X32 FILLER_93_377 ();
 FILLCELL_X32 FILLER_93_409 ();
 FILLCELL_X32 FILLER_93_441 ();
 FILLCELL_X32 FILLER_93_473 ();
 FILLCELL_X32 FILLER_93_505 ();
 FILLCELL_X32 FILLER_93_537 ();
 FILLCELL_X32 FILLER_93_569 ();
 FILLCELL_X8 FILLER_93_601 ();
 FILLCELL_X4 FILLER_93_609 ();
 FILLCELL_X2 FILLER_93_613 ();
 FILLCELL_X1 FILLER_93_615 ();
 FILLCELL_X4 FILLER_93_619 ();
 FILLCELL_X2 FILLER_93_623 ();
 FILLCELL_X1 FILLER_93_625 ();
 FILLCELL_X32 FILLER_93_640 ();
 FILLCELL_X32 FILLER_93_672 ();
 FILLCELL_X32 FILLER_93_704 ();
 FILLCELL_X32 FILLER_93_736 ();
 FILLCELL_X32 FILLER_93_768 ();
 FILLCELL_X32 FILLER_93_800 ();
 FILLCELL_X32 FILLER_93_832 ();
 FILLCELL_X32 FILLER_93_864 ();
 FILLCELL_X32 FILLER_93_896 ();
 FILLCELL_X32 FILLER_93_928 ();
 FILLCELL_X32 FILLER_93_960 ();
 FILLCELL_X32 FILLER_93_992 ();
 FILLCELL_X32 FILLER_93_1024 ();
 FILLCELL_X32 FILLER_93_1056 ();
 FILLCELL_X32 FILLER_93_1088 ();
 FILLCELL_X32 FILLER_93_1120 ();
 FILLCELL_X32 FILLER_93_1152 ();
 FILLCELL_X32 FILLER_93_1184 ();
 FILLCELL_X32 FILLER_93_1216 ();
 FILLCELL_X8 FILLER_93_1248 ();
 FILLCELL_X4 FILLER_93_1256 ();
 FILLCELL_X2 FILLER_93_1260 ();
 FILLCELL_X1 FILLER_93_1262 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X8 FILLER_93_1296 ();
 FILLCELL_X4 FILLER_93_1304 ();
 FILLCELL_X2 FILLER_93_1308 ();
 FILLCELL_X1 FILLER_93_1310 ();
 FILLCELL_X1 FILLER_93_1316 ();
 FILLCELL_X1 FILLER_93_1324 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X8 FILLER_94_65 ();
 FILLCELL_X4 FILLER_94_73 ();
 FILLCELL_X1 FILLER_94_77 ();
 FILLCELL_X4 FILLER_94_95 ();
 FILLCELL_X2 FILLER_94_99 ();
 FILLCELL_X8 FILLER_94_108 ();
 FILLCELL_X2 FILLER_94_116 ();
 FILLCELL_X1 FILLER_94_118 ();
 FILLCELL_X4 FILLER_94_136 ();
 FILLCELL_X2 FILLER_94_140 ();
 FILLCELL_X32 FILLER_94_145 ();
 FILLCELL_X16 FILLER_94_177 ();
 FILLCELL_X8 FILLER_94_193 ();
 FILLCELL_X2 FILLER_94_201 ();
 FILLCELL_X1 FILLER_94_203 ();
 FILLCELL_X32 FILLER_94_214 ();
 FILLCELL_X32 FILLER_94_246 ();
 FILLCELL_X32 FILLER_94_278 ();
 FILLCELL_X32 FILLER_94_310 ();
 FILLCELL_X32 FILLER_94_342 ();
 FILLCELL_X32 FILLER_94_374 ();
 FILLCELL_X32 FILLER_94_406 ();
 FILLCELL_X32 FILLER_94_438 ();
 FILLCELL_X32 FILLER_94_470 ();
 FILLCELL_X32 FILLER_94_502 ();
 FILLCELL_X32 FILLER_94_534 ();
 FILLCELL_X32 FILLER_94_566 ();
 FILLCELL_X16 FILLER_94_598 ();
 FILLCELL_X4 FILLER_94_614 ();
 FILLCELL_X1 FILLER_94_618 ();
 FILLCELL_X8 FILLER_94_635 ();
 FILLCELL_X4 FILLER_94_643 ();
 FILLCELL_X2 FILLER_94_647 ();
 FILLCELL_X1 FILLER_94_649 ();
 FILLCELL_X32 FILLER_94_654 ();
 FILLCELL_X32 FILLER_94_686 ();
 FILLCELL_X32 FILLER_94_718 ();
 FILLCELL_X32 FILLER_94_750 ();
 FILLCELL_X32 FILLER_94_782 ();
 FILLCELL_X32 FILLER_94_814 ();
 FILLCELL_X32 FILLER_94_846 ();
 FILLCELL_X32 FILLER_94_878 ();
 FILLCELL_X32 FILLER_94_910 ();
 FILLCELL_X32 FILLER_94_942 ();
 FILLCELL_X32 FILLER_94_974 ();
 FILLCELL_X32 FILLER_94_1006 ();
 FILLCELL_X32 FILLER_94_1038 ();
 FILLCELL_X32 FILLER_94_1070 ();
 FILLCELL_X32 FILLER_94_1102 ();
 FILLCELL_X32 FILLER_94_1134 ();
 FILLCELL_X32 FILLER_94_1166 ();
 FILLCELL_X32 FILLER_94_1198 ();
 FILLCELL_X32 FILLER_94_1230 ();
 FILLCELL_X32 FILLER_94_1262 ();
 FILLCELL_X16 FILLER_94_1294 ();
 FILLCELL_X4 FILLER_94_1310 ();
 FILLCELL_X2 FILLER_94_1316 ();
 FILLCELL_X1 FILLER_94_1318 ();
 FILLCELL_X1 FILLER_94_1324 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X16 FILLER_95_65 ();
 FILLCELL_X4 FILLER_95_81 ();
 FILLCELL_X2 FILLER_95_85 ();
 FILLCELL_X1 FILLER_95_87 ();
 FILLCELL_X32 FILLER_95_105 ();
 FILLCELL_X1 FILLER_95_137 ();
 FILLCELL_X32 FILLER_95_155 ();
 FILLCELL_X8 FILLER_95_187 ();
 FILLCELL_X4 FILLER_95_195 ();
 FILLCELL_X2 FILLER_95_199 ();
 FILLCELL_X1 FILLER_95_201 ();
 FILLCELL_X32 FILLER_95_216 ();
 FILLCELL_X32 FILLER_95_248 ();
 FILLCELL_X32 FILLER_95_280 ();
 FILLCELL_X32 FILLER_95_312 ();
 FILLCELL_X32 FILLER_95_344 ();
 FILLCELL_X32 FILLER_95_376 ();
 FILLCELL_X32 FILLER_95_408 ();
 FILLCELL_X32 FILLER_95_440 ();
 FILLCELL_X32 FILLER_95_472 ();
 FILLCELL_X32 FILLER_95_504 ();
 FILLCELL_X32 FILLER_95_536 ();
 FILLCELL_X32 FILLER_95_568 ();
 FILLCELL_X16 FILLER_95_600 ();
 FILLCELL_X8 FILLER_95_616 ();
 FILLCELL_X32 FILLER_95_643 ();
 FILLCELL_X32 FILLER_95_675 ();
 FILLCELL_X32 FILLER_95_707 ();
 FILLCELL_X32 FILLER_95_739 ();
 FILLCELL_X32 FILLER_95_771 ();
 FILLCELL_X32 FILLER_95_803 ();
 FILLCELL_X32 FILLER_95_835 ();
 FILLCELL_X32 FILLER_95_867 ();
 FILLCELL_X32 FILLER_95_899 ();
 FILLCELL_X32 FILLER_95_931 ();
 FILLCELL_X32 FILLER_95_963 ();
 FILLCELL_X32 FILLER_95_995 ();
 FILLCELL_X32 FILLER_95_1027 ();
 FILLCELL_X32 FILLER_95_1059 ();
 FILLCELL_X32 FILLER_95_1091 ();
 FILLCELL_X32 FILLER_95_1123 ();
 FILLCELL_X32 FILLER_95_1155 ();
 FILLCELL_X32 FILLER_95_1187 ();
 FILLCELL_X32 FILLER_95_1219 ();
 FILLCELL_X8 FILLER_95_1251 ();
 FILLCELL_X4 FILLER_95_1259 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X16 FILLER_95_1296 ();
 FILLCELL_X4 FILLER_95_1312 ();
 FILLCELL_X1 FILLER_95_1316 ();
 FILLCELL_X1 FILLER_95_1319 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X2 FILLER_96_609 ();
 FILLCELL_X1 FILLER_96_611 ();
 FILLCELL_X16 FILLER_96_632 ();
 FILLCELL_X8 FILLER_96_648 ();
 FILLCELL_X4 FILLER_96_656 ();
 FILLCELL_X32 FILLER_96_667 ();
 FILLCELL_X32 FILLER_96_699 ();
 FILLCELL_X32 FILLER_96_731 ();
 FILLCELL_X32 FILLER_96_763 ();
 FILLCELL_X32 FILLER_96_795 ();
 FILLCELL_X32 FILLER_96_827 ();
 FILLCELL_X32 FILLER_96_859 ();
 FILLCELL_X32 FILLER_96_891 ();
 FILLCELL_X32 FILLER_96_923 ();
 FILLCELL_X32 FILLER_96_955 ();
 FILLCELL_X32 FILLER_96_987 ();
 FILLCELL_X32 FILLER_96_1019 ();
 FILLCELL_X32 FILLER_96_1051 ();
 FILLCELL_X32 FILLER_96_1083 ();
 FILLCELL_X32 FILLER_96_1115 ();
 FILLCELL_X32 FILLER_96_1147 ();
 FILLCELL_X32 FILLER_96_1179 ();
 FILLCELL_X32 FILLER_96_1211 ();
 FILLCELL_X32 FILLER_96_1243 ();
 FILLCELL_X32 FILLER_96_1275 ();
 FILLCELL_X4 FILLER_96_1307 ();
 FILLCELL_X2 FILLER_96_1321 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X16 FILLER_97_161 ();
 FILLCELL_X2 FILLER_97_177 ();
 FILLCELL_X32 FILLER_97_188 ();
 FILLCELL_X32 FILLER_97_220 ();
 FILLCELL_X32 FILLER_97_252 ();
 FILLCELL_X32 FILLER_97_284 ();
 FILLCELL_X32 FILLER_97_316 ();
 FILLCELL_X32 FILLER_97_348 ();
 FILLCELL_X32 FILLER_97_380 ();
 FILLCELL_X32 FILLER_97_412 ();
 FILLCELL_X32 FILLER_97_444 ();
 FILLCELL_X32 FILLER_97_476 ();
 FILLCELL_X32 FILLER_97_508 ();
 FILLCELL_X32 FILLER_97_540 ();
 FILLCELL_X32 FILLER_97_572 ();
 FILLCELL_X32 FILLER_97_604 ();
 FILLCELL_X32 FILLER_97_636 ();
 FILLCELL_X32 FILLER_97_668 ();
 FILLCELL_X32 FILLER_97_700 ();
 FILLCELL_X32 FILLER_97_732 ();
 FILLCELL_X32 FILLER_97_764 ();
 FILLCELL_X32 FILLER_97_796 ();
 FILLCELL_X32 FILLER_97_828 ();
 FILLCELL_X32 FILLER_97_860 ();
 FILLCELL_X32 FILLER_97_892 ();
 FILLCELL_X32 FILLER_97_924 ();
 FILLCELL_X32 FILLER_97_956 ();
 FILLCELL_X32 FILLER_97_988 ();
 FILLCELL_X32 FILLER_97_1020 ();
 FILLCELL_X32 FILLER_97_1052 ();
 FILLCELL_X32 FILLER_97_1084 ();
 FILLCELL_X32 FILLER_97_1116 ();
 FILLCELL_X32 FILLER_97_1148 ();
 FILLCELL_X32 FILLER_97_1180 ();
 FILLCELL_X32 FILLER_97_1212 ();
 FILLCELL_X16 FILLER_97_1244 ();
 FILLCELL_X2 FILLER_97_1260 ();
 FILLCELL_X1 FILLER_97_1262 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X8 FILLER_97_1296 ();
 FILLCELL_X4 FILLER_97_1304 ();
 FILLCELL_X2 FILLER_97_1308 ();
 FILLCELL_X1 FILLER_97_1310 ();
 FILLCELL_X2 FILLER_97_1313 ();
 FILLCELL_X1 FILLER_97_1315 ();
 FILLCELL_X1 FILLER_97_1324 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X8 FILLER_98_161 ();
 FILLCELL_X4 FILLER_98_169 ();
 FILLCELL_X2 FILLER_98_173 ();
 FILLCELL_X32 FILLER_98_194 ();
 FILLCELL_X32 FILLER_98_226 ();
 FILLCELL_X32 FILLER_98_258 ();
 FILLCELL_X32 FILLER_98_290 ();
 FILLCELL_X32 FILLER_98_322 ();
 FILLCELL_X32 FILLER_98_354 ();
 FILLCELL_X32 FILLER_98_386 ();
 FILLCELL_X32 FILLER_98_418 ();
 FILLCELL_X32 FILLER_98_450 ();
 FILLCELL_X32 FILLER_98_482 ();
 FILLCELL_X32 FILLER_98_514 ();
 FILLCELL_X32 FILLER_98_546 ();
 FILLCELL_X32 FILLER_98_578 ();
 FILLCELL_X16 FILLER_98_610 ();
 FILLCELL_X4 FILLER_98_626 ();
 FILLCELL_X1 FILLER_98_630 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X8 FILLER_98_1304 ();
 FILLCELL_X2 FILLER_98_1312 ();
 FILLCELL_X1 FILLER_98_1319 ();
 FILLCELL_X1 FILLER_98_1327 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X8 FILLER_99_1296 ();
 FILLCELL_X4 FILLER_99_1304 ();
 FILLCELL_X2 FILLER_99_1308 ();
 FILLCELL_X1 FILLER_99_1310 ();
 FILLCELL_X1 FILLER_99_1318 ();
 FILLCELL_X1 FILLER_99_1324 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X16 FILLER_100_696 ();
 FILLCELL_X4 FILLER_100_712 ();
 FILLCELL_X2 FILLER_100_716 ();
 FILLCELL_X32 FILLER_100_732 ();
 FILLCELL_X32 FILLER_100_764 ();
 FILLCELL_X32 FILLER_100_796 ();
 FILLCELL_X32 FILLER_100_828 ();
 FILLCELL_X32 FILLER_100_860 ();
 FILLCELL_X32 FILLER_100_892 ();
 FILLCELL_X32 FILLER_100_924 ();
 FILLCELL_X32 FILLER_100_956 ();
 FILLCELL_X32 FILLER_100_988 ();
 FILLCELL_X32 FILLER_100_1020 ();
 FILLCELL_X32 FILLER_100_1052 ();
 FILLCELL_X32 FILLER_100_1084 ();
 FILLCELL_X32 FILLER_100_1116 ();
 FILLCELL_X32 FILLER_100_1148 ();
 FILLCELL_X32 FILLER_100_1180 ();
 FILLCELL_X32 FILLER_100_1212 ();
 FILLCELL_X32 FILLER_100_1244 ();
 FILLCELL_X32 FILLER_100_1276 ();
 FILLCELL_X8 FILLER_100_1308 ();
 FILLCELL_X2 FILLER_100_1321 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X8 FILLER_101_1296 ();
 FILLCELL_X4 FILLER_101_1304 ();
 FILLCELL_X2 FILLER_101_1308 ();
 FILLCELL_X1 FILLER_101_1310 ();
 FILLCELL_X1 FILLER_101_1316 ();
 FILLCELL_X1 FILLER_101_1327 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X8 FILLER_102_1304 ();
 FILLCELL_X4 FILLER_102_1312 ();
 FILLCELL_X1 FILLER_102_1323 ();
 FILLCELL_X1 FILLER_102_1327 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X8 FILLER_103_1296 ();
 FILLCELL_X4 FILLER_103_1304 ();
 FILLCELL_X2 FILLER_103_1308 ();
 FILLCELL_X1 FILLER_103_1310 ();
 FILLCELL_X2 FILLER_103_1318 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X4 FILLER_104_1304 ();
 FILLCELL_X2 FILLER_104_1308 ();
 FILLCELL_X1 FILLER_104_1310 ();
 FILLCELL_X2 FILLER_104_1313 ();
 FILLCELL_X1 FILLER_104_1315 ();
 FILLCELL_X4 FILLER_104_1319 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X32 FILLER_105_961 ();
 FILLCELL_X32 FILLER_105_993 ();
 FILLCELL_X32 FILLER_105_1025 ();
 FILLCELL_X32 FILLER_105_1057 ();
 FILLCELL_X32 FILLER_105_1089 ();
 FILLCELL_X32 FILLER_105_1121 ();
 FILLCELL_X32 FILLER_105_1153 ();
 FILLCELL_X32 FILLER_105_1185 ();
 FILLCELL_X32 FILLER_105_1217 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X8 FILLER_105_1296 ();
 FILLCELL_X4 FILLER_105_1304 ();
 FILLCELL_X2 FILLER_105_1308 ();
 FILLCELL_X1 FILLER_105_1310 ();
 FILLCELL_X1 FILLER_105_1313 ();
 FILLCELL_X1 FILLER_105_1324 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X8 FILLER_106_1304 ();
 FILLCELL_X4 FILLER_106_1312 ();
 FILLCELL_X2 FILLER_106_1321 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X32 FILLER_107_961 ();
 FILLCELL_X32 FILLER_107_993 ();
 FILLCELL_X32 FILLER_107_1025 ();
 FILLCELL_X32 FILLER_107_1057 ();
 FILLCELL_X32 FILLER_107_1089 ();
 FILLCELL_X32 FILLER_107_1121 ();
 FILLCELL_X32 FILLER_107_1153 ();
 FILLCELL_X32 FILLER_107_1185 ();
 FILLCELL_X32 FILLER_107_1217 ();
 FILLCELL_X8 FILLER_107_1249 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X8 FILLER_107_1296 ();
 FILLCELL_X4 FILLER_107_1304 ();
 FILLCELL_X2 FILLER_107_1308 ();
 FILLCELL_X1 FILLER_107_1310 ();
 FILLCELL_X2 FILLER_107_1313 ();
 FILLCELL_X1 FILLER_107_1315 ();
 FILLCELL_X1 FILLER_107_1324 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X16 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_751 ();
 FILLCELL_X32 FILLER_108_783 ();
 FILLCELL_X32 FILLER_108_815 ();
 FILLCELL_X32 FILLER_108_847 ();
 FILLCELL_X32 FILLER_108_879 ();
 FILLCELL_X32 FILLER_108_911 ();
 FILLCELL_X32 FILLER_108_943 ();
 FILLCELL_X32 FILLER_108_975 ();
 FILLCELL_X32 FILLER_108_1007 ();
 FILLCELL_X32 FILLER_108_1039 ();
 FILLCELL_X32 FILLER_108_1071 ();
 FILLCELL_X32 FILLER_108_1103 ();
 FILLCELL_X32 FILLER_108_1135 ();
 FILLCELL_X32 FILLER_108_1167 ();
 FILLCELL_X32 FILLER_108_1199 ();
 FILLCELL_X32 FILLER_108_1231 ();
 FILLCELL_X32 FILLER_108_1263 ();
 FILLCELL_X16 FILLER_108_1295 ();
 FILLCELL_X2 FILLER_108_1311 ();
 FILLCELL_X1 FILLER_108_1313 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X16 FILLER_109_1296 ();
 FILLCELL_X1 FILLER_109_1312 ();
 FILLCELL_X1 FILLER_109_1315 ();
 FILLCELL_X1 FILLER_109_1327 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X32 FILLER_110_952 ();
 FILLCELL_X32 FILLER_110_984 ();
 FILLCELL_X32 FILLER_110_1016 ();
 FILLCELL_X32 FILLER_110_1048 ();
 FILLCELL_X32 FILLER_110_1080 ();
 FILLCELL_X32 FILLER_110_1112 ();
 FILLCELL_X32 FILLER_110_1144 ();
 FILLCELL_X32 FILLER_110_1176 ();
 FILLCELL_X32 FILLER_110_1208 ();
 FILLCELL_X32 FILLER_110_1240 ();
 FILLCELL_X32 FILLER_110_1272 ();
 FILLCELL_X8 FILLER_110_1304 ();
 FILLCELL_X1 FILLER_110_1312 ();
 FILLCELL_X4 FILLER_110_1316 ();
 FILLCELL_X2 FILLER_110_1320 ();
 FILLCELL_X1 FILLER_110_1322 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X32 FILLER_111_961 ();
 FILLCELL_X32 FILLER_111_993 ();
 FILLCELL_X32 FILLER_111_1025 ();
 FILLCELL_X32 FILLER_111_1057 ();
 FILLCELL_X32 FILLER_111_1089 ();
 FILLCELL_X32 FILLER_111_1121 ();
 FILLCELL_X32 FILLER_111_1153 ();
 FILLCELL_X32 FILLER_111_1185 ();
 FILLCELL_X32 FILLER_111_1217 ();
 FILLCELL_X8 FILLER_111_1249 ();
 FILLCELL_X4 FILLER_111_1257 ();
 FILLCELL_X2 FILLER_111_1261 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X16 FILLER_111_1296 ();
 FILLCELL_X4 FILLER_111_1312 ();
 FILLCELL_X2 FILLER_111_1326 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X32 FILLER_112_952 ();
 FILLCELL_X32 FILLER_112_984 ();
 FILLCELL_X32 FILLER_112_1016 ();
 FILLCELL_X32 FILLER_112_1048 ();
 FILLCELL_X32 FILLER_112_1080 ();
 FILLCELL_X32 FILLER_112_1112 ();
 FILLCELL_X32 FILLER_112_1144 ();
 FILLCELL_X32 FILLER_112_1176 ();
 FILLCELL_X32 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_112_1240 ();
 FILLCELL_X16 FILLER_112_1272 ();
 FILLCELL_X4 FILLER_112_1288 ();
 FILLCELL_X2 FILLER_112_1292 ();
 FILLCELL_X1 FILLER_112_1294 ();
 FILLCELL_X4 FILLER_112_1298 ();
 FILLCELL_X2 FILLER_112_1302 ();
 FILLCELL_X8 FILLER_112_1308 ();
 FILLCELL_X2 FILLER_112_1321 ();
 FILLCELL_X16 FILLER_113_1 ();
 FILLCELL_X4 FILLER_113_17 ();
 FILLCELL_X2 FILLER_113_21 ();
 FILLCELL_X1 FILLER_113_23 ();
 FILLCELL_X32 FILLER_113_28 ();
 FILLCELL_X32 FILLER_113_60 ();
 FILLCELL_X32 FILLER_113_92 ();
 FILLCELL_X32 FILLER_113_124 ();
 FILLCELL_X32 FILLER_113_156 ();
 FILLCELL_X32 FILLER_113_188 ();
 FILLCELL_X32 FILLER_113_220 ();
 FILLCELL_X32 FILLER_113_252 ();
 FILLCELL_X32 FILLER_113_284 ();
 FILLCELL_X32 FILLER_113_316 ();
 FILLCELL_X32 FILLER_113_348 ();
 FILLCELL_X32 FILLER_113_380 ();
 FILLCELL_X32 FILLER_113_412 ();
 FILLCELL_X32 FILLER_113_444 ();
 FILLCELL_X32 FILLER_113_476 ();
 FILLCELL_X32 FILLER_113_508 ();
 FILLCELL_X32 FILLER_113_540 ();
 FILLCELL_X32 FILLER_113_572 ();
 FILLCELL_X32 FILLER_113_604 ();
 FILLCELL_X32 FILLER_113_636 ();
 FILLCELL_X32 FILLER_113_668 ();
 FILLCELL_X32 FILLER_113_700 ();
 FILLCELL_X32 FILLER_113_732 ();
 FILLCELL_X32 FILLER_113_764 ();
 FILLCELL_X32 FILLER_113_796 ();
 FILLCELL_X32 FILLER_113_828 ();
 FILLCELL_X32 FILLER_113_860 ();
 FILLCELL_X32 FILLER_113_892 ();
 FILLCELL_X32 FILLER_113_924 ();
 FILLCELL_X32 FILLER_113_956 ();
 FILLCELL_X32 FILLER_113_988 ();
 FILLCELL_X32 FILLER_113_1020 ();
 FILLCELL_X32 FILLER_113_1052 ();
 FILLCELL_X32 FILLER_113_1084 ();
 FILLCELL_X32 FILLER_113_1116 ();
 FILLCELL_X16 FILLER_113_1148 ();
 FILLCELL_X8 FILLER_113_1164 ();
 FILLCELL_X4 FILLER_113_1172 ();
 FILLCELL_X2 FILLER_113_1176 ();
 FILLCELL_X1 FILLER_113_1178 ();
 FILLCELL_X32 FILLER_113_1196 ();
 FILLCELL_X32 FILLER_113_1228 ();
 FILLCELL_X2 FILLER_113_1260 ();
 FILLCELL_X1 FILLER_113_1262 ();
 FILLCELL_X16 FILLER_113_1264 ();
 FILLCELL_X8 FILLER_113_1280 ();
 FILLCELL_X1 FILLER_113_1288 ();
 FILLCELL_X16 FILLER_113_1293 ();
 FILLCELL_X4 FILLER_113_1309 ();
 FILLCELL_X2 FILLER_113_1313 ();
 FILLCELL_X1 FILLER_113_1315 ();
 FILLCELL_X2 FILLER_113_1321 ();
 FILLCELL_X1 FILLER_113_1323 ();
 FILLCELL_X1 FILLER_113_1327 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X32 FILLER_114_952 ();
 FILLCELL_X32 FILLER_114_984 ();
 FILLCELL_X32 FILLER_114_1016 ();
 FILLCELL_X32 FILLER_114_1048 ();
 FILLCELL_X32 FILLER_114_1080 ();
 FILLCELL_X32 FILLER_114_1112 ();
 FILLCELL_X32 FILLER_114_1144 ();
 FILLCELL_X4 FILLER_114_1176 ();
 FILLCELL_X2 FILLER_114_1180 ();
 FILLCELL_X1 FILLER_114_1182 ();
 FILLCELL_X32 FILLER_114_1187 ();
 FILLCELL_X32 FILLER_114_1219 ();
 FILLCELL_X32 FILLER_114_1251 ();
 FILLCELL_X32 FILLER_114_1283 ();
 FILLCELL_X8 FILLER_114_1315 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X32 FILLER_115_801 ();
 FILLCELL_X32 FILLER_115_833 ();
 FILLCELL_X32 FILLER_115_865 ();
 FILLCELL_X32 FILLER_115_897 ();
 FILLCELL_X32 FILLER_115_929 ();
 FILLCELL_X32 FILLER_115_961 ();
 FILLCELL_X32 FILLER_115_993 ();
 FILLCELL_X32 FILLER_115_1025 ();
 FILLCELL_X32 FILLER_115_1057 ();
 FILLCELL_X32 FILLER_115_1089 ();
 FILLCELL_X8 FILLER_115_1121 ();
 FILLCELL_X4 FILLER_115_1129 ();
 FILLCELL_X32 FILLER_115_1150 ();
 FILLCELL_X4 FILLER_115_1182 ();
 FILLCELL_X2 FILLER_115_1186 ();
 FILLCELL_X1 FILLER_115_1188 ();
 FILLCELL_X2 FILLER_115_1193 ();
 FILLCELL_X1 FILLER_115_1195 ();
 FILLCELL_X32 FILLER_115_1213 ();
 FILLCELL_X16 FILLER_115_1245 ();
 FILLCELL_X2 FILLER_115_1261 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X16 FILLER_115_1296 ();
 FILLCELL_X1 FILLER_115_1312 ();
 FILLCELL_X2 FILLER_115_1321 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X32 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_888 ();
 FILLCELL_X32 FILLER_116_920 ();
 FILLCELL_X32 FILLER_116_952 ();
 FILLCELL_X32 FILLER_116_984 ();
 FILLCELL_X32 FILLER_116_1016 ();
 FILLCELL_X32 FILLER_116_1048 ();
 FILLCELL_X32 FILLER_116_1080 ();
 FILLCELL_X8 FILLER_116_1112 ();
 FILLCELL_X4 FILLER_116_1141 ();
 FILLCELL_X2 FILLER_116_1145 ();
 FILLCELL_X1 FILLER_116_1147 ();
 FILLCELL_X8 FILLER_116_1153 ();
 FILLCELL_X4 FILLER_116_1161 ();
 FILLCELL_X2 FILLER_116_1165 ();
 FILLCELL_X4 FILLER_116_1190 ();
 FILLCELL_X8 FILLER_116_1198 ();
 FILLCELL_X32 FILLER_116_1211 ();
 FILLCELL_X32 FILLER_116_1243 ();
 FILLCELL_X32 FILLER_116_1275 ();
 FILLCELL_X4 FILLER_116_1307 ();
 FILLCELL_X2 FILLER_116_1311 ();
 FILLCELL_X1 FILLER_116_1313 ();
 FILLCELL_X4 FILLER_116_1317 ();
 FILLCELL_X2 FILLER_116_1321 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X32 FILLER_117_801 ();
 FILLCELL_X32 FILLER_117_833 ();
 FILLCELL_X32 FILLER_117_865 ();
 FILLCELL_X32 FILLER_117_897 ();
 FILLCELL_X32 FILLER_117_929 ();
 FILLCELL_X32 FILLER_117_961 ();
 FILLCELL_X32 FILLER_117_993 ();
 FILLCELL_X32 FILLER_117_1025 ();
 FILLCELL_X32 FILLER_117_1057 ();
 FILLCELL_X32 FILLER_117_1089 ();
 FILLCELL_X8 FILLER_117_1121 ();
 FILLCELL_X4 FILLER_117_1129 ();
 FILLCELL_X1 FILLER_117_1133 ();
 FILLCELL_X1 FILLER_117_1142 ();
 FILLCELL_X16 FILLER_117_1147 ();
 FILLCELL_X4 FILLER_117_1163 ();
 FILLCELL_X2 FILLER_117_1167 ();
 FILLCELL_X1 FILLER_117_1181 ();
 FILLCELL_X2 FILLER_117_1195 ();
 FILLCELL_X1 FILLER_117_1197 ();
 FILLCELL_X32 FILLER_117_1207 ();
 FILLCELL_X8 FILLER_117_1239 ();
 FILLCELL_X1 FILLER_117_1247 ();
 FILLCELL_X4 FILLER_117_1258 ();
 FILLCELL_X1 FILLER_117_1262 ();
 FILLCELL_X8 FILLER_117_1264 ();
 FILLCELL_X4 FILLER_117_1272 ();
 FILLCELL_X2 FILLER_117_1276 ();
 FILLCELL_X1 FILLER_117_1278 ();
 FILLCELL_X16 FILLER_117_1289 ();
 FILLCELL_X8 FILLER_117_1305 ();
 FILLCELL_X2 FILLER_117_1313 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X16 FILLER_118_632 ();
 FILLCELL_X4 FILLER_118_648 ();
 FILLCELL_X2 FILLER_118_652 ();
 FILLCELL_X1 FILLER_118_654 ();
 FILLCELL_X32 FILLER_118_660 ();
 FILLCELL_X32 FILLER_118_692 ();
 FILLCELL_X32 FILLER_118_724 ();
 FILLCELL_X32 FILLER_118_756 ();
 FILLCELL_X32 FILLER_118_788 ();
 FILLCELL_X32 FILLER_118_820 ();
 FILLCELL_X32 FILLER_118_852 ();
 FILLCELL_X32 FILLER_118_884 ();
 FILLCELL_X32 FILLER_118_916 ();
 FILLCELL_X32 FILLER_118_948 ();
 FILLCELL_X32 FILLER_118_980 ();
 FILLCELL_X32 FILLER_118_1012 ();
 FILLCELL_X32 FILLER_118_1044 ();
 FILLCELL_X32 FILLER_118_1076 ();
 FILLCELL_X16 FILLER_118_1108 ();
 FILLCELL_X8 FILLER_118_1124 ();
 FILLCELL_X4 FILLER_118_1132 ();
 FILLCELL_X1 FILLER_118_1136 ();
 FILLCELL_X2 FILLER_118_1158 ();
 FILLCELL_X16 FILLER_118_1164 ();
 FILLCELL_X2 FILLER_118_1180 ();
 FILLCELL_X1 FILLER_118_1182 ();
 FILLCELL_X32 FILLER_118_1200 ();
 FILLCELL_X8 FILLER_118_1232 ();
 FILLCELL_X4 FILLER_118_1240 ();
 FILLCELL_X2 FILLER_118_1244 ();
 FILLCELL_X1 FILLER_118_1246 ();
 FILLCELL_X4 FILLER_118_1266 ();
 FILLCELL_X4 FILLER_118_1280 ();
 FILLCELL_X16 FILLER_118_1288 ();
 FILLCELL_X8 FILLER_118_1304 ();
 FILLCELL_X4 FILLER_118_1312 ();
 FILLCELL_X2 FILLER_118_1316 ();
 FILLCELL_X2 FILLER_118_1326 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X32 FILLER_119_993 ();
 FILLCELL_X32 FILLER_119_1025 ();
 FILLCELL_X32 FILLER_119_1057 ();
 FILLCELL_X16 FILLER_119_1089 ();
 FILLCELL_X4 FILLER_119_1105 ();
 FILLCELL_X2 FILLER_119_1109 ();
 FILLCELL_X1 FILLER_119_1111 ();
 FILLCELL_X8 FILLER_119_1131 ();
 FILLCELL_X1 FILLER_119_1139 ();
 FILLCELL_X1 FILLER_119_1147 ();
 FILLCELL_X16 FILLER_119_1161 ();
 FILLCELL_X1 FILLER_119_1206 ();
 FILLCELL_X2 FILLER_119_1211 ();
 FILLCELL_X1 FILLER_119_1213 ();
 FILLCELL_X16 FILLER_119_1235 ();
 FILLCELL_X8 FILLER_119_1251 ();
 FILLCELL_X4 FILLER_119_1259 ();
 FILLCELL_X1 FILLER_119_1264 ();
 FILLCELL_X2 FILLER_119_1269 ();
 FILLCELL_X1 FILLER_119_1271 ();
 FILLCELL_X8 FILLER_119_1301 ();
 FILLCELL_X4 FILLER_119_1309 ();
 FILLCELL_X2 FILLER_119_1313 ();
 FILLCELL_X1 FILLER_119_1315 ();
 FILLCELL_X2 FILLER_119_1321 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X32 FILLER_120_984 ();
 FILLCELL_X32 FILLER_120_1016 ();
 FILLCELL_X32 FILLER_120_1048 ();
 FILLCELL_X16 FILLER_120_1080 ();
 FILLCELL_X8 FILLER_120_1096 ();
 FILLCELL_X2 FILLER_120_1104 ();
 FILLCELL_X1 FILLER_120_1129 ();
 FILLCELL_X4 FILLER_120_1134 ();
 FILLCELL_X2 FILLER_120_1138 ();
 FILLCELL_X16 FILLER_120_1165 ();
 FILLCELL_X8 FILLER_120_1181 ();
 FILLCELL_X1 FILLER_120_1189 ();
 FILLCELL_X1 FILLER_120_1195 ();
 FILLCELL_X2 FILLER_120_1208 ();
 FILLCELL_X32 FILLER_120_1218 ();
 FILLCELL_X16 FILLER_120_1250 ();
 FILLCELL_X4 FILLER_120_1266 ();
 FILLCELL_X2 FILLER_120_1270 ();
 FILLCELL_X1 FILLER_120_1272 ();
 FILLCELL_X8 FILLER_120_1284 ();
 FILLCELL_X1 FILLER_120_1292 ();
 FILLCELL_X8 FILLER_120_1296 ();
 FILLCELL_X4 FILLER_120_1304 ();
 FILLCELL_X2 FILLER_120_1308 ();
 FILLCELL_X1 FILLER_120_1310 ();
 FILLCELL_X2 FILLER_120_1326 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X32 FILLER_121_993 ();
 FILLCELL_X32 FILLER_121_1025 ();
 FILLCELL_X32 FILLER_121_1057 ();
 FILLCELL_X16 FILLER_121_1089 ();
 FILLCELL_X8 FILLER_121_1105 ();
 FILLCELL_X4 FILLER_121_1113 ();
 FILLCELL_X8 FILLER_121_1124 ();
 FILLCELL_X2 FILLER_121_1139 ();
 FILLCELL_X32 FILLER_121_1151 ();
 FILLCELL_X2 FILLER_121_1183 ();
 FILLCELL_X32 FILLER_121_1208 ();
 FILLCELL_X16 FILLER_121_1240 ();
 FILLCELL_X4 FILLER_121_1256 ();
 FILLCELL_X2 FILLER_121_1260 ();
 FILLCELL_X1 FILLER_121_1262 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X16 FILLER_121_1296 ();
 FILLCELL_X4 FILLER_121_1312 ();
 FILLCELL_X2 FILLER_121_1316 ();
 FILLCELL_X1 FILLER_121_1318 ();
 FILLCELL_X1 FILLER_121_1322 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X32 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_122_1048 ();
 FILLCELL_X32 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1112 ();
 FILLCELL_X32 FILLER_122_1144 ();
 FILLCELL_X32 FILLER_122_1176 ();
 FILLCELL_X4 FILLER_122_1208 ();
 FILLCELL_X2 FILLER_122_1212 ();
 FILLCELL_X1 FILLER_122_1214 ();
 FILLCELL_X4 FILLER_122_1232 ();
 FILLCELL_X1 FILLER_122_1236 ();
 FILLCELL_X16 FILLER_122_1286 ();
 FILLCELL_X4 FILLER_122_1302 ();
 FILLCELL_X1 FILLER_122_1306 ();
 FILLCELL_X8 FILLER_122_1311 ();
 FILLCELL_X4 FILLER_122_1319 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X32 FILLER_123_993 ();
 FILLCELL_X32 FILLER_123_1025 ();
 FILLCELL_X32 FILLER_123_1057 ();
 FILLCELL_X16 FILLER_123_1089 ();
 FILLCELL_X4 FILLER_123_1105 ();
 FILLCELL_X1 FILLER_123_1109 ();
 FILLCELL_X16 FILLER_123_1133 ();
 FILLCELL_X2 FILLER_123_1149 ();
 FILLCELL_X1 FILLER_123_1151 ();
 FILLCELL_X32 FILLER_123_1185 ();
 FILLCELL_X1 FILLER_123_1221 ();
 FILLCELL_X4 FILLER_123_1225 ();
 FILLCELL_X2 FILLER_123_1229 ();
 FILLCELL_X8 FILLER_123_1234 ();
 FILLCELL_X16 FILLER_123_1288 ();
 FILLCELL_X2 FILLER_123_1304 ();
 FILLCELL_X1 FILLER_123_1306 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X4 FILLER_124_1144 ();
 FILLCELL_X1 FILLER_124_1148 ();
 FILLCELL_X4 FILLER_124_1170 ();
 FILLCELL_X2 FILLER_124_1174 ();
 FILLCELL_X1 FILLER_124_1176 ();
 FILLCELL_X16 FILLER_124_1186 ();
 FILLCELL_X1 FILLER_124_1202 ();
 FILLCELL_X2 FILLER_124_1209 ();
 FILLCELL_X8 FILLER_124_1230 ();
 FILLCELL_X4 FILLER_124_1238 ();
 FILLCELL_X1 FILLER_124_1242 ();
 FILLCELL_X8 FILLER_124_1253 ();
 FILLCELL_X4 FILLER_124_1261 ();
 FILLCELL_X1 FILLER_124_1265 ();
 FILLCELL_X2 FILLER_124_1269 ();
 FILLCELL_X1 FILLER_124_1312 ();
 FILLCELL_X1 FILLER_124_1321 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X32 FILLER_125_961 ();
 FILLCELL_X32 FILLER_125_993 ();
 FILLCELL_X32 FILLER_125_1025 ();
 FILLCELL_X32 FILLER_125_1057 ();
 FILLCELL_X16 FILLER_125_1089 ();
 FILLCELL_X8 FILLER_125_1105 ();
 FILLCELL_X4 FILLER_125_1113 ();
 FILLCELL_X2 FILLER_125_1117 ();
 FILLCELL_X4 FILLER_125_1131 ();
 FILLCELL_X16 FILLER_125_1179 ();
 FILLCELL_X4 FILLER_125_1195 ();
 FILLCELL_X1 FILLER_125_1199 ();
 FILLCELL_X4 FILLER_125_1210 ();
 FILLCELL_X2 FILLER_125_1214 ();
 FILLCELL_X1 FILLER_125_1216 ();
 FILLCELL_X2 FILLER_125_1220 ();
 FILLCELL_X32 FILLER_125_1226 ();
 FILLCELL_X4 FILLER_125_1258 ();
 FILLCELL_X1 FILLER_125_1262 ();
 FILLCELL_X8 FILLER_125_1264 ();
 FILLCELL_X4 FILLER_125_1272 ();
 FILLCELL_X2 FILLER_125_1304 ();
 FILLCELL_X1 FILLER_125_1306 ();
 FILLCELL_X4 FILLER_125_1310 ();
 FILLCELL_X2 FILLER_125_1314 ();
 FILLCELL_X1 FILLER_125_1316 ();
 FILLCELL_X8 FILLER_125_1320 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_126_1048 ();
 FILLCELL_X32 FILLER_126_1080 ();
 FILLCELL_X2 FILLER_126_1112 ();
 FILLCELL_X1 FILLER_126_1114 ();
 FILLCELL_X8 FILLER_126_1118 ();
 FILLCELL_X2 FILLER_126_1126 ();
 FILLCELL_X1 FILLER_126_1128 ();
 FILLCELL_X1 FILLER_126_1150 ();
 FILLCELL_X1 FILLER_126_1172 ();
 FILLCELL_X2 FILLER_126_1190 ();
 FILLCELL_X4 FILLER_126_1194 ();
 FILLCELL_X2 FILLER_126_1198 ();
 FILLCELL_X1 FILLER_126_1200 ();
 FILLCELL_X32 FILLER_126_1224 ();
 FILLCELL_X32 FILLER_126_1256 ();
 FILLCELL_X16 FILLER_126_1288 ();
 FILLCELL_X2 FILLER_126_1314 ();
 FILLCELL_X1 FILLER_126_1316 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X4 FILLER_127_1089 ();
 FILLCELL_X1 FILLER_127_1093 ();
 FILLCELL_X8 FILLER_127_1099 ();
 FILLCELL_X4 FILLER_127_1107 ();
 FILLCELL_X1 FILLER_127_1111 ();
 FILLCELL_X16 FILLER_127_1129 ();
 FILLCELL_X4 FILLER_127_1145 ();
 FILLCELL_X1 FILLER_127_1149 ();
 FILLCELL_X8 FILLER_127_1155 ();
 FILLCELL_X4 FILLER_127_1163 ();
 FILLCELL_X1 FILLER_127_1167 ();
 FILLCELL_X32 FILLER_127_1173 ();
 FILLCELL_X8 FILLER_127_1205 ();
 FILLCELL_X2 FILLER_127_1213 ();
 FILLCELL_X4 FILLER_127_1228 ();
 FILLCELL_X2 FILLER_127_1232 ();
 FILLCELL_X1 FILLER_127_1234 ();
 FILLCELL_X1 FILLER_127_1239 ();
 FILLCELL_X4 FILLER_127_1245 ();
 FILLCELL_X2 FILLER_127_1249 ();
 FILLCELL_X1 FILLER_127_1251 ();
 FILLCELL_X4 FILLER_127_1258 ();
 FILLCELL_X1 FILLER_127_1262 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X4 FILLER_127_1296 ();
 FILLCELL_X1 FILLER_127_1300 ();
 FILLCELL_X8 FILLER_127_1304 ();
 FILLCELL_X1 FILLER_127_1312 ();
 FILLCELL_X4 FILLER_127_1316 ();
 FILLCELL_X2 FILLER_127_1320 ();
 FILLCELL_X1 FILLER_127_1322 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X32 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_128_1048 ();
 FILLCELL_X32 FILLER_128_1080 ();
 FILLCELL_X16 FILLER_128_1112 ();
 FILLCELL_X4 FILLER_128_1128 ();
 FILLCELL_X2 FILLER_128_1132 ();
 FILLCELL_X1 FILLER_128_1134 ();
 FILLCELL_X32 FILLER_128_1151 ();
 FILLCELL_X16 FILLER_128_1183 ();
 FILLCELL_X4 FILLER_128_1199 ();
 FILLCELL_X8 FILLER_128_1208 ();
 FILLCELL_X4 FILLER_128_1216 ();
 FILLCELL_X2 FILLER_128_1220 ();
 FILLCELL_X1 FILLER_128_1222 ();
 FILLCELL_X1 FILLER_128_1232 ();
 FILLCELL_X4 FILLER_128_1237 ();
 FILLCELL_X1 FILLER_128_1244 ();
 FILLCELL_X16 FILLER_128_1262 ();
 FILLCELL_X4 FILLER_128_1278 ();
 FILLCELL_X2 FILLER_128_1282 ();
 FILLCELL_X1 FILLER_128_1284 ();
 FILLCELL_X1 FILLER_128_1297 ();
 FILLCELL_X16 FILLER_128_1300 ();
 FILLCELL_X4 FILLER_128_1316 ();
 FILLCELL_X2 FILLER_128_1320 ();
 FILLCELL_X1 FILLER_128_1322 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_993 ();
 FILLCELL_X32 FILLER_129_1025 ();
 FILLCELL_X32 FILLER_129_1057 ();
 FILLCELL_X16 FILLER_129_1089 ();
 FILLCELL_X16 FILLER_129_1136 ();
 FILLCELL_X4 FILLER_129_1157 ();
 FILLCELL_X2 FILLER_129_1161 ();
 FILLCELL_X1 FILLER_129_1163 ();
 FILLCELL_X16 FILLER_129_1171 ();
 FILLCELL_X4 FILLER_129_1187 ();
 FILLCELL_X2 FILLER_129_1191 ();
 FILLCELL_X1 FILLER_129_1193 ();
 FILLCELL_X4 FILLER_129_1215 ();
 FILLCELL_X1 FILLER_129_1219 ();
 FILLCELL_X16 FILLER_129_1234 ();
 FILLCELL_X8 FILLER_129_1250 ();
 FILLCELL_X4 FILLER_129_1258 ();
 FILLCELL_X1 FILLER_129_1262 ();
 FILLCELL_X16 FILLER_129_1264 ();
 FILLCELL_X2 FILLER_129_1280 ();
 FILLCELL_X1 FILLER_129_1282 ();
 FILLCELL_X2 FILLER_129_1299 ();
 FILLCELL_X1 FILLER_129_1301 ();
 FILLCELL_X8 FILLER_129_1305 ();
 FILLCELL_X4 FILLER_129_1313 ();
 FILLCELL_X1 FILLER_129_1317 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X32 FILLER_130_1016 ();
 FILLCELL_X32 FILLER_130_1048 ();
 FILLCELL_X4 FILLER_130_1080 ();
 FILLCELL_X2 FILLER_130_1084 ();
 FILLCELL_X32 FILLER_130_1095 ();
 FILLCELL_X4 FILLER_130_1127 ();
 FILLCELL_X1 FILLER_130_1131 ();
 FILLCELL_X16 FILLER_130_1137 ();
 FILLCELL_X4 FILLER_130_1153 ();
 FILLCELL_X4 FILLER_130_1161 ();
 FILLCELL_X2 FILLER_130_1165 ();
 FILLCELL_X32 FILLER_130_1172 ();
 FILLCELL_X4 FILLER_130_1204 ();
 FILLCELL_X2 FILLER_130_1224 ();
 FILLCELL_X32 FILLER_130_1232 ();
 FILLCELL_X16 FILLER_130_1264 ();
 FILLCELL_X2 FILLER_130_1280 ();
 FILLCELL_X8 FILLER_130_1286 ();
 FILLCELL_X8 FILLER_130_1297 ();
 FILLCELL_X2 FILLER_130_1308 ();
 FILLCELL_X2 FILLER_130_1313 ();
 FILLCELL_X1 FILLER_130_1315 ();
 FILLCELL_X2 FILLER_130_1321 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_584 ();
 FILLCELL_X32 FILLER_131_616 ();
 FILLCELL_X32 FILLER_131_648 ();
 FILLCELL_X32 FILLER_131_680 ();
 FILLCELL_X32 FILLER_131_712 ();
 FILLCELL_X32 FILLER_131_744 ();
 FILLCELL_X32 FILLER_131_776 ();
 FILLCELL_X32 FILLER_131_808 ();
 FILLCELL_X32 FILLER_131_840 ();
 FILLCELL_X32 FILLER_131_872 ();
 FILLCELL_X32 FILLER_131_904 ();
 FILLCELL_X32 FILLER_131_936 ();
 FILLCELL_X32 FILLER_131_968 ();
 FILLCELL_X32 FILLER_131_1000 ();
 FILLCELL_X32 FILLER_131_1032 ();
 FILLCELL_X32 FILLER_131_1064 ();
 FILLCELL_X32 FILLER_131_1096 ();
 FILLCELL_X16 FILLER_131_1133 ();
 FILLCELL_X4 FILLER_131_1149 ();
 FILLCELL_X32 FILLER_131_1175 ();
 FILLCELL_X32 FILLER_131_1207 ();
 FILLCELL_X2 FILLER_131_1239 ();
 FILLCELL_X4 FILLER_131_1248 ();
 FILLCELL_X2 FILLER_131_1252 ();
 FILLCELL_X1 FILLER_131_1254 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X4 FILLER_131_1264 ();
 FILLCELL_X2 FILLER_131_1268 ();
 FILLCELL_X16 FILLER_131_1298 ();
 FILLCELL_X4 FILLER_131_1314 ();
 FILLCELL_X1 FILLER_131_1318 ();
 FILLCELL_X1 FILLER_131_1322 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X4 FILLER_132_577 ();
 FILLCELL_X2 FILLER_132_581 ();
 FILLCELL_X32 FILLER_132_590 ();
 FILLCELL_X8 FILLER_132_622 ();
 FILLCELL_X1 FILLER_132_630 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X32 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_132_1048 ();
 FILLCELL_X16 FILLER_132_1080 ();
 FILLCELL_X8 FILLER_132_1096 ();
 FILLCELL_X2 FILLER_132_1104 ();
 FILLCELL_X1 FILLER_132_1106 ();
 FILLCELL_X32 FILLER_132_1112 ();
 FILLCELL_X4 FILLER_132_1144 ();
 FILLCELL_X2 FILLER_132_1148 ();
 FILLCELL_X1 FILLER_132_1150 ();
 FILLCELL_X1 FILLER_132_1158 ();
 FILLCELL_X4 FILLER_132_1162 ();
 FILLCELL_X2 FILLER_132_1166 ();
 FILLCELL_X1 FILLER_132_1168 ();
 FILLCELL_X8 FILLER_132_1174 ();
 FILLCELL_X1 FILLER_132_1182 ();
 FILLCELL_X16 FILLER_132_1187 ();
 FILLCELL_X2 FILLER_132_1203 ();
 FILLCELL_X1 FILLER_132_1205 ();
 FILLCELL_X4 FILLER_132_1217 ();
 FILLCELL_X1 FILLER_132_1221 ();
 FILLCELL_X4 FILLER_132_1231 ();
 FILLCELL_X1 FILLER_132_1235 ();
 FILLCELL_X8 FILLER_132_1263 ();
 FILLCELL_X4 FILLER_132_1271 ();
 FILLCELL_X2 FILLER_132_1275 ();
 FILLCELL_X16 FILLER_132_1297 ();
 FILLCELL_X1 FILLER_132_1313 ();
 FILLCELL_X1 FILLER_132_1327 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X32 FILLER_133_993 ();
 FILLCELL_X32 FILLER_133_1025 ();
 FILLCELL_X32 FILLER_133_1057 ();
 FILLCELL_X32 FILLER_133_1089 ();
 FILLCELL_X4 FILLER_133_1121 ();
 FILLCELL_X1 FILLER_133_1125 ();
 FILLCELL_X32 FILLER_133_1128 ();
 FILLCELL_X16 FILLER_133_1160 ();
 FILLCELL_X8 FILLER_133_1176 ();
 FILLCELL_X4 FILLER_133_1208 ();
 FILLCELL_X2 FILLER_133_1212 ();
 FILLCELL_X32 FILLER_133_1228 ();
 FILLCELL_X2 FILLER_133_1260 ();
 FILLCELL_X1 FILLER_133_1262 ();
 FILLCELL_X8 FILLER_133_1264 ();
 FILLCELL_X4 FILLER_133_1272 ();
 FILLCELL_X2 FILLER_133_1276 ();
 FILLCELL_X2 FILLER_133_1289 ();
 FILLCELL_X1 FILLER_133_1291 ();
 FILLCELL_X16 FILLER_133_1296 ();
 FILLCELL_X2 FILLER_133_1312 ();
 FILLCELL_X1 FILLER_133_1314 ();
 FILLCELL_X1 FILLER_133_1325 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X16 FILLER_134_696 ();
 FILLCELL_X2 FILLER_134_712 ();
 FILLCELL_X1 FILLER_134_714 ();
 FILLCELL_X32 FILLER_134_722 ();
 FILLCELL_X32 FILLER_134_754 ();
 FILLCELL_X32 FILLER_134_786 ();
 FILLCELL_X32 FILLER_134_818 ();
 FILLCELL_X32 FILLER_134_850 ();
 FILLCELL_X32 FILLER_134_882 ();
 FILLCELL_X32 FILLER_134_914 ();
 FILLCELL_X32 FILLER_134_946 ();
 FILLCELL_X32 FILLER_134_978 ();
 FILLCELL_X32 FILLER_134_1010 ();
 FILLCELL_X32 FILLER_134_1042 ();
 FILLCELL_X8 FILLER_134_1074 ();
 FILLCELL_X1 FILLER_134_1082 ();
 FILLCELL_X2 FILLER_134_1092 ();
 FILLCELL_X2 FILLER_134_1098 ();
 FILLCELL_X1 FILLER_134_1120 ();
 FILLCELL_X32 FILLER_134_1150 ();
 FILLCELL_X4 FILLER_134_1182 ();
 FILLCELL_X2 FILLER_134_1186 ();
 FILLCELL_X16 FILLER_134_1192 ();
 FILLCELL_X2 FILLER_134_1208 ();
 FILLCELL_X1 FILLER_134_1210 ();
 FILLCELL_X1 FILLER_134_1221 ();
 FILLCELL_X4 FILLER_134_1225 ();
 FILLCELL_X1 FILLER_134_1229 ();
 FILLCELL_X32 FILLER_134_1236 ();
 FILLCELL_X8 FILLER_134_1268 ();
 FILLCELL_X4 FILLER_134_1276 ();
 FILLCELL_X16 FILLER_134_1293 ();
 FILLCELL_X8 FILLER_134_1315 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X16 FILLER_135_641 ();
 FILLCELL_X8 FILLER_135_657 ();
 FILLCELL_X4 FILLER_135_665 ();
 FILLCELL_X1 FILLER_135_669 ();
 FILLCELL_X16 FILLER_135_687 ();
 FILLCELL_X1 FILLER_135_703 ();
 FILLCELL_X1 FILLER_135_730 ();
 FILLCELL_X32 FILLER_135_736 ();
 FILLCELL_X32 FILLER_135_768 ();
 FILLCELL_X32 FILLER_135_800 ();
 FILLCELL_X32 FILLER_135_832 ();
 FILLCELL_X32 FILLER_135_864 ();
 FILLCELL_X32 FILLER_135_896 ();
 FILLCELL_X32 FILLER_135_928 ();
 FILLCELL_X32 FILLER_135_960 ();
 FILLCELL_X32 FILLER_135_992 ();
 FILLCELL_X32 FILLER_135_1024 ();
 FILLCELL_X4 FILLER_135_1056 ();
 FILLCELL_X8 FILLER_135_1079 ();
 FILLCELL_X4 FILLER_135_1087 ();
 FILLCELL_X2 FILLER_135_1091 ();
 FILLCELL_X16 FILLER_135_1108 ();
 FILLCELL_X8 FILLER_135_1124 ();
 FILLCELL_X4 FILLER_135_1132 ();
 FILLCELL_X2 FILLER_135_1136 ();
 FILLCELL_X32 FILLER_135_1151 ();
 FILLCELL_X16 FILLER_135_1183 ();
 FILLCELL_X4 FILLER_135_1199 ();
 FILLCELL_X2 FILLER_135_1203 ();
 FILLCELL_X1 FILLER_135_1205 ();
 FILLCELL_X16 FILLER_135_1223 ();
 FILLCELL_X8 FILLER_135_1239 ();
 FILLCELL_X2 FILLER_135_1247 ();
 FILLCELL_X1 FILLER_135_1249 ();
 FILLCELL_X2 FILLER_135_1260 ();
 FILLCELL_X1 FILLER_135_1262 ();
 FILLCELL_X2 FILLER_135_1264 ();
 FILLCELL_X1 FILLER_135_1266 ();
 FILLCELL_X32 FILLER_135_1285 ();
 FILLCELL_X1 FILLER_135_1327 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X16 FILLER_136_545 ();
 FILLCELL_X2 FILLER_136_561 ();
 FILLCELL_X1 FILLER_136_563 ();
 FILLCELL_X32 FILLER_136_571 ();
 FILLCELL_X16 FILLER_136_603 ();
 FILLCELL_X8 FILLER_136_619 ();
 FILLCELL_X4 FILLER_136_627 ();
 FILLCELL_X16 FILLER_136_632 ();
 FILLCELL_X8 FILLER_136_648 ();
 FILLCELL_X2 FILLER_136_656 ();
 FILLCELL_X4 FILLER_136_662 ();
 FILLCELL_X2 FILLER_136_666 ();
 FILLCELL_X8 FILLER_136_675 ();
 FILLCELL_X1 FILLER_136_683 ();
 FILLCELL_X4 FILLER_136_689 ();
 FILLCELL_X1 FILLER_136_693 ();
 FILLCELL_X4 FILLER_136_707 ();
 FILLCELL_X2 FILLER_136_711 ();
 FILLCELL_X8 FILLER_136_718 ();
 FILLCELL_X4 FILLER_136_726 ();
 FILLCELL_X1 FILLER_136_730 ();
 FILLCELL_X32 FILLER_136_755 ();
 FILLCELL_X32 FILLER_136_787 ();
 FILLCELL_X32 FILLER_136_819 ();
 FILLCELL_X32 FILLER_136_851 ();
 FILLCELL_X32 FILLER_136_883 ();
 FILLCELL_X32 FILLER_136_915 ();
 FILLCELL_X32 FILLER_136_947 ();
 FILLCELL_X32 FILLER_136_979 ();
 FILLCELL_X32 FILLER_136_1011 ();
 FILLCELL_X32 FILLER_136_1043 ();
 FILLCELL_X1 FILLER_136_1075 ();
 FILLCELL_X32 FILLER_136_1104 ();
 FILLCELL_X8 FILLER_136_1136 ();
 FILLCELL_X8 FILLER_136_1162 ();
 FILLCELL_X32 FILLER_136_1175 ();
 FILLCELL_X32 FILLER_136_1207 ();
 FILLCELL_X16 FILLER_136_1239 ();
 FILLCELL_X1 FILLER_136_1255 ();
 FILLCELL_X16 FILLER_136_1283 ();
 FILLCELL_X8 FILLER_136_1299 ();
 FILLCELL_X4 FILLER_136_1307 ();
 FILLCELL_X1 FILLER_136_1316 ();
 FILLCELL_X2 FILLER_136_1322 ();
 FILLCELL_X1 FILLER_136_1327 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X16 FILLER_137_641 ();
 FILLCELL_X8 FILLER_137_673 ();
 FILLCELL_X4 FILLER_137_681 ();
 FILLCELL_X1 FILLER_137_685 ();
 FILLCELL_X4 FILLER_137_692 ();
 FILLCELL_X1 FILLER_137_696 ();
 FILLCELL_X1 FILLER_137_712 ();
 FILLCELL_X1 FILLER_137_717 ();
 FILLCELL_X32 FILLER_137_723 ();
 FILLCELL_X32 FILLER_137_755 ();
 FILLCELL_X32 FILLER_137_787 ();
 FILLCELL_X32 FILLER_137_819 ();
 FILLCELL_X32 FILLER_137_851 ();
 FILLCELL_X32 FILLER_137_883 ();
 FILLCELL_X32 FILLER_137_915 ();
 FILLCELL_X32 FILLER_137_947 ();
 FILLCELL_X32 FILLER_137_979 ();
 FILLCELL_X32 FILLER_137_1011 ();
 FILLCELL_X8 FILLER_137_1043 ();
 FILLCELL_X4 FILLER_137_1051 ();
 FILLCELL_X16 FILLER_137_1069 ();
 FILLCELL_X2 FILLER_137_1085 ();
 FILLCELL_X1 FILLER_137_1087 ();
 FILLCELL_X32 FILLER_137_1102 ();
 FILLCELL_X16 FILLER_137_1134 ();
 FILLCELL_X2 FILLER_137_1150 ();
 FILLCELL_X1 FILLER_137_1152 ();
 FILLCELL_X4 FILLER_137_1157 ();
 FILLCELL_X2 FILLER_137_1161 ();
 FILLCELL_X1 FILLER_137_1163 ();
 FILLCELL_X2 FILLER_137_1186 ();
 FILLCELL_X1 FILLER_137_1192 ();
 FILLCELL_X32 FILLER_137_1196 ();
 FILLCELL_X16 FILLER_137_1237 ();
 FILLCELL_X8 FILLER_137_1253 ();
 FILLCELL_X2 FILLER_137_1261 ();
 FILLCELL_X2 FILLER_137_1268 ();
 FILLCELL_X16 FILLER_137_1284 ();
 FILLCELL_X8 FILLER_137_1300 ();
 FILLCELL_X2 FILLER_137_1308 ();
 FILLCELL_X1 FILLER_137_1310 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X8 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_617 ();
 FILLCELL_X2 FILLER_138_628 ();
 FILLCELL_X1 FILLER_138_630 ();
 FILLCELL_X4 FILLER_138_636 ();
 FILLCELL_X4 FILLER_138_662 ();
 FILLCELL_X1 FILLER_138_666 ();
 FILLCELL_X16 FILLER_138_670 ();
 FILLCELL_X4 FILLER_138_686 ();
 FILLCELL_X2 FILLER_138_690 ();
 FILLCELL_X4 FILLER_138_697 ();
 FILLCELL_X1 FILLER_138_701 ();
 FILLCELL_X32 FILLER_138_710 ();
 FILLCELL_X32 FILLER_138_742 ();
 FILLCELL_X32 FILLER_138_774 ();
 FILLCELL_X32 FILLER_138_806 ();
 FILLCELL_X32 FILLER_138_838 ();
 FILLCELL_X32 FILLER_138_870 ();
 FILLCELL_X32 FILLER_138_902 ();
 FILLCELL_X32 FILLER_138_934 ();
 FILLCELL_X32 FILLER_138_966 ();
 FILLCELL_X32 FILLER_138_998 ();
 FILLCELL_X32 FILLER_138_1030 ();
 FILLCELL_X32 FILLER_138_1062 ();
 FILLCELL_X32 FILLER_138_1094 ();
 FILLCELL_X4 FILLER_138_1126 ();
 FILLCELL_X2 FILLER_138_1130 ();
 FILLCELL_X1 FILLER_138_1132 ();
 FILLCELL_X1 FILLER_138_1145 ();
 FILLCELL_X8 FILLER_138_1159 ();
 FILLCELL_X4 FILLER_138_1167 ();
 FILLCELL_X2 FILLER_138_1171 ();
 FILLCELL_X2 FILLER_138_1177 ();
 FILLCELL_X1 FILLER_138_1179 ();
 FILLCELL_X2 FILLER_138_1191 ();
 FILLCELL_X1 FILLER_138_1193 ();
 FILLCELL_X8 FILLER_138_1200 ();
 FILLCELL_X4 FILLER_138_1208 ();
 FILLCELL_X2 FILLER_138_1212 ();
 FILLCELL_X1 FILLER_138_1214 ();
 FILLCELL_X4 FILLER_138_1227 ();
 FILLCELL_X2 FILLER_138_1234 ();
 FILLCELL_X1 FILLER_138_1236 ();
 FILLCELL_X16 FILLER_138_1247 ();
 FILLCELL_X2 FILLER_138_1284 ();
 FILLCELL_X2 FILLER_138_1296 ();
 FILLCELL_X1 FILLER_138_1298 ();
 FILLCELL_X4 FILLER_138_1302 ();
 FILLCELL_X1 FILLER_138_1306 ();
 FILLCELL_X4 FILLER_138_1309 ();
 FILLCELL_X1 FILLER_138_1313 ();
 FILLCELL_X2 FILLER_138_1317 ();
 FILLCELL_X4 FILLER_138_1324 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X16 FILLER_139_577 ();
 FILLCELL_X4 FILLER_139_593 ();
 FILLCELL_X2 FILLER_139_597 ();
 FILLCELL_X1 FILLER_139_599 ();
 FILLCELL_X8 FILLER_139_642 ();
 FILLCELL_X32 FILLER_139_669 ();
 FILLCELL_X4 FILLER_139_701 ();
 FILLCELL_X8 FILLER_139_707 ();
 FILLCELL_X4 FILLER_139_715 ();
 FILLCELL_X2 FILLER_139_719 ();
 FILLCELL_X1 FILLER_139_721 ();
 FILLCELL_X32 FILLER_139_727 ();
 FILLCELL_X32 FILLER_139_759 ();
 FILLCELL_X32 FILLER_139_791 ();
 FILLCELL_X32 FILLER_139_823 ();
 FILLCELL_X32 FILLER_139_855 ();
 FILLCELL_X32 FILLER_139_887 ();
 FILLCELL_X32 FILLER_139_919 ();
 FILLCELL_X32 FILLER_139_951 ();
 FILLCELL_X32 FILLER_139_983 ();
 FILLCELL_X32 FILLER_139_1015 ();
 FILLCELL_X32 FILLER_139_1047 ();
 FILLCELL_X32 FILLER_139_1079 ();
 FILLCELL_X8 FILLER_139_1111 ();
 FILLCELL_X2 FILLER_139_1119 ();
 FILLCELL_X2 FILLER_139_1138 ();
 FILLCELL_X2 FILLER_139_1146 ();
 FILLCELL_X1 FILLER_139_1148 ();
 FILLCELL_X16 FILLER_139_1163 ();
 FILLCELL_X1 FILLER_139_1179 ();
 FILLCELL_X16 FILLER_139_1201 ();
 FILLCELL_X4 FILLER_139_1217 ();
 FILLCELL_X16 FILLER_139_1240 ();
 FILLCELL_X4 FILLER_139_1256 ();
 FILLCELL_X2 FILLER_139_1260 ();
 FILLCELL_X1 FILLER_139_1262 ();
 FILLCELL_X2 FILLER_139_1268 ();
 FILLCELL_X1 FILLER_139_1270 ();
 FILLCELL_X8 FILLER_139_1282 ();
 FILLCELL_X4 FILLER_139_1290 ();
 FILLCELL_X16 FILLER_139_1296 ();
 FILLCELL_X8 FILLER_139_1312 ();
 FILLCELL_X2 FILLER_139_1320 ();
 FILLCELL_X1 FILLER_139_1322 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X16 FILLER_140_632 ();
 FILLCELL_X4 FILLER_140_648 ();
 FILLCELL_X2 FILLER_140_652 ();
 FILLCELL_X1 FILLER_140_654 ();
 FILLCELL_X4 FILLER_140_660 ();
 FILLCELL_X1 FILLER_140_664 ();
 FILLCELL_X8 FILLER_140_670 ();
 FILLCELL_X8 FILLER_140_695 ();
 FILLCELL_X4 FILLER_140_703 ();
 FILLCELL_X32 FILLER_140_724 ();
 FILLCELL_X32 FILLER_140_756 ();
 FILLCELL_X32 FILLER_140_788 ();
 FILLCELL_X32 FILLER_140_820 ();
 FILLCELL_X32 FILLER_140_852 ();
 FILLCELL_X32 FILLER_140_884 ();
 FILLCELL_X32 FILLER_140_916 ();
 FILLCELL_X32 FILLER_140_948 ();
 FILLCELL_X32 FILLER_140_980 ();
 FILLCELL_X32 FILLER_140_1012 ();
 FILLCELL_X32 FILLER_140_1044 ();
 FILLCELL_X32 FILLER_140_1076 ();
 FILLCELL_X32 FILLER_140_1108 ();
 FILLCELL_X8 FILLER_140_1140 ();
 FILLCELL_X1 FILLER_140_1148 ();
 FILLCELL_X32 FILLER_140_1159 ();
 FILLCELL_X16 FILLER_140_1191 ();
 FILLCELL_X8 FILLER_140_1207 ();
 FILLCELL_X4 FILLER_140_1215 ();
 FILLCELL_X8 FILLER_140_1222 ();
 FILLCELL_X4 FILLER_140_1230 ();
 FILLCELL_X16 FILLER_140_1243 ();
 FILLCELL_X2 FILLER_140_1259 ();
 FILLCELL_X16 FILLER_140_1296 ();
 FILLCELL_X4 FILLER_140_1312 ();
 FILLCELL_X1 FILLER_140_1316 ();
 FILLCELL_X1 FILLER_140_1327 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X32 FILLER_141_993 ();
 FILLCELL_X32 FILLER_141_1025 ();
 FILLCELL_X32 FILLER_141_1057 ();
 FILLCELL_X32 FILLER_141_1089 ();
 FILLCELL_X16 FILLER_141_1121 ();
 FILLCELL_X2 FILLER_141_1137 ();
 FILLCELL_X1 FILLER_141_1139 ();
 FILLCELL_X1 FILLER_141_1144 ();
 FILLCELL_X1 FILLER_141_1160 ();
 FILLCELL_X32 FILLER_141_1167 ();
 FILLCELL_X32 FILLER_141_1199 ();
 FILLCELL_X2 FILLER_141_1231 ();
 FILLCELL_X1 FILLER_141_1233 ();
 FILLCELL_X16 FILLER_141_1237 ();
 FILLCELL_X8 FILLER_141_1253 ();
 FILLCELL_X2 FILLER_141_1261 ();
 FILLCELL_X8 FILLER_141_1264 ();
 FILLCELL_X4 FILLER_141_1272 ();
 FILLCELL_X2 FILLER_141_1276 ();
 FILLCELL_X1 FILLER_141_1278 ();
 FILLCELL_X16 FILLER_141_1293 ();
 FILLCELL_X2 FILLER_141_1309 ();
 FILLCELL_X2 FILLER_141_1316 ();
 FILLCELL_X1 FILLER_141_1318 ();
 FILLCELL_X1 FILLER_141_1321 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X2 FILLER_142_1132 ();
 FILLCELL_X1 FILLER_142_1141 ();
 FILLCELL_X16 FILLER_142_1170 ();
 FILLCELL_X8 FILLER_142_1186 ();
 FILLCELL_X1 FILLER_142_1194 ();
 FILLCELL_X16 FILLER_142_1204 ();
 FILLCELL_X2 FILLER_142_1220 ();
 FILLCELL_X4 FILLER_142_1229 ();
 FILLCELL_X1 FILLER_142_1233 ();
 FILLCELL_X8 FILLER_142_1244 ();
 FILLCELL_X4 FILLER_142_1252 ();
 FILLCELL_X16 FILLER_142_1262 ();
 FILLCELL_X4 FILLER_142_1278 ();
 FILLCELL_X2 FILLER_142_1282 ();
 FILLCELL_X1 FILLER_142_1284 ();
 FILLCELL_X8 FILLER_142_1295 ();
 FILLCELL_X4 FILLER_142_1303 ();
 FILLCELL_X2 FILLER_142_1307 ();
 FILLCELL_X2 FILLER_142_1315 ();
 FILLCELL_X1 FILLER_142_1317 ();
 FILLCELL_X2 FILLER_142_1323 ();
 FILLCELL_X1 FILLER_142_1325 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X8 FILLER_143_641 ();
 FILLCELL_X2 FILLER_143_649 ();
 FILLCELL_X1 FILLER_143_651 ();
 FILLCELL_X32 FILLER_143_669 ();
 FILLCELL_X32 FILLER_143_701 ();
 FILLCELL_X32 FILLER_143_733 ();
 FILLCELL_X32 FILLER_143_765 ();
 FILLCELL_X32 FILLER_143_797 ();
 FILLCELL_X32 FILLER_143_829 ();
 FILLCELL_X32 FILLER_143_861 ();
 FILLCELL_X32 FILLER_143_893 ();
 FILLCELL_X32 FILLER_143_925 ();
 FILLCELL_X32 FILLER_143_957 ();
 FILLCELL_X32 FILLER_143_989 ();
 FILLCELL_X32 FILLER_143_1021 ();
 FILLCELL_X32 FILLER_143_1053 ();
 FILLCELL_X32 FILLER_143_1085 ();
 FILLCELL_X32 FILLER_143_1117 ();
 FILLCELL_X4 FILLER_143_1149 ();
 FILLCELL_X2 FILLER_143_1153 ();
 FILLCELL_X1 FILLER_143_1155 ();
 FILLCELL_X32 FILLER_143_1163 ();
 FILLCELL_X4 FILLER_143_1195 ();
 FILLCELL_X2 FILLER_143_1199 ();
 FILLCELL_X1 FILLER_143_1201 ();
 FILLCELL_X8 FILLER_143_1215 ();
 FILLCELL_X2 FILLER_143_1223 ();
 FILLCELL_X8 FILLER_143_1227 ();
 FILLCELL_X4 FILLER_143_1235 ();
 FILLCELL_X1 FILLER_143_1239 ();
 FILLCELL_X16 FILLER_143_1244 ();
 FILLCELL_X2 FILLER_143_1260 ();
 FILLCELL_X1 FILLER_143_1262 ();
 FILLCELL_X32 FILLER_143_1274 ();
 FILLCELL_X8 FILLER_143_1306 ();
 FILLCELL_X2 FILLER_143_1314 ();
 FILLCELL_X1 FILLER_143_1316 ();
 FILLCELL_X1 FILLER_143_1324 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X8 FILLER_144_1144 ();
 FILLCELL_X2 FILLER_144_1152 ();
 FILLCELL_X1 FILLER_144_1154 ();
 FILLCELL_X8 FILLER_144_1162 ();
 FILLCELL_X4 FILLER_144_1170 ();
 FILLCELL_X1 FILLER_144_1174 ();
 FILLCELL_X4 FILLER_144_1177 ();
 FILLCELL_X1 FILLER_144_1191 ();
 FILLCELL_X1 FILLER_144_1201 ();
 FILLCELL_X2 FILLER_144_1213 ();
 FILLCELL_X2 FILLER_144_1223 ();
 FILLCELL_X1 FILLER_144_1225 ();
 FILLCELL_X4 FILLER_144_1238 ();
 FILLCELL_X2 FILLER_144_1242 ();
 FILLCELL_X1 FILLER_144_1244 ();
 FILLCELL_X32 FILLER_144_1266 ();
 FILLCELL_X16 FILLER_144_1298 ();
 FILLCELL_X2 FILLER_144_1316 ();
 FILLCELL_X2 FILLER_144_1321 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X16 FILLER_145_1121 ();
 FILLCELL_X1 FILLER_145_1137 ();
 FILLCELL_X8 FILLER_145_1159 ();
 FILLCELL_X4 FILLER_145_1167 ();
 FILLCELL_X2 FILLER_145_1171 ();
 FILLCELL_X8 FILLER_145_1186 ();
 FILLCELL_X4 FILLER_145_1194 ();
 FILLCELL_X4 FILLER_145_1211 ();
 FILLCELL_X2 FILLER_145_1215 ();
 FILLCELL_X1 FILLER_145_1217 ();
 FILLCELL_X1 FILLER_145_1234 ();
 FILLCELL_X8 FILLER_145_1238 ();
 FILLCELL_X8 FILLER_145_1255 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X8 FILLER_145_1296 ();
 FILLCELL_X4 FILLER_145_1304 ();
 FILLCELL_X2 FILLER_145_1308 ();
 FILLCELL_X1 FILLER_145_1310 ();
 FILLCELL_X2 FILLER_145_1321 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X8 FILLER_146_1144 ();
 FILLCELL_X2 FILLER_146_1152 ();
 FILLCELL_X1 FILLER_146_1154 ();
 FILLCELL_X8 FILLER_146_1176 ();
 FILLCELL_X4 FILLER_146_1184 ();
 FILLCELL_X2 FILLER_146_1188 ();
 FILLCELL_X8 FILLER_146_1209 ();
 FILLCELL_X4 FILLER_146_1221 ();
 FILLCELL_X2 FILLER_146_1225 ();
 FILLCELL_X32 FILLER_146_1235 ();
 FILLCELL_X32 FILLER_146_1267 ();
 FILLCELL_X16 FILLER_146_1299 ();
 FILLCELL_X2 FILLER_146_1315 ();
 FILLCELL_X1 FILLER_146_1317 ();
 FILLCELL_X1 FILLER_146_1321 ();
 FILLCELL_X1 FILLER_146_1327 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X16 FILLER_147_1185 ();
 FILLCELL_X8 FILLER_147_1201 ();
 FILLCELL_X2 FILLER_147_1209 ();
 FILLCELL_X1 FILLER_147_1211 ();
 FILLCELL_X8 FILLER_147_1248 ();
 FILLCELL_X4 FILLER_147_1256 ();
 FILLCELL_X2 FILLER_147_1260 ();
 FILLCELL_X1 FILLER_147_1262 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X8 FILLER_147_1296 ();
 FILLCELL_X4 FILLER_147_1304 ();
 FILLCELL_X2 FILLER_147_1308 ();
 FILLCELL_X1 FILLER_147_1310 ();
 FILLCELL_X1 FILLER_147_1316 ();
 FILLCELL_X1 FILLER_147_1324 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X4 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_238 ();
 FILLCELL_X32 FILLER_148_270 ();
 FILLCELL_X32 FILLER_148_302 ();
 FILLCELL_X32 FILLER_148_334 ();
 FILLCELL_X32 FILLER_148_366 ();
 FILLCELL_X32 FILLER_148_398 ();
 FILLCELL_X32 FILLER_148_430 ();
 FILLCELL_X32 FILLER_148_462 ();
 FILLCELL_X32 FILLER_148_494 ();
 FILLCELL_X32 FILLER_148_526 ();
 FILLCELL_X32 FILLER_148_558 ();
 FILLCELL_X32 FILLER_148_590 ();
 FILLCELL_X8 FILLER_148_622 ();
 FILLCELL_X1 FILLER_148_630 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X16 FILLER_148_1208 ();
 FILLCELL_X2 FILLER_148_1224 ();
 FILLCELL_X32 FILLER_148_1230 ();
 FILLCELL_X32 FILLER_148_1262 ();
 FILLCELL_X16 FILLER_148_1294 ();
 FILLCELL_X2 FILLER_148_1310 ();
 FILLCELL_X1 FILLER_148_1324 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X16 FILLER_149_1296 ();
 FILLCELL_X4 FILLER_149_1312 ();
 FILLCELL_X1 FILLER_149_1318 ();
 FILLCELL_X1 FILLER_149_1327 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X2 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_468 ();
 FILLCELL_X32 FILLER_150_500 ();
 FILLCELL_X32 FILLER_150_532 ();
 FILLCELL_X32 FILLER_150_564 ();
 FILLCELL_X32 FILLER_150_596 ();
 FILLCELL_X2 FILLER_150_628 ();
 FILLCELL_X1 FILLER_150_630 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X8 FILLER_150_1304 ();
 FILLCELL_X2 FILLER_150_1312 ();
 FILLCELL_X1 FILLER_150_1324 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X16 FILLER_151_193 ();
 FILLCELL_X8 FILLER_151_209 ();
 FILLCELL_X32 FILLER_151_230 ();
 FILLCELL_X32 FILLER_151_262 ();
 FILLCELL_X32 FILLER_151_294 ();
 FILLCELL_X32 FILLER_151_326 ();
 FILLCELL_X32 FILLER_151_358 ();
 FILLCELL_X32 FILLER_151_390 ();
 FILLCELL_X32 FILLER_151_422 ();
 FILLCELL_X8 FILLER_151_454 ();
 FILLCELL_X4 FILLER_151_462 ();
 FILLCELL_X1 FILLER_151_470 ();
 FILLCELL_X8 FILLER_151_488 ();
 FILLCELL_X2 FILLER_151_496 ();
 FILLCELL_X2 FILLER_151_532 ();
 FILLCELL_X1 FILLER_151_534 ();
 FILLCELL_X32 FILLER_151_552 ();
 FILLCELL_X32 FILLER_151_584 ();
 FILLCELL_X32 FILLER_151_616 ();
 FILLCELL_X32 FILLER_151_648 ();
 FILLCELL_X32 FILLER_151_680 ();
 FILLCELL_X32 FILLER_151_712 ();
 FILLCELL_X32 FILLER_151_744 ();
 FILLCELL_X32 FILLER_151_776 ();
 FILLCELL_X32 FILLER_151_808 ();
 FILLCELL_X32 FILLER_151_840 ();
 FILLCELL_X32 FILLER_151_872 ();
 FILLCELL_X32 FILLER_151_904 ();
 FILLCELL_X32 FILLER_151_936 ();
 FILLCELL_X32 FILLER_151_968 ();
 FILLCELL_X32 FILLER_151_1000 ();
 FILLCELL_X32 FILLER_151_1032 ();
 FILLCELL_X32 FILLER_151_1064 ();
 FILLCELL_X32 FILLER_151_1096 ();
 FILLCELL_X32 FILLER_151_1128 ();
 FILLCELL_X32 FILLER_151_1160 ();
 FILLCELL_X32 FILLER_151_1192 ();
 FILLCELL_X32 FILLER_151_1224 ();
 FILLCELL_X4 FILLER_151_1256 ();
 FILLCELL_X2 FILLER_151_1260 ();
 FILLCELL_X1 FILLER_151_1262 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X8 FILLER_151_1296 ();
 FILLCELL_X1 FILLER_151_1304 ();
 FILLCELL_X8 FILLER_151_1308 ();
 FILLCELL_X2 FILLER_151_1316 ();
 FILLCELL_X1 FILLER_151_1318 ();
 FILLCELL_X1 FILLER_151_1321 ();
 FILLCELL_X1 FILLER_151_1325 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X4 FILLER_152_385 ();
 FILLCELL_X2 FILLER_152_389 ();
 FILLCELL_X1 FILLER_152_391 ();
 FILLCELL_X16 FILLER_152_409 ();
 FILLCELL_X8 FILLER_152_425 ();
 FILLCELL_X16 FILLER_152_450 ();
 FILLCELL_X1 FILLER_152_466 ();
 FILLCELL_X2 FILLER_152_474 ();
 FILLCELL_X1 FILLER_152_476 ();
 FILLCELL_X4 FILLER_152_479 ();
 FILLCELL_X2 FILLER_152_483 ();
 FILLCELL_X16 FILLER_152_489 ();
 FILLCELL_X2 FILLER_152_505 ();
 FILLCELL_X1 FILLER_152_507 ();
 FILLCELL_X2 FILLER_152_512 ();
 FILLCELL_X1 FILLER_152_514 ();
 FILLCELL_X2 FILLER_152_518 ();
 FILLCELL_X1 FILLER_152_520 ();
 FILLCELL_X2 FILLER_152_525 ();
 FILLCELL_X1 FILLER_152_527 ();
 FILLCELL_X4 FILLER_152_532 ();
 FILLCELL_X1 FILLER_152_536 ();
 FILLCELL_X32 FILLER_152_548 ();
 FILLCELL_X32 FILLER_152_580 ();
 FILLCELL_X16 FILLER_152_612 ();
 FILLCELL_X2 FILLER_152_628 ();
 FILLCELL_X1 FILLER_152_630 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X4 FILLER_152_1304 ();
 FILLCELL_X2 FILLER_152_1308 ();
 FILLCELL_X1 FILLER_152_1310 ();
 FILLCELL_X4 FILLER_152_1316 ();
 FILLCELL_X2 FILLER_152_1320 ();
 FILLCELL_X1 FILLER_152_1322 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X8 FILLER_153_385 ();
 FILLCELL_X4 FILLER_153_402 ();
 FILLCELL_X2 FILLER_153_406 ();
 FILLCELL_X8 FILLER_153_429 ();
 FILLCELL_X2 FILLER_153_437 ();
 FILLCELL_X1 FILLER_153_439 ();
 FILLCELL_X1 FILLER_153_447 ();
 FILLCELL_X16 FILLER_153_452 ();
 FILLCELL_X1 FILLER_153_475 ();
 FILLCELL_X16 FILLER_153_488 ();
 FILLCELL_X4 FILLER_153_504 ();
 FILLCELL_X2 FILLER_153_508 ();
 FILLCELL_X1 FILLER_153_510 ();
 FILLCELL_X4 FILLER_153_518 ();
 FILLCELL_X2 FILLER_153_522 ();
 FILLCELL_X2 FILLER_153_531 ();
 FILLCELL_X1 FILLER_153_533 ();
 FILLCELL_X4 FILLER_153_550 ();
 FILLCELL_X2 FILLER_153_554 ();
 FILLCELL_X1 FILLER_153_556 ();
 FILLCELL_X4 FILLER_153_574 ();
 FILLCELL_X2 FILLER_153_578 ();
 FILLCELL_X1 FILLER_153_580 ();
 FILLCELL_X32 FILLER_153_585 ();
 FILLCELL_X32 FILLER_153_617 ();
 FILLCELL_X32 FILLER_153_649 ();
 FILLCELL_X32 FILLER_153_681 ();
 FILLCELL_X32 FILLER_153_713 ();
 FILLCELL_X32 FILLER_153_745 ();
 FILLCELL_X32 FILLER_153_777 ();
 FILLCELL_X32 FILLER_153_809 ();
 FILLCELL_X32 FILLER_153_841 ();
 FILLCELL_X32 FILLER_153_873 ();
 FILLCELL_X32 FILLER_153_905 ();
 FILLCELL_X32 FILLER_153_937 ();
 FILLCELL_X32 FILLER_153_969 ();
 FILLCELL_X32 FILLER_153_1001 ();
 FILLCELL_X32 FILLER_153_1033 ();
 FILLCELL_X32 FILLER_153_1065 ();
 FILLCELL_X32 FILLER_153_1097 ();
 FILLCELL_X32 FILLER_153_1129 ();
 FILLCELL_X32 FILLER_153_1161 ();
 FILLCELL_X32 FILLER_153_1193 ();
 FILLCELL_X32 FILLER_153_1225 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X8 FILLER_153_1296 ();
 FILLCELL_X4 FILLER_153_1304 ();
 FILLCELL_X2 FILLER_153_1308 ();
 FILLCELL_X1 FILLER_153_1310 ();
 FILLCELL_X1 FILLER_153_1318 ();
 FILLCELL_X1 FILLER_153_1324 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X8 FILLER_154_385 ();
 FILLCELL_X1 FILLER_154_393 ();
 FILLCELL_X8 FILLER_154_402 ();
 FILLCELL_X2 FILLER_154_410 ();
 FILLCELL_X1 FILLER_154_412 ();
 FILLCELL_X2 FILLER_154_416 ();
 FILLCELL_X1 FILLER_154_418 ();
 FILLCELL_X16 FILLER_154_423 ();
 FILLCELL_X1 FILLER_154_439 ();
 FILLCELL_X32 FILLER_154_450 ();
 FILLCELL_X16 FILLER_154_482 ();
 FILLCELL_X8 FILLER_154_498 ();
 FILLCELL_X4 FILLER_154_506 ();
 FILLCELL_X2 FILLER_154_510 ();
 FILLCELL_X1 FILLER_154_512 ();
 FILLCELL_X16 FILLER_154_534 ();
 FILLCELL_X8 FILLER_154_550 ();
 FILLCELL_X4 FILLER_154_558 ();
 FILLCELL_X1 FILLER_154_562 ();
 FILLCELL_X2 FILLER_154_567 ();
 FILLCELL_X1 FILLER_154_569 ();
 FILLCELL_X1 FILLER_154_576 ();
 FILLCELL_X16 FILLER_154_612 ();
 FILLCELL_X2 FILLER_154_628 ();
 FILLCELL_X1 FILLER_154_630 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X8 FILLER_154_1304 ();
 FILLCELL_X2 FILLER_154_1312 ();
 FILLCELL_X1 FILLER_154_1314 ();
 FILLCELL_X2 FILLER_154_1320 ();
 FILLCELL_X1 FILLER_154_1322 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X4 FILLER_155_396 ();
 FILLCELL_X2 FILLER_155_400 ();
 FILLCELL_X32 FILLER_155_415 ();
 FILLCELL_X16 FILLER_155_447 ();
 FILLCELL_X8 FILLER_155_463 ();
 FILLCELL_X4 FILLER_155_471 ();
 FILLCELL_X16 FILLER_155_496 ();
 FILLCELL_X4 FILLER_155_512 ();
 FILLCELL_X2 FILLER_155_516 ();
 FILLCELL_X1 FILLER_155_518 ();
 FILLCELL_X4 FILLER_155_535 ();
 FILLCELL_X8 FILLER_155_544 ();
 FILLCELL_X4 FILLER_155_552 ();
 FILLCELL_X2 FILLER_155_556 ();
 FILLCELL_X1 FILLER_155_558 ();
 FILLCELL_X4 FILLER_155_567 ();
 FILLCELL_X2 FILLER_155_571 ();
 FILLCELL_X1 FILLER_155_573 ();
 FILLCELL_X32 FILLER_155_589 ();
 FILLCELL_X32 FILLER_155_621 ();
 FILLCELL_X32 FILLER_155_653 ();
 FILLCELL_X32 FILLER_155_685 ();
 FILLCELL_X32 FILLER_155_717 ();
 FILLCELL_X32 FILLER_155_749 ();
 FILLCELL_X32 FILLER_155_781 ();
 FILLCELL_X32 FILLER_155_813 ();
 FILLCELL_X32 FILLER_155_845 ();
 FILLCELL_X32 FILLER_155_877 ();
 FILLCELL_X32 FILLER_155_909 ();
 FILLCELL_X32 FILLER_155_941 ();
 FILLCELL_X32 FILLER_155_973 ();
 FILLCELL_X32 FILLER_155_1005 ();
 FILLCELL_X32 FILLER_155_1037 ();
 FILLCELL_X32 FILLER_155_1069 ();
 FILLCELL_X32 FILLER_155_1101 ();
 FILLCELL_X32 FILLER_155_1133 ();
 FILLCELL_X32 FILLER_155_1165 ();
 FILLCELL_X32 FILLER_155_1197 ();
 FILLCELL_X32 FILLER_155_1229 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X8 FILLER_155_1296 ();
 FILLCELL_X4 FILLER_155_1304 ();
 FILLCELL_X2 FILLER_155_1311 ();
 FILLCELL_X1 FILLER_155_1313 ();
 FILLCELL_X2 FILLER_155_1319 ();
 FILLCELL_X2 FILLER_155_1326 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X16 FILLER_156_353 ();
 FILLCELL_X4 FILLER_156_373 ();
 FILLCELL_X2 FILLER_156_377 ();
 FILLCELL_X2 FILLER_156_389 ();
 FILLCELL_X1 FILLER_156_391 ();
 FILLCELL_X8 FILLER_156_413 ();
 FILLCELL_X4 FILLER_156_421 ();
 FILLCELL_X1 FILLER_156_425 ();
 FILLCELL_X16 FILLER_156_429 ();
 FILLCELL_X2 FILLER_156_454 ();
 FILLCELL_X1 FILLER_156_480 ();
 FILLCELL_X8 FILLER_156_486 ();
 FILLCELL_X4 FILLER_156_494 ();
 FILLCELL_X1 FILLER_156_498 ();
 FILLCELL_X8 FILLER_156_506 ();
 FILLCELL_X2 FILLER_156_514 ();
 FILLCELL_X2 FILLER_156_528 ();
 FILLCELL_X16 FILLER_156_535 ();
 FILLCELL_X4 FILLER_156_551 ();
 FILLCELL_X2 FILLER_156_555 ();
 FILLCELL_X1 FILLER_156_557 ();
 FILLCELL_X32 FILLER_156_565 ();
 FILLCELL_X16 FILLER_156_597 ();
 FILLCELL_X8 FILLER_156_613 ();
 FILLCELL_X2 FILLER_156_621 ();
 FILLCELL_X2 FILLER_156_628 ();
 FILLCELL_X1 FILLER_156_630 ();
 FILLCELL_X32 FILLER_156_637 ();
 FILLCELL_X32 FILLER_156_669 ();
 FILLCELL_X32 FILLER_156_701 ();
 FILLCELL_X32 FILLER_156_733 ();
 FILLCELL_X32 FILLER_156_765 ();
 FILLCELL_X32 FILLER_156_797 ();
 FILLCELL_X32 FILLER_156_829 ();
 FILLCELL_X32 FILLER_156_861 ();
 FILLCELL_X32 FILLER_156_893 ();
 FILLCELL_X32 FILLER_156_925 ();
 FILLCELL_X32 FILLER_156_957 ();
 FILLCELL_X32 FILLER_156_989 ();
 FILLCELL_X32 FILLER_156_1021 ();
 FILLCELL_X32 FILLER_156_1053 ();
 FILLCELL_X32 FILLER_156_1085 ();
 FILLCELL_X32 FILLER_156_1117 ();
 FILLCELL_X32 FILLER_156_1149 ();
 FILLCELL_X32 FILLER_156_1181 ();
 FILLCELL_X32 FILLER_156_1213 ();
 FILLCELL_X32 FILLER_156_1245 ();
 FILLCELL_X32 FILLER_156_1277 ();
 FILLCELL_X1 FILLER_156_1309 ();
 FILLCELL_X4 FILLER_156_1313 ();
 FILLCELL_X1 FILLER_156_1324 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X16 FILLER_157_353 ();
 FILLCELL_X1 FILLER_157_369 ();
 FILLCELL_X16 FILLER_157_377 ();
 FILLCELL_X2 FILLER_157_393 ();
 FILLCELL_X2 FILLER_157_403 ();
 FILLCELL_X1 FILLER_157_405 ();
 FILLCELL_X2 FILLER_157_413 ();
 FILLCELL_X32 FILLER_157_425 ();
 FILLCELL_X4 FILLER_157_457 ();
 FILLCELL_X2 FILLER_157_470 ();
 FILLCELL_X1 FILLER_157_472 ();
 FILLCELL_X1 FILLER_157_478 ();
 FILLCELL_X16 FILLER_157_489 ();
 FILLCELL_X1 FILLER_157_505 ();
 FILLCELL_X16 FILLER_157_534 ();
 FILLCELL_X4 FILLER_157_550 ();
 FILLCELL_X2 FILLER_157_554 ();
 FILLCELL_X1 FILLER_157_556 ();
 FILLCELL_X2 FILLER_157_567 ();
 FILLCELL_X1 FILLER_157_569 ();
 FILLCELL_X1 FILLER_157_573 ();
 FILLCELL_X2 FILLER_157_581 ();
 FILLCELL_X32 FILLER_157_587 ();
 FILLCELL_X32 FILLER_157_619 ();
 FILLCELL_X32 FILLER_157_651 ();
 FILLCELL_X32 FILLER_157_683 ();
 FILLCELL_X32 FILLER_157_715 ();
 FILLCELL_X32 FILLER_157_747 ();
 FILLCELL_X32 FILLER_157_779 ();
 FILLCELL_X32 FILLER_157_811 ();
 FILLCELL_X32 FILLER_157_843 ();
 FILLCELL_X32 FILLER_157_875 ();
 FILLCELL_X32 FILLER_157_907 ();
 FILLCELL_X32 FILLER_157_939 ();
 FILLCELL_X32 FILLER_157_971 ();
 FILLCELL_X32 FILLER_157_1003 ();
 FILLCELL_X32 FILLER_157_1035 ();
 FILLCELL_X32 FILLER_157_1067 ();
 FILLCELL_X32 FILLER_157_1099 ();
 FILLCELL_X32 FILLER_157_1131 ();
 FILLCELL_X32 FILLER_157_1163 ();
 FILLCELL_X32 FILLER_157_1195 ();
 FILLCELL_X32 FILLER_157_1227 ();
 FILLCELL_X4 FILLER_157_1259 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X16 FILLER_157_1296 ();
 FILLCELL_X2 FILLER_157_1312 ();
 FILLCELL_X1 FILLER_157_1319 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X16 FILLER_158_321 ();
 FILLCELL_X4 FILLER_158_337 ();
 FILLCELL_X1 FILLER_158_362 ();
 FILLCELL_X4 FILLER_158_372 ();
 FILLCELL_X2 FILLER_158_376 ();
 FILLCELL_X1 FILLER_158_378 ();
 FILLCELL_X1 FILLER_158_387 ();
 FILLCELL_X32 FILLER_158_393 ();
 FILLCELL_X32 FILLER_158_425 ();
 FILLCELL_X2 FILLER_158_461 ();
 FILLCELL_X1 FILLER_158_463 ();
 FILLCELL_X2 FILLER_158_494 ();
 FILLCELL_X1 FILLER_158_501 ();
 FILLCELL_X8 FILLER_158_520 ();
 FILLCELL_X4 FILLER_158_528 ();
 FILLCELL_X2 FILLER_158_539 ();
 FILLCELL_X16 FILLER_158_545 ();
 FILLCELL_X4 FILLER_158_561 ();
 FILLCELL_X1 FILLER_158_565 ();
 FILLCELL_X4 FILLER_158_573 ();
 FILLCELL_X4 FILLER_158_588 ();
 FILLCELL_X1 FILLER_158_592 ();
 FILLCELL_X8 FILLER_158_617 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X16 FILLER_158_1304 ();
 FILLCELL_X2 FILLER_158_1320 ();
 FILLCELL_X1 FILLER_158_1322 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X16 FILLER_159_321 ();
 FILLCELL_X2 FILLER_159_337 ();
 FILLCELL_X1 FILLER_159_339 ();
 FILLCELL_X4 FILLER_159_343 ();
 FILLCELL_X1 FILLER_159_347 ();
 FILLCELL_X8 FILLER_159_358 ();
 FILLCELL_X4 FILLER_159_366 ();
 FILLCELL_X32 FILLER_159_376 ();
 FILLCELL_X2 FILLER_159_408 ();
 FILLCELL_X1 FILLER_159_410 ();
 FILLCELL_X8 FILLER_159_429 ();
 FILLCELL_X4 FILLER_159_437 ();
 FILLCELL_X1 FILLER_159_458 ();
 FILLCELL_X1 FILLER_159_474 ();
 FILLCELL_X8 FILLER_159_481 ();
 FILLCELL_X1 FILLER_159_489 ();
 FILLCELL_X16 FILLER_159_510 ();
 FILLCELL_X8 FILLER_159_526 ();
 FILLCELL_X2 FILLER_159_534 ();
 FILLCELL_X1 FILLER_159_536 ();
 FILLCELL_X16 FILLER_159_544 ();
 FILLCELL_X8 FILLER_159_560 ();
 FILLCELL_X2 FILLER_159_568 ();
 FILLCELL_X16 FILLER_159_574 ();
 FILLCELL_X32 FILLER_159_600 ();
 FILLCELL_X32 FILLER_159_632 ();
 FILLCELL_X32 FILLER_159_664 ();
 FILLCELL_X32 FILLER_159_696 ();
 FILLCELL_X32 FILLER_159_728 ();
 FILLCELL_X32 FILLER_159_760 ();
 FILLCELL_X32 FILLER_159_792 ();
 FILLCELL_X32 FILLER_159_824 ();
 FILLCELL_X32 FILLER_159_856 ();
 FILLCELL_X32 FILLER_159_888 ();
 FILLCELL_X32 FILLER_159_920 ();
 FILLCELL_X32 FILLER_159_952 ();
 FILLCELL_X32 FILLER_159_984 ();
 FILLCELL_X32 FILLER_159_1016 ();
 FILLCELL_X32 FILLER_159_1048 ();
 FILLCELL_X32 FILLER_159_1080 ();
 FILLCELL_X32 FILLER_159_1112 ();
 FILLCELL_X32 FILLER_159_1144 ();
 FILLCELL_X32 FILLER_159_1176 ();
 FILLCELL_X32 FILLER_159_1208 ();
 FILLCELL_X16 FILLER_159_1240 ();
 FILLCELL_X4 FILLER_159_1256 ();
 FILLCELL_X2 FILLER_159_1260 ();
 FILLCELL_X1 FILLER_159_1262 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X16 FILLER_159_1296 ();
 FILLCELL_X2 FILLER_159_1312 ();
 FILLCELL_X1 FILLER_159_1314 ();
 FILLCELL_X8 FILLER_159_1320 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X4 FILLER_160_321 ();
 FILLCELL_X1 FILLER_160_325 ();
 FILLCELL_X1 FILLER_160_350 ();
 FILLCELL_X2 FILLER_160_356 ();
 FILLCELL_X2 FILLER_160_362 ();
 FILLCELL_X1 FILLER_160_364 ();
 FILLCELL_X4 FILLER_160_386 ();
 FILLCELL_X4 FILLER_160_401 ();
 FILLCELL_X2 FILLER_160_405 ();
 FILLCELL_X32 FILLER_160_425 ();
 FILLCELL_X4 FILLER_160_457 ();
 FILLCELL_X2 FILLER_160_461 ();
 FILLCELL_X32 FILLER_160_487 ();
 FILLCELL_X8 FILLER_160_519 ();
 FILLCELL_X1 FILLER_160_527 ();
 FILLCELL_X16 FILLER_160_555 ();
 FILLCELL_X2 FILLER_160_571 ();
 FILLCELL_X1 FILLER_160_581 ();
 FILLCELL_X32 FILLER_160_592 ();
 FILLCELL_X4 FILLER_160_624 ();
 FILLCELL_X2 FILLER_160_628 ();
 FILLCELL_X1 FILLER_160_630 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X16 FILLER_160_1304 ();
 FILLCELL_X8 FILLER_160_1320 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X2 FILLER_161_353 ();
 FILLCELL_X1 FILLER_161_355 ();
 FILLCELL_X1 FILLER_161_361 ();
 FILLCELL_X8 FILLER_161_380 ();
 FILLCELL_X4 FILLER_161_388 ();
 FILLCELL_X2 FILLER_161_392 ();
 FILLCELL_X8 FILLER_161_403 ();
 FILLCELL_X2 FILLER_161_411 ();
 FILLCELL_X32 FILLER_161_426 ();
 FILLCELL_X4 FILLER_161_458 ();
 FILLCELL_X2 FILLER_161_462 ();
 FILLCELL_X32 FILLER_161_469 ();
 FILLCELL_X16 FILLER_161_501 ();
 FILLCELL_X8 FILLER_161_517 ();
 FILLCELL_X2 FILLER_161_525 ();
 FILLCELL_X1 FILLER_161_527 ();
 FILLCELL_X32 FILLER_161_542 ();
 FILLCELL_X2 FILLER_161_574 ();
 FILLCELL_X1 FILLER_161_576 ();
 FILLCELL_X32 FILLER_161_602 ();
 FILLCELL_X32 FILLER_161_634 ();
 FILLCELL_X32 FILLER_161_666 ();
 FILLCELL_X32 FILLER_161_698 ();
 FILLCELL_X32 FILLER_161_730 ();
 FILLCELL_X32 FILLER_161_762 ();
 FILLCELL_X32 FILLER_161_794 ();
 FILLCELL_X32 FILLER_161_826 ();
 FILLCELL_X32 FILLER_161_858 ();
 FILLCELL_X32 FILLER_161_890 ();
 FILLCELL_X32 FILLER_161_922 ();
 FILLCELL_X32 FILLER_161_954 ();
 FILLCELL_X32 FILLER_161_986 ();
 FILLCELL_X32 FILLER_161_1018 ();
 FILLCELL_X32 FILLER_161_1050 ();
 FILLCELL_X32 FILLER_161_1082 ();
 FILLCELL_X32 FILLER_161_1114 ();
 FILLCELL_X32 FILLER_161_1146 ();
 FILLCELL_X32 FILLER_161_1178 ();
 FILLCELL_X32 FILLER_161_1210 ();
 FILLCELL_X16 FILLER_161_1242 ();
 FILLCELL_X4 FILLER_161_1258 ();
 FILLCELL_X1 FILLER_161_1262 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X16 FILLER_162_321 ();
 FILLCELL_X8 FILLER_162_337 ();
 FILLCELL_X4 FILLER_162_345 ();
 FILLCELL_X8 FILLER_162_372 ();
 FILLCELL_X4 FILLER_162_380 ();
 FILLCELL_X2 FILLER_162_384 ();
 FILLCELL_X1 FILLER_162_386 ();
 FILLCELL_X16 FILLER_162_395 ();
 FILLCELL_X4 FILLER_162_411 ();
 FILLCELL_X2 FILLER_162_415 ();
 FILLCELL_X32 FILLER_162_440 ();
 FILLCELL_X32 FILLER_162_472 ();
 FILLCELL_X16 FILLER_162_504 ();
 FILLCELL_X2 FILLER_162_520 ();
 FILLCELL_X1 FILLER_162_522 ();
 FILLCELL_X32 FILLER_162_525 ();
 FILLCELL_X32 FILLER_162_557 ();
 FILLCELL_X2 FILLER_162_589 ();
 FILLCELL_X1 FILLER_162_591 ();
 FILLCELL_X32 FILLER_162_597 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X16 FILLER_162_1304 ();
 FILLCELL_X8 FILLER_162_1320 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X8 FILLER_163_321 ();
 FILLCELL_X4 FILLER_163_329 ();
 FILLCELL_X2 FILLER_163_333 ();
 FILLCELL_X1 FILLER_163_335 ();
 FILLCELL_X32 FILLER_163_368 ();
 FILLCELL_X8 FILLER_163_400 ();
 FILLCELL_X4 FILLER_163_408 ();
 FILLCELL_X1 FILLER_163_412 ();
 FILLCELL_X4 FILLER_163_441 ();
 FILLCELL_X1 FILLER_163_445 ();
 FILLCELL_X2 FILLER_163_449 ();
 FILLCELL_X1 FILLER_163_451 ();
 FILLCELL_X1 FILLER_163_459 ();
 FILLCELL_X1 FILLER_163_462 ();
 FILLCELL_X1 FILLER_163_472 ();
 FILLCELL_X4 FILLER_163_480 ();
 FILLCELL_X4 FILLER_163_503 ();
 FILLCELL_X2 FILLER_163_529 ();
 FILLCELL_X1 FILLER_163_531 ();
 FILLCELL_X32 FILLER_163_542 ();
 FILLCELL_X32 FILLER_163_574 ();
 FILLCELL_X32 FILLER_163_606 ();
 FILLCELL_X32 FILLER_163_638 ();
 FILLCELL_X32 FILLER_163_670 ();
 FILLCELL_X32 FILLER_163_702 ();
 FILLCELL_X32 FILLER_163_734 ();
 FILLCELL_X32 FILLER_163_766 ();
 FILLCELL_X32 FILLER_163_798 ();
 FILLCELL_X32 FILLER_163_830 ();
 FILLCELL_X32 FILLER_163_862 ();
 FILLCELL_X32 FILLER_163_894 ();
 FILLCELL_X32 FILLER_163_926 ();
 FILLCELL_X32 FILLER_163_958 ();
 FILLCELL_X32 FILLER_163_990 ();
 FILLCELL_X32 FILLER_163_1022 ();
 FILLCELL_X32 FILLER_163_1054 ();
 FILLCELL_X32 FILLER_163_1086 ();
 FILLCELL_X32 FILLER_163_1118 ();
 FILLCELL_X32 FILLER_163_1150 ();
 FILLCELL_X32 FILLER_163_1182 ();
 FILLCELL_X32 FILLER_163_1214 ();
 FILLCELL_X16 FILLER_163_1246 ();
 FILLCELL_X1 FILLER_163_1262 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X16 FILLER_164_225 ();
 FILLCELL_X8 FILLER_164_241 ();
 FILLCELL_X4 FILLER_164_249 ();
 FILLCELL_X32 FILLER_164_260 ();
 FILLCELL_X32 FILLER_164_292 ();
 FILLCELL_X32 FILLER_164_324 ();
 FILLCELL_X2 FILLER_164_360 ();
 FILLCELL_X1 FILLER_164_362 ();
 FILLCELL_X16 FILLER_164_370 ();
 FILLCELL_X4 FILLER_164_386 ();
 FILLCELL_X32 FILLER_164_407 ();
 FILLCELL_X4 FILLER_164_439 ();
 FILLCELL_X4 FILLER_164_453 ();
 FILLCELL_X2 FILLER_164_457 ();
 FILLCELL_X4 FILLER_164_464 ();
 FILLCELL_X2 FILLER_164_468 ();
 FILLCELL_X1 FILLER_164_470 ();
 FILLCELL_X2 FILLER_164_475 ();
 FILLCELL_X1 FILLER_164_477 ();
 FILLCELL_X32 FILLER_164_493 ();
 FILLCELL_X16 FILLER_164_525 ();
 FILLCELL_X8 FILLER_164_541 ();
 FILLCELL_X8 FILLER_164_575 ();
 FILLCELL_X4 FILLER_164_583 ();
 FILLCELL_X2 FILLER_164_587 ();
 FILLCELL_X16 FILLER_164_612 ();
 FILLCELL_X2 FILLER_164_628 ();
 FILLCELL_X1 FILLER_164_630 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X16 FILLER_164_1304 ();
 FILLCELL_X8 FILLER_164_1320 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X2 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_240 ();
 FILLCELL_X32 FILLER_165_272 ();
 FILLCELL_X16 FILLER_165_304 ();
 FILLCELL_X1 FILLER_165_320 ();
 FILLCELL_X4 FILLER_165_342 ();
 FILLCELL_X1 FILLER_165_346 ();
 FILLCELL_X16 FILLER_165_372 ();
 FILLCELL_X8 FILLER_165_388 ();
 FILLCELL_X2 FILLER_165_396 ();
 FILLCELL_X16 FILLER_165_411 ();
 FILLCELL_X2 FILLER_165_427 ();
 FILLCELL_X16 FILLER_165_434 ();
 FILLCELL_X4 FILLER_165_450 ();
 FILLCELL_X4 FILLER_165_471 ();
 FILLCELL_X32 FILLER_165_478 ();
 FILLCELL_X4 FILLER_165_510 ();
 FILLCELL_X2 FILLER_165_514 ();
 FILLCELL_X1 FILLER_165_516 ();
 FILLCELL_X8 FILLER_165_521 ();
 FILLCELL_X8 FILLER_165_531 ();
 FILLCELL_X2 FILLER_165_543 ();
 FILLCELL_X16 FILLER_165_578 ();
 FILLCELL_X8 FILLER_165_594 ();
 FILLCELL_X4 FILLER_165_602 ();
 FILLCELL_X2 FILLER_165_606 ();
 FILLCELL_X4 FILLER_165_612 ();
 FILLCELL_X1 FILLER_165_616 ();
 FILLCELL_X4 FILLER_165_636 ();
 FILLCELL_X1 FILLER_165_640 ();
 FILLCELL_X32 FILLER_165_644 ();
 FILLCELL_X32 FILLER_165_676 ();
 FILLCELL_X32 FILLER_165_708 ();
 FILLCELL_X32 FILLER_165_740 ();
 FILLCELL_X32 FILLER_165_772 ();
 FILLCELL_X32 FILLER_165_804 ();
 FILLCELL_X32 FILLER_165_836 ();
 FILLCELL_X32 FILLER_165_868 ();
 FILLCELL_X32 FILLER_165_900 ();
 FILLCELL_X32 FILLER_165_932 ();
 FILLCELL_X32 FILLER_165_964 ();
 FILLCELL_X32 FILLER_165_996 ();
 FILLCELL_X32 FILLER_165_1028 ();
 FILLCELL_X32 FILLER_165_1060 ();
 FILLCELL_X32 FILLER_165_1092 ();
 FILLCELL_X32 FILLER_165_1124 ();
 FILLCELL_X32 FILLER_165_1156 ();
 FILLCELL_X32 FILLER_165_1188 ();
 FILLCELL_X32 FILLER_165_1220 ();
 FILLCELL_X8 FILLER_165_1252 ();
 FILLCELL_X2 FILLER_165_1260 ();
 FILLCELL_X1 FILLER_165_1262 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X4 FILLER_166_321 ();
 FILLCELL_X1 FILLER_166_325 ();
 FILLCELL_X4 FILLER_166_347 ();
 FILLCELL_X1 FILLER_166_372 ();
 FILLCELL_X16 FILLER_166_375 ();
 FILLCELL_X4 FILLER_166_391 ();
 FILLCELL_X2 FILLER_166_395 ();
 FILLCELL_X32 FILLER_166_405 ();
 FILLCELL_X16 FILLER_166_437 ();
 FILLCELL_X8 FILLER_166_453 ();
 FILLCELL_X1 FILLER_166_461 ();
 FILLCELL_X4 FILLER_166_468 ();
 FILLCELL_X16 FILLER_166_483 ();
 FILLCELL_X8 FILLER_166_499 ();
 FILLCELL_X4 FILLER_166_507 ();
 FILLCELL_X2 FILLER_166_511 ();
 FILLCELL_X16 FILLER_166_532 ();
 FILLCELL_X8 FILLER_166_548 ();
 FILLCELL_X4 FILLER_166_556 ();
 FILLCELL_X2 FILLER_166_560 ();
 FILLCELL_X1 FILLER_166_562 ();
 FILLCELL_X1 FILLER_166_569 ();
 FILLCELL_X16 FILLER_166_592 ();
 FILLCELL_X8 FILLER_166_608 ();
 FILLCELL_X2 FILLER_166_616 ();
 FILLCELL_X2 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_649 ();
 FILLCELL_X32 FILLER_166_681 ();
 FILLCELL_X32 FILLER_166_713 ();
 FILLCELL_X32 FILLER_166_745 ();
 FILLCELL_X32 FILLER_166_777 ();
 FILLCELL_X32 FILLER_166_809 ();
 FILLCELL_X32 FILLER_166_841 ();
 FILLCELL_X32 FILLER_166_873 ();
 FILLCELL_X32 FILLER_166_905 ();
 FILLCELL_X32 FILLER_166_937 ();
 FILLCELL_X32 FILLER_166_969 ();
 FILLCELL_X32 FILLER_166_1001 ();
 FILLCELL_X32 FILLER_166_1033 ();
 FILLCELL_X32 FILLER_166_1065 ();
 FILLCELL_X32 FILLER_166_1097 ();
 FILLCELL_X32 FILLER_166_1129 ();
 FILLCELL_X32 FILLER_166_1161 ();
 FILLCELL_X32 FILLER_166_1193 ();
 FILLCELL_X32 FILLER_166_1225 ();
 FILLCELL_X32 FILLER_166_1257 ();
 FILLCELL_X32 FILLER_166_1289 ();
 FILLCELL_X4 FILLER_166_1321 ();
 FILLCELL_X2 FILLER_166_1325 ();
 FILLCELL_X1 FILLER_166_1327 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X4 FILLER_167_353 ();
 FILLCELL_X8 FILLER_167_370 ();
 FILLCELL_X4 FILLER_167_378 ();
 FILLCELL_X2 FILLER_167_382 ();
 FILLCELL_X1 FILLER_167_384 ();
 FILLCELL_X2 FILLER_167_411 ();
 FILLCELL_X1 FILLER_167_413 ();
 FILLCELL_X32 FILLER_167_424 ();
 FILLCELL_X16 FILLER_167_456 ();
 FILLCELL_X1 FILLER_167_472 ();
 FILLCELL_X16 FILLER_167_490 ();
 FILLCELL_X4 FILLER_167_506 ();
 FILLCELL_X2 FILLER_167_510 ();
 FILLCELL_X1 FILLER_167_530 ();
 FILLCELL_X16 FILLER_167_548 ();
 FILLCELL_X1 FILLER_167_564 ();
 FILLCELL_X32 FILLER_167_572 ();
 FILLCELL_X16 FILLER_167_604 ();
 FILLCELL_X2 FILLER_167_620 ();
 FILLCELL_X1 FILLER_167_622 ();
 FILLCELL_X8 FILLER_167_627 ();
 FILLCELL_X32 FILLER_167_652 ();
 FILLCELL_X32 FILLER_167_684 ();
 FILLCELL_X32 FILLER_167_716 ();
 FILLCELL_X32 FILLER_167_748 ();
 FILLCELL_X32 FILLER_167_780 ();
 FILLCELL_X32 FILLER_167_812 ();
 FILLCELL_X32 FILLER_167_844 ();
 FILLCELL_X32 FILLER_167_876 ();
 FILLCELL_X32 FILLER_167_908 ();
 FILLCELL_X32 FILLER_167_940 ();
 FILLCELL_X32 FILLER_167_972 ();
 FILLCELL_X32 FILLER_167_1004 ();
 FILLCELL_X32 FILLER_167_1036 ();
 FILLCELL_X32 FILLER_167_1068 ();
 FILLCELL_X32 FILLER_167_1100 ();
 FILLCELL_X32 FILLER_167_1132 ();
 FILLCELL_X32 FILLER_167_1164 ();
 FILLCELL_X32 FILLER_167_1196 ();
 FILLCELL_X32 FILLER_167_1228 ();
 FILLCELL_X2 FILLER_167_1260 ();
 FILLCELL_X1 FILLER_167_1262 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X4 FILLER_168_353 ();
 FILLCELL_X4 FILLER_168_361 ();
 FILLCELL_X2 FILLER_168_370 ();
 FILLCELL_X1 FILLER_168_372 ();
 FILLCELL_X16 FILLER_168_379 ();
 FILLCELL_X4 FILLER_168_395 ();
 FILLCELL_X2 FILLER_168_399 ();
 FILLCELL_X1 FILLER_168_401 ();
 FILLCELL_X2 FILLER_168_437 ();
 FILLCELL_X32 FILLER_168_446 ();
 FILLCELL_X32 FILLER_168_478 ();
 FILLCELL_X32 FILLER_168_510 ();
 FILLCELL_X8 FILLER_168_542 ();
 FILLCELL_X4 FILLER_168_550 ();
 FILLCELL_X2 FILLER_168_560 ();
 FILLCELL_X32 FILLER_168_576 ();
 FILLCELL_X16 FILLER_168_608 ();
 FILLCELL_X4 FILLER_168_624 ();
 FILLCELL_X2 FILLER_168_628 ();
 FILLCELL_X1 FILLER_168_630 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X32 FILLER_168_1176 ();
 FILLCELL_X32 FILLER_168_1208 ();
 FILLCELL_X32 FILLER_168_1240 ();
 FILLCELL_X32 FILLER_168_1272 ();
 FILLCELL_X16 FILLER_168_1304 ();
 FILLCELL_X8 FILLER_168_1320 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X4 FILLER_169_353 ();
 FILLCELL_X1 FILLER_169_357 ();
 FILLCELL_X32 FILLER_169_372 ();
 FILLCELL_X4 FILLER_169_404 ();
 FILLCELL_X1 FILLER_169_408 ();
 FILLCELL_X4 FILLER_169_427 ();
 FILLCELL_X2 FILLER_169_431 ();
 FILLCELL_X1 FILLER_169_433 ();
 FILLCELL_X32 FILLER_169_453 ();
 FILLCELL_X16 FILLER_169_485 ();
 FILLCELL_X8 FILLER_169_501 ();
 FILLCELL_X4 FILLER_169_509 ();
 FILLCELL_X2 FILLER_169_513 ();
 FILLCELL_X1 FILLER_169_515 ();
 FILLCELL_X16 FILLER_169_523 ();
 FILLCELL_X8 FILLER_169_539 ();
 FILLCELL_X2 FILLER_169_547 ();
 FILLCELL_X8 FILLER_169_556 ();
 FILLCELL_X4 FILLER_169_564 ();
 FILLCELL_X4 FILLER_169_582 ();
 FILLCELL_X32 FILLER_169_589 ();
 FILLCELL_X16 FILLER_169_621 ();
 FILLCELL_X4 FILLER_169_637 ();
 FILLCELL_X32 FILLER_169_645 ();
 FILLCELL_X32 FILLER_169_677 ();
 FILLCELL_X32 FILLER_169_709 ();
 FILLCELL_X32 FILLER_169_741 ();
 FILLCELL_X32 FILLER_169_773 ();
 FILLCELL_X32 FILLER_169_805 ();
 FILLCELL_X32 FILLER_169_837 ();
 FILLCELL_X32 FILLER_169_869 ();
 FILLCELL_X32 FILLER_169_901 ();
 FILLCELL_X32 FILLER_169_933 ();
 FILLCELL_X32 FILLER_169_965 ();
 FILLCELL_X32 FILLER_169_997 ();
 FILLCELL_X32 FILLER_169_1029 ();
 FILLCELL_X32 FILLER_169_1061 ();
 FILLCELL_X32 FILLER_169_1093 ();
 FILLCELL_X32 FILLER_169_1125 ();
 FILLCELL_X32 FILLER_169_1157 ();
 FILLCELL_X32 FILLER_169_1189 ();
 FILLCELL_X32 FILLER_169_1221 ();
 FILLCELL_X8 FILLER_169_1253 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X16 FILLER_170_321 ();
 FILLCELL_X1 FILLER_170_337 ();
 FILLCELL_X8 FILLER_170_342 ();
 FILLCELL_X1 FILLER_170_350 ();
 FILLCELL_X1 FILLER_170_355 ();
 FILLCELL_X32 FILLER_170_366 ();
 FILLCELL_X4 FILLER_170_398 ();
 FILLCELL_X2 FILLER_170_402 ();
 FILLCELL_X1 FILLER_170_404 ();
 FILLCELL_X4 FILLER_170_413 ();
 FILLCELL_X32 FILLER_170_426 ();
 FILLCELL_X16 FILLER_170_458 ();
 FILLCELL_X1 FILLER_170_474 ();
 FILLCELL_X8 FILLER_170_495 ();
 FILLCELL_X4 FILLER_170_503 ();
 FILLCELL_X1 FILLER_170_507 ();
 FILLCELL_X4 FILLER_170_531 ();
 FILLCELL_X4 FILLER_170_540 ();
 FILLCELL_X2 FILLER_170_544 ();
 FILLCELL_X1 FILLER_170_546 ();
 FILLCELL_X4 FILLER_170_555 ();
 FILLCELL_X2 FILLER_170_559 ();
 FILLCELL_X1 FILLER_170_561 ();
 FILLCELL_X4 FILLER_170_566 ();
 FILLCELL_X1 FILLER_170_570 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X2 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_644 ();
 FILLCELL_X32 FILLER_170_676 ();
 FILLCELL_X32 FILLER_170_708 ();
 FILLCELL_X32 FILLER_170_740 ();
 FILLCELL_X32 FILLER_170_772 ();
 FILLCELL_X32 FILLER_170_804 ();
 FILLCELL_X32 FILLER_170_836 ();
 FILLCELL_X32 FILLER_170_868 ();
 FILLCELL_X32 FILLER_170_900 ();
 FILLCELL_X32 FILLER_170_932 ();
 FILLCELL_X32 FILLER_170_964 ();
 FILLCELL_X32 FILLER_170_996 ();
 FILLCELL_X32 FILLER_170_1028 ();
 FILLCELL_X32 FILLER_170_1060 ();
 FILLCELL_X32 FILLER_170_1092 ();
 FILLCELL_X32 FILLER_170_1124 ();
 FILLCELL_X32 FILLER_170_1156 ();
 FILLCELL_X32 FILLER_170_1188 ();
 FILLCELL_X32 FILLER_170_1220 ();
 FILLCELL_X32 FILLER_170_1252 ();
 FILLCELL_X32 FILLER_170_1284 ();
 FILLCELL_X8 FILLER_170_1316 ();
 FILLCELL_X4 FILLER_170_1324 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X8 FILLER_171_321 ();
 FILLCELL_X4 FILLER_171_329 ();
 FILLCELL_X32 FILLER_171_350 ();
 FILLCELL_X16 FILLER_171_382 ();
 FILLCELL_X2 FILLER_171_398 ();
 FILLCELL_X1 FILLER_171_400 ();
 FILLCELL_X8 FILLER_171_422 ();
 FILLCELL_X4 FILLER_171_430 ();
 FILLCELL_X2 FILLER_171_434 ();
 FILLCELL_X1 FILLER_171_436 ();
 FILLCELL_X32 FILLER_171_439 ();
 FILLCELL_X1 FILLER_171_471 ();
 FILLCELL_X16 FILLER_171_489 ();
 FILLCELL_X4 FILLER_171_505 ();
 FILLCELL_X2 FILLER_171_509 ();
 FILLCELL_X1 FILLER_171_511 ();
 FILLCELL_X4 FILLER_171_525 ();
 FILLCELL_X8 FILLER_171_546 ();
 FILLCELL_X4 FILLER_171_554 ();
 FILLCELL_X1 FILLER_171_558 ();
 FILLCELL_X1 FILLER_171_561 ();
 FILLCELL_X32 FILLER_171_566 ();
 FILLCELL_X16 FILLER_171_598 ();
 FILLCELL_X8 FILLER_171_614 ();
 FILLCELL_X1 FILLER_171_622 ();
 FILLCELL_X2 FILLER_171_655 ();
 FILLCELL_X32 FILLER_171_674 ();
 FILLCELL_X32 FILLER_171_706 ();
 FILLCELL_X32 FILLER_171_738 ();
 FILLCELL_X32 FILLER_171_770 ();
 FILLCELL_X32 FILLER_171_802 ();
 FILLCELL_X32 FILLER_171_834 ();
 FILLCELL_X32 FILLER_171_866 ();
 FILLCELL_X32 FILLER_171_898 ();
 FILLCELL_X32 FILLER_171_930 ();
 FILLCELL_X32 FILLER_171_962 ();
 FILLCELL_X32 FILLER_171_994 ();
 FILLCELL_X32 FILLER_171_1026 ();
 FILLCELL_X32 FILLER_171_1058 ();
 FILLCELL_X32 FILLER_171_1090 ();
 FILLCELL_X32 FILLER_171_1122 ();
 FILLCELL_X32 FILLER_171_1154 ();
 FILLCELL_X32 FILLER_171_1186 ();
 FILLCELL_X32 FILLER_171_1218 ();
 FILLCELL_X8 FILLER_171_1250 ();
 FILLCELL_X4 FILLER_171_1258 ();
 FILLCELL_X1 FILLER_171_1262 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X1 FILLER_172_353 ();
 FILLCELL_X1 FILLER_172_368 ();
 FILLCELL_X32 FILLER_172_391 ();
 FILLCELL_X32 FILLER_172_423 ();
 FILLCELL_X8 FILLER_172_455 ();
 FILLCELL_X2 FILLER_172_480 ();
 FILLCELL_X1 FILLER_172_482 ();
 FILLCELL_X32 FILLER_172_487 ();
 FILLCELL_X1 FILLER_172_519 ();
 FILLCELL_X32 FILLER_172_537 ();
 FILLCELL_X32 FILLER_172_569 ();
 FILLCELL_X1 FILLER_172_601 ();
 FILLCELL_X16 FILLER_172_606 ();
 FILLCELL_X8 FILLER_172_622 ();
 FILLCELL_X1 FILLER_172_630 ();
 FILLCELL_X2 FILLER_172_632 ();
 FILLCELL_X1 FILLER_172_634 ();
 FILLCELL_X32 FILLER_172_645 ();
 FILLCELL_X32 FILLER_172_677 ();
 FILLCELL_X32 FILLER_172_709 ();
 FILLCELL_X32 FILLER_172_741 ();
 FILLCELL_X32 FILLER_172_773 ();
 FILLCELL_X32 FILLER_172_805 ();
 FILLCELL_X32 FILLER_172_837 ();
 FILLCELL_X32 FILLER_172_869 ();
 FILLCELL_X32 FILLER_172_901 ();
 FILLCELL_X32 FILLER_172_933 ();
 FILLCELL_X32 FILLER_172_965 ();
 FILLCELL_X32 FILLER_172_997 ();
 FILLCELL_X32 FILLER_172_1029 ();
 FILLCELL_X32 FILLER_172_1061 ();
 FILLCELL_X32 FILLER_172_1093 ();
 FILLCELL_X32 FILLER_172_1125 ();
 FILLCELL_X32 FILLER_172_1157 ();
 FILLCELL_X32 FILLER_172_1189 ();
 FILLCELL_X32 FILLER_172_1221 ();
 FILLCELL_X32 FILLER_172_1253 ();
 FILLCELL_X32 FILLER_172_1285 ();
 FILLCELL_X8 FILLER_172_1317 ();
 FILLCELL_X2 FILLER_172_1325 ();
 FILLCELL_X1 FILLER_172_1327 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X16 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_383 ();
 FILLCELL_X16 FILLER_173_415 ();
 FILLCELL_X4 FILLER_173_431 ();
 FILLCELL_X2 FILLER_173_435 ();
 FILLCELL_X1 FILLER_173_437 ();
 FILLCELL_X16 FILLER_173_460 ();
 FILLCELL_X8 FILLER_173_476 ();
 FILLCELL_X16 FILLER_173_491 ();
 FILLCELL_X2 FILLER_173_507 ();
 FILLCELL_X32 FILLER_173_517 ();
 FILLCELL_X1 FILLER_173_549 ();
 FILLCELL_X4 FILLER_173_554 ();
 FILLCELL_X4 FILLER_173_566 ();
 FILLCELL_X2 FILLER_173_570 ();
 FILLCELL_X1 FILLER_173_572 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X16 FILLER_173_609 ();
 FILLCELL_X4 FILLER_173_625 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X32 FILLER_173_1089 ();
 FILLCELL_X32 FILLER_173_1121 ();
 FILLCELL_X32 FILLER_173_1153 ();
 FILLCELL_X32 FILLER_173_1185 ();
 FILLCELL_X32 FILLER_173_1217 ();
 FILLCELL_X8 FILLER_173_1249 ();
 FILLCELL_X4 FILLER_173_1257 ();
 FILLCELL_X2 FILLER_173_1261 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X16 FILLER_174_353 ();
 FILLCELL_X8 FILLER_174_369 ();
 FILLCELL_X8 FILLER_174_384 ();
 FILLCELL_X4 FILLER_174_392 ();
 FILLCELL_X1 FILLER_174_396 ();
 FILLCELL_X2 FILLER_174_400 ();
 FILLCELL_X4 FILLER_174_404 ();
 FILLCELL_X16 FILLER_174_415 ();
 FILLCELL_X2 FILLER_174_431 ();
 FILLCELL_X1 FILLER_174_433 ();
 FILLCELL_X1 FILLER_174_448 ();
 FILLCELL_X2 FILLER_174_460 ();
 FILLCELL_X8 FILLER_174_472 ();
 FILLCELL_X2 FILLER_174_480 ();
 FILLCELL_X1 FILLER_174_482 ();
 FILLCELL_X8 FILLER_174_492 ();
 FILLCELL_X1 FILLER_174_500 ();
 FILLCELL_X32 FILLER_174_516 ();
 FILLCELL_X8 FILLER_174_548 ();
 FILLCELL_X2 FILLER_174_556 ();
 FILLCELL_X1 FILLER_174_558 ();
 FILLCELL_X4 FILLER_174_576 ();
 FILLCELL_X32 FILLER_174_597 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X16 FILLER_174_1304 ();
 FILLCELL_X8 FILLER_174_1320 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X4 FILLER_175_385 ();
 FILLCELL_X2 FILLER_175_389 ();
 FILLCELL_X1 FILLER_175_391 ();
 FILLCELL_X2 FILLER_175_414 ();
 FILLCELL_X1 FILLER_175_416 ();
 FILLCELL_X2 FILLER_175_434 ();
 FILLCELL_X32 FILLER_175_447 ();
 FILLCELL_X16 FILLER_175_479 ();
 FILLCELL_X8 FILLER_175_495 ();
 FILLCELL_X4 FILLER_175_503 ();
 FILLCELL_X32 FILLER_175_521 ();
 FILLCELL_X32 FILLER_175_553 ();
 FILLCELL_X1 FILLER_175_585 ();
 FILLCELL_X16 FILLER_175_596 ();
 FILLCELL_X8 FILLER_175_612 ();
 FILLCELL_X4 FILLER_175_620 ();
 FILLCELL_X2 FILLER_175_624 ();
 FILLCELL_X32 FILLER_175_643 ();
 FILLCELL_X32 FILLER_175_675 ();
 FILLCELL_X32 FILLER_175_707 ();
 FILLCELL_X32 FILLER_175_739 ();
 FILLCELL_X32 FILLER_175_771 ();
 FILLCELL_X32 FILLER_175_803 ();
 FILLCELL_X32 FILLER_175_835 ();
 FILLCELL_X32 FILLER_175_867 ();
 FILLCELL_X32 FILLER_175_899 ();
 FILLCELL_X32 FILLER_175_931 ();
 FILLCELL_X32 FILLER_175_963 ();
 FILLCELL_X32 FILLER_175_995 ();
 FILLCELL_X32 FILLER_175_1027 ();
 FILLCELL_X32 FILLER_175_1059 ();
 FILLCELL_X32 FILLER_175_1091 ();
 FILLCELL_X32 FILLER_175_1123 ();
 FILLCELL_X32 FILLER_175_1155 ();
 FILLCELL_X32 FILLER_175_1187 ();
 FILLCELL_X32 FILLER_175_1219 ();
 FILLCELL_X8 FILLER_175_1251 ();
 FILLCELL_X4 FILLER_175_1259 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X8 FILLER_176_353 ();
 FILLCELL_X4 FILLER_176_361 ();
 FILLCELL_X4 FILLER_176_385 ();
 FILLCELL_X8 FILLER_176_401 ();
 FILLCELL_X4 FILLER_176_409 ();
 FILLCELL_X2 FILLER_176_413 ();
 FILLCELL_X2 FILLER_176_424 ();
 FILLCELL_X2 FILLER_176_433 ();
 FILLCELL_X16 FILLER_176_445 ();
 FILLCELL_X4 FILLER_176_461 ();
 FILLCELL_X2 FILLER_176_465 ();
 FILLCELL_X1 FILLER_176_467 ();
 FILLCELL_X2 FILLER_176_478 ();
 FILLCELL_X1 FILLER_176_480 ();
 FILLCELL_X16 FILLER_176_491 ();
 FILLCELL_X1 FILLER_176_507 ();
 FILLCELL_X1 FILLER_176_517 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X4 FILLER_176_577 ();
 FILLCELL_X2 FILLER_176_581 ();
 FILLCELL_X1 FILLER_176_583 ();
 FILLCELL_X1 FILLER_176_588 ();
 FILLCELL_X16 FILLER_176_602 ();
 FILLCELL_X8 FILLER_176_618 ();
 FILLCELL_X4 FILLER_176_626 ();
 FILLCELL_X1 FILLER_176_630 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X32 FILLER_176_1112 ();
 FILLCELL_X32 FILLER_176_1144 ();
 FILLCELL_X32 FILLER_176_1176 ();
 FILLCELL_X32 FILLER_176_1208 ();
 FILLCELL_X32 FILLER_176_1240 ();
 FILLCELL_X32 FILLER_176_1272 ();
 FILLCELL_X16 FILLER_176_1304 ();
 FILLCELL_X8 FILLER_176_1320 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X16 FILLER_177_353 ();
 FILLCELL_X4 FILLER_177_369 ();
 FILLCELL_X2 FILLER_177_373 ();
 FILLCELL_X1 FILLER_177_393 ();
 FILLCELL_X8 FILLER_177_401 ();
 FILLCELL_X1 FILLER_177_409 ();
 FILLCELL_X4 FILLER_177_424 ();
 FILLCELL_X1 FILLER_177_428 ();
 FILLCELL_X16 FILLER_177_439 ();
 FILLCELL_X8 FILLER_177_455 ();
 FILLCELL_X4 FILLER_177_463 ();
 FILLCELL_X2 FILLER_177_467 ();
 FILLCELL_X1 FILLER_177_469 ();
 FILLCELL_X1 FILLER_177_480 ();
 FILLCELL_X8 FILLER_177_504 ();
 FILLCELL_X4 FILLER_177_512 ();
 FILLCELL_X1 FILLER_177_525 ();
 FILLCELL_X4 FILLER_177_540 ();
 FILLCELL_X2 FILLER_177_544 ();
 FILLCELL_X32 FILLER_177_550 ();
 FILLCELL_X1 FILLER_177_595 ();
 FILLCELL_X4 FILLER_177_644 ();
 FILLCELL_X32 FILLER_177_665 ();
 FILLCELL_X32 FILLER_177_697 ();
 FILLCELL_X32 FILLER_177_729 ();
 FILLCELL_X32 FILLER_177_761 ();
 FILLCELL_X32 FILLER_177_793 ();
 FILLCELL_X32 FILLER_177_825 ();
 FILLCELL_X32 FILLER_177_857 ();
 FILLCELL_X32 FILLER_177_889 ();
 FILLCELL_X32 FILLER_177_921 ();
 FILLCELL_X32 FILLER_177_953 ();
 FILLCELL_X32 FILLER_177_985 ();
 FILLCELL_X32 FILLER_177_1017 ();
 FILLCELL_X32 FILLER_177_1049 ();
 FILLCELL_X32 FILLER_177_1081 ();
 FILLCELL_X32 FILLER_177_1113 ();
 FILLCELL_X32 FILLER_177_1145 ();
 FILLCELL_X32 FILLER_177_1177 ();
 FILLCELL_X32 FILLER_177_1209 ();
 FILLCELL_X16 FILLER_177_1241 ();
 FILLCELL_X4 FILLER_177_1257 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X1 FILLER_178_385 ();
 FILLCELL_X16 FILLER_178_396 ();
 FILLCELL_X4 FILLER_178_412 ();
 FILLCELL_X2 FILLER_178_416 ();
 FILLCELL_X32 FILLER_178_432 ();
 FILLCELL_X4 FILLER_178_464 ();
 FILLCELL_X2 FILLER_178_474 ();
 FILLCELL_X4 FILLER_178_480 ();
 FILLCELL_X2 FILLER_178_484 ();
 FILLCELL_X16 FILLER_178_493 ();
 FILLCELL_X4 FILLER_178_509 ();
 FILLCELL_X2 FILLER_178_513 ();
 FILLCELL_X1 FILLER_178_515 ();
 FILLCELL_X1 FILLER_178_519 ();
 FILLCELL_X8 FILLER_178_534 ();
 FILLCELL_X2 FILLER_178_542 ();
 FILLCELL_X1 FILLER_178_544 ();
 FILLCELL_X32 FILLER_178_562 ();
 FILLCELL_X4 FILLER_178_607 ();
 FILLCELL_X2 FILLER_178_611 ();
 FILLCELL_X1 FILLER_178_613 ();
 FILLCELL_X16 FILLER_178_632 ();
 FILLCELL_X8 FILLER_178_648 ();
 FILLCELL_X4 FILLER_178_656 ();
 FILLCELL_X32 FILLER_178_663 ();
 FILLCELL_X32 FILLER_178_695 ();
 FILLCELL_X32 FILLER_178_727 ();
 FILLCELL_X32 FILLER_178_759 ();
 FILLCELL_X32 FILLER_178_791 ();
 FILLCELL_X32 FILLER_178_823 ();
 FILLCELL_X32 FILLER_178_855 ();
 FILLCELL_X32 FILLER_178_887 ();
 FILLCELL_X32 FILLER_178_919 ();
 FILLCELL_X32 FILLER_178_951 ();
 FILLCELL_X32 FILLER_178_983 ();
 FILLCELL_X32 FILLER_178_1015 ();
 FILLCELL_X32 FILLER_178_1047 ();
 FILLCELL_X32 FILLER_178_1079 ();
 FILLCELL_X32 FILLER_178_1111 ();
 FILLCELL_X32 FILLER_178_1143 ();
 FILLCELL_X32 FILLER_178_1175 ();
 FILLCELL_X32 FILLER_178_1207 ();
 FILLCELL_X32 FILLER_178_1239 ();
 FILLCELL_X32 FILLER_178_1271 ();
 FILLCELL_X16 FILLER_178_1303 ();
 FILLCELL_X8 FILLER_178_1319 ();
 FILLCELL_X1 FILLER_178_1327 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X8 FILLER_179_353 ();
 FILLCELL_X2 FILLER_179_361 ();
 FILLCELL_X2 FILLER_179_366 ();
 FILLCELL_X1 FILLER_179_368 ();
 FILLCELL_X8 FILLER_179_375 ();
 FILLCELL_X16 FILLER_179_395 ();
 FILLCELL_X4 FILLER_179_411 ();
 FILLCELL_X2 FILLER_179_415 ();
 FILLCELL_X2 FILLER_179_420 ();
 FILLCELL_X1 FILLER_179_422 ();
 FILLCELL_X4 FILLER_179_429 ();
 FILLCELL_X2 FILLER_179_433 ();
 FILLCELL_X8 FILLER_179_441 ();
 FILLCELL_X1 FILLER_179_449 ();
 FILLCELL_X8 FILLER_179_459 ();
 FILLCELL_X2 FILLER_179_467 ();
 FILLCELL_X2 FILLER_179_481 ();
 FILLCELL_X8 FILLER_179_491 ();
 FILLCELL_X1 FILLER_179_499 ();
 FILLCELL_X16 FILLER_179_503 ();
 FILLCELL_X2 FILLER_179_525 ();
 FILLCELL_X4 FILLER_179_533 ();
 FILLCELL_X2 FILLER_179_537 ();
 FILLCELL_X1 FILLER_179_539 ();
 FILLCELL_X1 FILLER_179_550 ();
 FILLCELL_X2 FILLER_179_563 ();
 FILLCELL_X1 FILLER_179_565 ();
 FILLCELL_X8 FILLER_179_570 ();
 FILLCELL_X1 FILLER_179_578 ();
 FILLCELL_X2 FILLER_179_582 ();
 FILLCELL_X1 FILLER_179_584 ();
 FILLCELL_X2 FILLER_179_597 ();
 FILLCELL_X4 FILLER_179_602 ();
 FILLCELL_X1 FILLER_179_606 ();
 FILLCELL_X8 FILLER_179_616 ();
 FILLCELL_X2 FILLER_179_632 ();
 FILLCELL_X1 FILLER_179_640 ();
 FILLCELL_X4 FILLER_179_644 ();
 FILLCELL_X2 FILLER_179_648 ();
 FILLCELL_X4 FILLER_179_661 ();
 FILLCELL_X2 FILLER_179_665 ();
 FILLCELL_X2 FILLER_179_670 ();
 FILLCELL_X8 FILLER_179_675 ();
 FILLCELL_X32 FILLER_179_688 ();
 FILLCELL_X32 FILLER_179_720 ();
 FILLCELL_X32 FILLER_179_752 ();
 FILLCELL_X16 FILLER_179_784 ();
 FILLCELL_X8 FILLER_179_800 ();
 FILLCELL_X32 FILLER_179_816 ();
 FILLCELL_X32 FILLER_179_848 ();
 FILLCELL_X32 FILLER_179_880 ();
 FILLCELL_X32 FILLER_179_912 ();
 FILLCELL_X32 FILLER_179_944 ();
 FILLCELL_X32 FILLER_179_981 ();
 FILLCELL_X2 FILLER_179_1013 ();
 FILLCELL_X1 FILLER_179_1015 ();
 FILLCELL_X1 FILLER_179_1018 ();
 FILLCELL_X8 FILLER_179_1027 ();
 FILLCELL_X1 FILLER_179_1040 ();
 FILLCELL_X1 FILLER_179_1054 ();
 FILLCELL_X8 FILLER_179_1057 ();
 FILLCELL_X2 FILLER_179_1065 ();
 FILLCELL_X4 FILLER_179_1072 ();
 FILLCELL_X2 FILLER_179_1076 ();
 FILLCELL_X1 FILLER_179_1078 ();
 FILLCELL_X1 FILLER_179_1092 ();
 FILLCELL_X16 FILLER_179_1095 ();
 FILLCELL_X4 FILLER_179_1111 ();
 FILLCELL_X2 FILLER_179_1115 ();
 FILLCELL_X32 FILLER_179_1122 ();
 FILLCELL_X32 FILLER_179_1154 ();
 FILLCELL_X32 FILLER_179_1186 ();
 FILLCELL_X32 FILLER_179_1218 ();
 FILLCELL_X8 FILLER_179_1250 ();
 FILLCELL_X4 FILLER_179_1258 ();
 FILLCELL_X32 FILLER_179_1263 ();
 FILLCELL_X32 FILLER_179_1295 ();
 FILLCELL_X1 FILLER_179_1327 ();
endmodule
