module bist_controller (bist_done,
    bist_pass,
    bist_start,
    clk,
    mem_enable,
    mem_write,
    rst_n,
    error_addr,
    error_count,
    mem_addr,
    mem_rdata,
    mem_wdata);
 output bist_done;
 output bist_pass;
 input bist_start;
 input clk;
 output mem_enable;
 output mem_write;
 input rst_n;
 output [4:0] error_addr;
 output [31:0] error_count;
 output [4:0] mem_addr;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire phase_complete;
 wire read_phase;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 BUF_X2 _0538_ (.A(net74),
    .Z(_0054_));
 NAND3_X2 _0539_ (.A1(net75),
    .A2(_0054_),
    .A3(_0529_),
    .ZN(_0532_));
 INV_X1 _0540_ (.A(_0532_),
    .ZN(_0535_));
 BUF_X4 _0541_ (.A(rst_n),
    .Z(_0055_));
 INV_X1 _0542_ (.A(_0055_),
    .ZN(_0056_));
 CLKBUF_X3 _0543_ (.A(_0056_),
    .Z(_0057_));
 CLKBUF_X3 _0544_ (.A(_0057_),
    .Z(_0058_));
 BUF_X1 _0545_ (.A(net72),
    .Z(_0059_));
 CLKBUF_X3 _0546_ (.A(\state[0] ),
    .Z(_0060_));
 BUF_X4 _0547_ (.A(_0060_),
    .Z(_0061_));
 CLKBUF_X2 _0548_ (.A(\state[3] ),
    .Z(_0062_));
 INV_X2 _0549_ (.A(_0062_),
    .ZN(_0063_));
 NAND2_X1 _0550_ (.A1(_0061_),
    .A2(_0063_),
    .ZN(_0064_));
 BUF_X4 _0551_ (.A(\state[2] ),
    .Z(_0065_));
 CLKBUF_X2 _0552_ (.A(_0001_),
    .Z(_0066_));
 NAND2_X1 _0553_ (.A1(_0065_),
    .A2(_0066_),
    .ZN(_0067_));
 CLKBUF_X3 _0554_ (.A(\state[1] ),
    .Z(_0068_));
 BUF_X4 _0555_ (.A(_0068_),
    .Z(_0069_));
 CLKBUF_X2 _0556_ (.A(_0000_),
    .Z(_0070_));
 INV_X1 _0557_ (.A(_0070_),
    .ZN(_0071_));
 BUF_X4 _0558_ (.A(_0062_),
    .Z(_0072_));
 CLKBUF_X3 _0559_ (.A(_0072_),
    .Z(_0073_));
 INV_X2 _0560_ (.A(_0065_),
    .ZN(_0074_));
 BUF_X2 _0561_ (.A(phase_complete),
    .Z(_0075_));
 CLKBUF_X3 _0562_ (.A(read_phase),
    .Z(_0076_));
 OR2_X1 _0563_ (.A1(_0075_),
    .A2(_0076_),
    .ZN(_0077_));
 NOR3_X1 _0564_ (.A1(_0073_),
    .A2(_0074_),
    .A3(_0077_),
    .ZN(_0078_));
 OAI21_X1 _0565_ (.A(_0069_),
    .B1(_0071_),
    .B2(_0078_),
    .ZN(_0079_));
 AOI21_X2 _0566_ (.A(_0064_),
    .B1(_0067_),
    .B2(_0079_),
    .ZN(_0080_));
 CLKBUF_X2 _0567_ (.A(bist_start),
    .Z(_0081_));
 NOR4_X2 _0568_ (.A1(_0061_),
    .A2(_0069_),
    .A3(_0065_),
    .A4(_0081_),
    .ZN(_0082_));
 NOR2_X2 _0569_ (.A1(_0072_),
    .A2(_0082_),
    .ZN(_0083_));
 INV_X2 _0570_ (.A(_0068_),
    .ZN(_0084_));
 NOR2_X1 _0571_ (.A1(_0084_),
    .A2(_0072_),
    .ZN(_0085_));
 BUF_X4 _0572_ (.A(_0065_),
    .Z(_0086_));
 OAI21_X1 _0573_ (.A(_0067_),
    .B1(_0075_),
    .B2(_0086_),
    .ZN(_0087_));
 NOR2_X4 _0574_ (.A1(_0060_),
    .A2(_0068_),
    .ZN(_0088_));
 AND3_X2 _0575_ (.A1(_0063_),
    .A2(_0065_),
    .A3(_0088_),
    .ZN(_0089_));
 CLKBUF_X2 _0576_ (.A(net110),
    .Z(_0090_));
 INV_X1 _0577_ (.A(_0090_),
    .ZN(_0091_));
 AOI21_X1 _0578_ (.A(_0077_),
    .B1(_0066_),
    .B2(_0091_),
    .ZN(_0092_));
 AOI22_X2 _0579_ (.A1(_0085_),
    .A2(_0087_),
    .B1(_0089_),
    .B2(_0092_),
    .ZN(_0093_));
 AOI21_X2 _0580_ (.A(_0065_),
    .B1(_0069_),
    .B2(_0061_),
    .ZN(_0094_));
 NOR2_X2 _0581_ (.A1(_0072_),
    .A2(_0094_),
    .ZN(_0095_));
 AOI21_X1 _0582_ (.A(_0065_),
    .B1(_0076_),
    .B2(_0091_),
    .ZN(_0096_));
 NAND2_X2 _0583_ (.A1(_0061_),
    .A2(_0069_),
    .ZN(_0097_));
 INV_X1 _0584_ (.A(_0066_),
    .ZN(_0098_));
 NAND2_X1 _0585_ (.A1(_0091_),
    .A2(_0098_),
    .ZN(_0099_));
 OAI221_X2 _0586_ (.A(_0095_),
    .B1(_0096_),
    .B2(_0097_),
    .C1(_0076_),
    .C2(_0099_),
    .ZN(_0100_));
 NAND3_X1 _0587_ (.A1(_0083_),
    .A2(_0093_),
    .A3(_0100_),
    .ZN(_0101_));
 OAI21_X1 _0588_ (.A(_0059_),
    .B1(_0080_),
    .B2(_0101_),
    .ZN(_0102_));
 INV_X1 _0589_ (.A(_0064_),
    .ZN(_0103_));
 NOR2_X1 _0590_ (.A1(_0074_),
    .A2(_0098_),
    .ZN(_0104_));
 OR3_X1 _0591_ (.A1(_0072_),
    .A2(_0074_),
    .A3(_0077_),
    .ZN(_0105_));
 AOI21_X1 _0592_ (.A(_0084_),
    .B1(_0070_),
    .B2(_0105_),
    .ZN(_0106_));
 OAI21_X2 _0593_ (.A(_0103_),
    .B1(_0104_),
    .B2(_0106_),
    .ZN(_0107_));
 AND3_X2 _0594_ (.A1(_0083_),
    .A2(_0093_),
    .A3(_0100_),
    .ZN(_0108_));
 NOR2_X1 _0595_ (.A1(_0069_),
    .A2(_0086_),
    .ZN(_0109_));
 OR2_X1 _0596_ (.A1(_0073_),
    .A2(_0109_),
    .ZN(_0110_));
 NOR3_X2 _0597_ (.A1(_0072_),
    .A2(_0074_),
    .A3(_0088_),
    .ZN(_0111_));
 INV_X1 _0598_ (.A(_0527_),
    .ZN(_0112_));
 OR3_X2 _0599_ (.A1(net75),
    .A2(_0054_),
    .A3(_0112_),
    .ZN(_0113_));
 INV_X1 _0600_ (.A(_0531_),
    .ZN(_0114_));
 OAI21_X4 _0601_ (.A(_0111_),
    .B1(_0113_),
    .B2(_0114_),
    .ZN(_0115_));
 NOR3_X4 _0602_ (.A1(_0084_),
    .A2(_0072_),
    .A3(_0086_),
    .ZN(_0116_));
 INV_X1 _0603_ (.A(_0536_),
    .ZN(_0117_));
 AOI21_X2 _0604_ (.A(_0089_),
    .B1(_0116_),
    .B2(_0117_),
    .ZN(_0118_));
 NAND2_X1 _0605_ (.A1(_0536_),
    .A2(_0088_),
    .ZN(_0119_));
 AOI221_X1 _0606_ (.A(_0110_),
    .B1(_0115_),
    .B2(_0118_),
    .C1(_0119_),
    .C2(_0059_),
    .ZN(_0120_));
 NAND3_X1 _0607_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0120_),
    .ZN(_0121_));
 AOI21_X1 _0608_ (.A(_0058_),
    .B1(_0102_),
    .B2(_0121_),
    .ZN(_0003_));
 AOI21_X1 _0609_ (.A(net73),
    .B1(_0107_),
    .B2(_0108_),
    .ZN(_0122_));
 NAND2_X1 _0610_ (.A1(_0536_),
    .A2(_0089_),
    .ZN(_0123_));
 MUX2_X1 _0611_ (.A(_0115_),
    .B(_0118_),
    .S(_0528_),
    .Z(_0124_));
 AND4_X1 _0612_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0123_),
    .A4(_0124_),
    .ZN(_0125_));
 NOR3_X1 _0613_ (.A1(_0058_),
    .A2(_0122_),
    .A3(_0125_),
    .ZN(_0004_));
 OAI221_X1 _0614_ (.A(_0054_),
    .B1(_0527_),
    .B2(_0115_),
    .C1(_0118_),
    .C2(_0529_),
    .ZN(_0126_));
 INV_X1 _0615_ (.A(_0529_),
    .ZN(_0127_));
 OAI22_X1 _0616_ (.A1(_0112_),
    .A2(_0115_),
    .B1(_0118_),
    .B2(_0127_),
    .ZN(_0128_));
 OAI21_X1 _0617_ (.A(_0126_),
    .B1(_0128_),
    .B2(_0054_),
    .ZN(_0129_));
 AND3_X1 _0618_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0123_),
    .ZN(_0130_));
 NAND2_X1 _0619_ (.A1(_0107_),
    .A2(_0108_),
    .ZN(_0131_));
 INV_X1 _0620_ (.A(_0054_),
    .ZN(_0132_));
 AOI221_X1 _0621_ (.A(_0057_),
    .B1(_0129_),
    .B2(_0130_),
    .C1(_0131_),
    .C2(_0132_),
    .ZN(_0005_));
 AOI21_X1 _0622_ (.A(net75),
    .B1(_0107_),
    .B2(_0108_),
    .ZN(_0133_));
 NOR3_X1 _0623_ (.A1(_0054_),
    .A2(_0059_),
    .A3(net73),
    .ZN(_0134_));
 XOR2_X1 _0624_ (.A(_0002_),
    .B(_0134_),
    .Z(_0135_));
 NAND3_X1 _0625_ (.A1(_0054_),
    .A2(_0059_),
    .A3(net73),
    .ZN(_0136_));
 XOR2_X1 _0626_ (.A(_0002_),
    .B(_0136_),
    .Z(_0137_));
 NOR2_X1 _0627_ (.A1(_0536_),
    .A2(_0137_),
    .ZN(_0138_));
 OAI22_X1 _0628_ (.A1(_0115_),
    .A2(_0135_),
    .B1(_0138_),
    .B2(_0118_),
    .ZN(_0139_));
 NOR3_X1 _0629_ (.A1(_0080_),
    .A2(_0101_),
    .A3(_0139_),
    .ZN(_0140_));
 NOR3_X1 _0630_ (.A1(_0058_),
    .A2(_0133_),
    .A3(_0140_),
    .ZN(_0006_));
 AOI21_X1 _0631_ (.A(net76),
    .B1(_0107_),
    .B2(_0108_),
    .ZN(_0141_));
 NAND2_X1 _0632_ (.A1(_0534_),
    .A2(_0116_),
    .ZN(_0142_));
 INV_X1 _0633_ (.A(_0533_),
    .ZN(_0143_));
 NOR2_X1 _0634_ (.A1(_0531_),
    .A2(_0088_),
    .ZN(_0144_));
 AOI22_X1 _0635_ (.A1(_0143_),
    .A2(_0088_),
    .B1(_0113_),
    .B2(_0144_),
    .ZN(_0145_));
 NAND2_X1 _0636_ (.A1(_0063_),
    .A2(_0086_),
    .ZN(_0146_));
 OAI21_X1 _0637_ (.A(_0142_),
    .B1(_0145_),
    .B2(_0146_),
    .ZN(_0147_));
 NOR3_X1 _0638_ (.A1(_0080_),
    .A2(_0101_),
    .A3(_0147_),
    .ZN(_0148_));
 NOR3_X1 _0639_ (.A1(_0058_),
    .A2(_0141_),
    .A3(_0148_),
    .ZN(_0007_));
 NOR3_X2 _0640_ (.A1(_0061_),
    .A2(_0069_),
    .A3(_0065_),
    .ZN(_0149_));
 NAND2_X1 _0641_ (.A1(_0073_),
    .A2(_0149_),
    .ZN(_0150_));
 NAND2_X1 _0642_ (.A1(_0081_),
    .A2(_0149_),
    .ZN(_0151_));
 NAND2_X1 _0643_ (.A1(net33),
    .A2(_0151_),
    .ZN(_0152_));
 AOI21_X1 _0644_ (.A(_0058_),
    .B1(_0150_),
    .B2(_0152_),
    .ZN(_0008_));
 INV_X1 _0645_ (.A(_0521_),
    .ZN(_0153_));
 NOR4_X1 _0646_ (.A1(net58),
    .A2(net63),
    .A3(net64),
    .A4(_0153_),
    .ZN(_0154_));
 BUF_X1 _0647_ (.A(net60),
    .Z(_0155_));
 NOR4_X1 _0648_ (.A1(net49),
    .A2(net59),
    .A3(_0155_),
    .A4(net61),
    .ZN(_0156_));
 BUF_X1 _0649_ (.A(net56),
    .Z(_0157_));
 BUF_X1 _0650_ (.A(net57),
    .Z(_0158_));
 NOR4_X1 _0651_ (.A1(net54),
    .A2(net55),
    .A3(_0157_),
    .A4(_0158_),
    .ZN(_0159_));
 BUF_X1 _0652_ (.A(net50),
    .Z(_0160_));
 BUF_X1 _0653_ (.A(net53),
    .Z(_0161_));
 NOR3_X1 _0654_ (.A1(_0160_),
    .A2(net52),
    .A3(_0161_),
    .ZN(_0162_));
 NAND4_X1 _0655_ (.A1(_0154_),
    .A2(_0156_),
    .A3(_0159_),
    .A4(_0162_),
    .ZN(_0163_));
 BUF_X2 _0656_ (.A(net68),
    .Z(_0164_));
 BUF_X4 _0657_ (.A(net69),
    .Z(_0165_));
 BUF_X1 _0658_ (.A(net70),
    .Z(_0166_));
 CLKBUF_X2 _0659_ (.A(net71),
    .Z(_0167_));
 NOR4_X1 _0660_ (.A1(_0164_),
    .A2(_0165_),
    .A3(_0166_),
    .A4(_0167_),
    .ZN(_0168_));
 CLKBUF_X2 _0661_ (.A(net62),
    .Z(_0169_));
 CLKBUF_X2 _0662_ (.A(net65),
    .Z(_0170_));
 CLKBUF_X2 _0663_ (.A(net66),
    .Z(_0171_));
 CLKBUF_X2 _0664_ (.A(net67),
    .Z(_0172_));
 NOR4_X1 _0665_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0171_),
    .A4(_0172_),
    .ZN(_0173_));
 BUF_X4 _0666_ (.A(net41),
    .Z(_0174_));
 NOR4_X1 _0667_ (.A1(_0174_),
    .A2(net45),
    .A3(net46),
    .A4(net47),
    .ZN(_0175_));
 BUF_X1 _0668_ (.A(net43),
    .Z(_0176_));
 CLKBUF_X2 _0669_ (.A(net48),
    .Z(_0177_));
 NOR4_X1 _0670_ (.A1(net42),
    .A2(_0176_),
    .A3(net44),
    .A4(_0177_),
    .ZN(_0178_));
 NAND4_X1 _0671_ (.A1(_0168_),
    .A2(_0173_),
    .A3(_0175_),
    .A4(_0178_),
    .ZN(_0179_));
 NOR3_X1 _0672_ (.A1(_0150_),
    .A2(_0163_),
    .A3(_0179_),
    .ZN(_0180_));
 OAI21_X1 _0673_ (.A(_0149_),
    .B1(_0081_),
    .B2(_0073_),
    .ZN(_0181_));
 AOI21_X1 _0674_ (.A(_0180_),
    .B1(_0181_),
    .B2(net34),
    .ZN(_0182_));
 NOR2_X1 _0675_ (.A1(_0058_),
    .A2(_0182_),
    .ZN(_0009_));
 BUF_X2 _0676_ (.A(_0055_),
    .Z(_0183_));
 AND2_X1 _0677_ (.A1(net35),
    .A2(_0183_),
    .ZN(_0184_));
 AND2_X1 _0678_ (.A1(_0059_),
    .A2(_0183_),
    .ZN(_0185_));
 OR2_X2 _0679_ (.A1(_0072_),
    .A2(_0094_),
    .ZN(_0186_));
 NAND3_X2 _0680_ (.A1(_0060_),
    .A2(_0068_),
    .A3(\state[2] ),
    .ZN(_0187_));
 NOR4_X2 _0681_ (.A1(_0072_),
    .A2(_0075_),
    .A3(_0076_),
    .A4(_0187_),
    .ZN(_0188_));
 AND2_X1 _0682_ (.A1(_0060_),
    .A2(_0068_),
    .ZN(_0189_));
 XNOR2_X1 _0683_ (.A(_0074_),
    .B(_0189_),
    .ZN(_0190_));
 NOR4_X2 _0684_ (.A1(_0072_),
    .A2(_0076_),
    .A3(_0090_),
    .A4(_0098_),
    .ZN(_0191_));
 AOI21_X2 _0685_ (.A(_0188_),
    .B1(_0190_),
    .B2(_0191_),
    .ZN(_0192_));
 NAND4_X1 _0686_ (.A1(net9),
    .A2(net13),
    .A3(net16),
    .A4(net15),
    .ZN(_0193_));
 NAND4_X1 _0687_ (.A1(net8),
    .A2(net11),
    .A3(net10),
    .A4(net14),
    .ZN(_0194_));
 NAND4_X1 _0688_ (.A1(net18),
    .A2(net21),
    .A3(net25),
    .A4(net24),
    .ZN(_0195_));
 NAND4_X1 _0689_ (.A1(net17),
    .A2(net20),
    .A3(net19),
    .A4(net22),
    .ZN(_0196_));
 NOR4_X1 _0690_ (.A1(_0193_),
    .A2(_0194_),
    .A3(_0195_),
    .A4(_0196_),
    .ZN(_0197_));
 NAND4_X1 _0691_ (.A1(net28),
    .A2(net27),
    .A3(net30),
    .A4(net6),
    .ZN(_0198_));
 NAND4_X1 _0692_ (.A1(net12),
    .A2(net1),
    .A3(net26),
    .A4(net23),
    .ZN(_0199_));
 NAND4_X1 _0693_ (.A1(net29),
    .A2(net5),
    .A3(net4),
    .A4(net7),
    .ZN(_0200_));
 NAND4_X1 _0694_ (.A1(net32),
    .A2(net31),
    .A3(net3),
    .A4(net2),
    .ZN(_0201_));
 NOR4_X1 _0695_ (.A1(_0198_),
    .A2(_0199_),
    .A3(_0200_),
    .A4(_0201_),
    .ZN(_0202_));
 AOI21_X1 _0696_ (.A(_0070_),
    .B1(_0197_),
    .B2(_0202_),
    .ZN(_0203_));
 NOR3_X1 _0697_ (.A1(_0076_),
    .A2(_0090_),
    .A3(_0098_),
    .ZN(_0204_));
 NOR2_X2 _0698_ (.A1(_0060_),
    .A2(_0062_),
    .ZN(_0205_));
 NAND2_X1 _0699_ (.A1(_0065_),
    .A2(_0205_),
    .ZN(_0206_));
 OR2_X1 _0700_ (.A1(_0204_),
    .A2(_0206_),
    .ZN(_0207_));
 OAI21_X2 _0701_ (.A(_0192_),
    .B1(_0203_),
    .B2(_0207_),
    .ZN(_0208_));
 INV_X1 _0702_ (.A(_0076_),
    .ZN(_0209_));
 NOR4_X1 _0703_ (.A1(net18),
    .A2(net17),
    .A3(net20),
    .A4(net24),
    .ZN(_0210_));
 NOR4_X1 _0704_ (.A1(net19),
    .A2(net22),
    .A3(net21),
    .A4(net25),
    .ZN(_0211_));
 NAND2_X1 _0705_ (.A1(_0210_),
    .A2(_0211_),
    .ZN(_0212_));
 NOR4_X1 _0706_ (.A1(net9),
    .A2(net8),
    .A3(net11),
    .A4(net15),
    .ZN(_0213_));
 NOR4_X1 _0707_ (.A1(net10),
    .A2(net14),
    .A3(net13),
    .A4(net16),
    .ZN(_0214_));
 NAND2_X1 _0708_ (.A1(_0213_),
    .A2(_0214_),
    .ZN(_0215_));
 NOR4_X1 _0709_ (.A1(net28),
    .A2(net27),
    .A3(net30),
    .A4(net6),
    .ZN(_0216_));
 NOR4_X1 _0710_ (.A1(net12),
    .A2(net1),
    .A3(net26),
    .A4(net23),
    .ZN(_0217_));
 NAND2_X1 _0711_ (.A1(_0216_),
    .A2(_0217_),
    .ZN(_0218_));
 NOR4_X1 _0712_ (.A1(net29),
    .A2(net5),
    .A3(net4),
    .A4(net7),
    .ZN(_0219_));
 NOR4_X1 _0713_ (.A1(net32),
    .A2(net31),
    .A3(net3),
    .A4(net2),
    .ZN(_0220_));
 NAND2_X1 _0714_ (.A1(_0219_),
    .A2(_0220_),
    .ZN(_0221_));
 OR4_X1 _0715_ (.A1(_0212_),
    .A2(_0215_),
    .A3(_0218_),
    .A4(_0221_),
    .ZN(_0222_));
 OAI21_X1 _0716_ (.A(_0071_),
    .B1(_0209_),
    .B2(_0222_),
    .ZN(_0223_));
 AOI211_X2 _0717_ (.A(_0186_),
    .B(_0208_),
    .C1(_0223_),
    .C2(_0206_),
    .ZN(_0224_));
 MUX2_X1 _0718_ (.A(_0184_),
    .B(_0185_),
    .S(_0224_),
    .Z(_0010_));
 AND2_X1 _0719_ (.A1(net36),
    .A2(_0183_),
    .ZN(_0225_));
 AND2_X1 _0720_ (.A1(net73),
    .A2(_0183_),
    .ZN(_0226_));
 MUX2_X1 _0721_ (.A(_0225_),
    .B(_0226_),
    .S(_0224_),
    .Z(_0011_));
 AND2_X1 _0722_ (.A1(net37),
    .A2(_0183_),
    .ZN(_0227_));
 NOR2_X1 _0723_ (.A1(_0132_),
    .A2(_0057_),
    .ZN(_0228_));
 MUX2_X1 _0724_ (.A(_0227_),
    .B(_0228_),
    .S(_0224_),
    .Z(_0012_));
 AND2_X1 _0725_ (.A1(net38),
    .A2(_0183_),
    .ZN(_0229_));
 AND2_X1 _0726_ (.A1(net75),
    .A2(_0183_),
    .ZN(_0230_));
 MUX2_X1 _0727_ (.A(_0229_),
    .B(_0230_),
    .S(_0224_),
    .Z(_0013_));
 AND2_X1 _0728_ (.A1(net39),
    .A2(_0183_),
    .ZN(_0231_));
 AND2_X1 _0729_ (.A1(net76),
    .A2(_0183_),
    .ZN(_0232_));
 MUX2_X1 _0730_ (.A(_0231_),
    .B(_0232_),
    .S(_0224_),
    .Z(_0014_));
 OAI21_X2 _0731_ (.A(_0055_),
    .B1(_0151_),
    .B2(_0073_),
    .ZN(_0233_));
 CLKBUF_X3 _0732_ (.A(_0233_),
    .Z(_0234_));
 BUF_X4 _0733_ (.A(_0208_),
    .Z(_0235_));
 CLKBUF_X3 _0734_ (.A(_0235_),
    .Z(_0236_));
 NOR2_X1 _0735_ (.A1(_0070_),
    .A2(_0094_),
    .ZN(_0237_));
 AOI21_X1 _0736_ (.A(_0065_),
    .B1(_0081_),
    .B2(_0084_),
    .ZN(_0238_));
 NOR2_X1 _0737_ (.A1(_0061_),
    .A2(_0238_),
    .ZN(_0239_));
 OAI21_X1 _0738_ (.A(_0061_),
    .B1(_0069_),
    .B2(_0086_),
    .ZN(_0240_));
 OAI221_X2 _0739_ (.A(_0063_),
    .B1(_0237_),
    .B2(_0239_),
    .C1(_0240_),
    .C2(_0222_),
    .ZN(_0241_));
 CLKBUF_X3 _0740_ (.A(_0241_),
    .Z(_0242_));
 CLKBUF_X3 _0741_ (.A(_0242_),
    .Z(_0243_));
 OAI21_X1 _0742_ (.A(net40),
    .B1(_0236_),
    .B2(_0243_),
    .ZN(_0244_));
 BUF_X4 _0743_ (.A(_0242_),
    .Z(_0245_));
 OR3_X1 _0744_ (.A1(net40),
    .A2(_0235_),
    .A3(_0245_),
    .ZN(_0246_));
 AOI21_X1 _0745_ (.A(_0234_),
    .B1(_0244_),
    .B2(_0246_),
    .ZN(_0015_));
 OR3_X2 _0746_ (.A1(_0186_),
    .A2(_0208_),
    .A3(_0241_),
    .ZN(_0247_));
 CLKBUF_X3 _0747_ (.A(_0247_),
    .Z(_0248_));
 INV_X1 _0748_ (.A(_0164_),
    .ZN(_0249_));
 INV_X1 _0749_ (.A(_0165_),
    .ZN(_0250_));
 NAND3_X2 _0750_ (.A1(_0523_),
    .A2(_0169_),
    .A3(_0170_),
    .ZN(_0251_));
 NAND2_X2 _0751_ (.A1(_0171_),
    .A2(_0172_),
    .ZN(_0252_));
 NOR4_X4 _0752_ (.A1(_0249_),
    .A2(_0250_),
    .A3(_0251_),
    .A4(_0252_),
    .ZN(_0253_));
 INV_X1 _0753_ (.A(_0166_),
    .ZN(_0254_));
 INV_X1 _0754_ (.A(_0167_),
    .ZN(_0255_));
 NOR2_X1 _0755_ (.A1(_0254_),
    .A2(_0255_),
    .ZN(_0256_));
 NOR2_X1 _0756_ (.A1(_0174_),
    .A2(_0057_),
    .ZN(_0257_));
 NAND3_X1 _0757_ (.A1(_0253_),
    .A2(_0256_),
    .A3(_0257_),
    .ZN(_0258_));
 CLKBUF_X3 _0758_ (.A(_0055_),
    .Z(_0259_));
 NAND2_X1 _0759_ (.A1(_0174_),
    .A2(_0259_),
    .ZN(_0260_));
 BUF_X4 _0760_ (.A(_0235_),
    .Z(_0261_));
 BUF_X4 _0761_ (.A(_0242_),
    .Z(_0262_));
 BUF_X4 _0762_ (.A(_0186_),
    .Z(_0263_));
 AOI21_X1 _0763_ (.A(_0263_),
    .B1(_0253_),
    .B2(_0256_),
    .ZN(_0264_));
 NOR3_X1 _0764_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0264_),
    .ZN(_0265_));
 OAI22_X1 _0765_ (.A1(_0248_),
    .A2(_0258_),
    .B1(_0260_),
    .B2(_0265_),
    .ZN(_0016_));
 NOR2_X1 _0766_ (.A1(_0073_),
    .A2(_0151_),
    .ZN(_0266_));
 NOR2_X1 _0767_ (.A1(_0056_),
    .A2(_0266_),
    .ZN(_0267_));
 BUF_X2 _0768_ (.A(_0267_),
    .Z(_0268_));
 AND2_X1 _0769_ (.A1(net42),
    .A2(_0268_),
    .ZN(_0269_));
 NOR2_X1 _0770_ (.A1(net42),
    .A2(_0234_),
    .ZN(_0270_));
 CLKBUF_X3 _0771_ (.A(_0235_),
    .Z(_0271_));
 NAND2_X2 _0772_ (.A1(net40),
    .A2(net51),
    .ZN(_0272_));
 NAND4_X1 _0773_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0171_),
    .A4(_0172_),
    .ZN(_0273_));
 NOR2_X1 _0774_ (.A1(_0272_),
    .A2(_0273_),
    .ZN(_0274_));
 AND4_X1 _0775_ (.A1(_0164_),
    .A2(_0165_),
    .A3(_0166_),
    .A4(_0274_),
    .ZN(_0275_));
 NAND3_X1 _0776_ (.A1(_0167_),
    .A2(_0174_),
    .A3(_0275_),
    .ZN(_0276_));
 NOR3_X1 _0777_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0276_),
    .ZN(_0277_));
 MUX2_X1 _0778_ (.A(_0269_),
    .B(_0270_),
    .S(_0277_),
    .Z(_0017_));
 NAND2_X1 _0779_ (.A1(_0166_),
    .A2(_0167_),
    .ZN(_0278_));
 NAND4_X2 _0780_ (.A1(_0164_),
    .A2(_0165_),
    .A3(_0174_),
    .A4(net42),
    .ZN(_0279_));
 OR4_X4 _0781_ (.A1(_0251_),
    .A2(_0252_),
    .A3(_0278_),
    .A4(_0279_),
    .ZN(_0280_));
 AND2_X1 _0782_ (.A1(_0095_),
    .A2(_0280_),
    .ZN(_0281_));
 NOR3_X1 _0783_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0281_),
    .ZN(_0282_));
 BUF_X4 _0784_ (.A(_0183_),
    .Z(_0283_));
 NAND2_X1 _0785_ (.A1(_0176_),
    .A2(_0283_),
    .ZN(_0284_));
 OR3_X1 _0786_ (.A1(_0176_),
    .A2(_0057_),
    .A3(_0280_),
    .ZN(_0285_));
 OAI22_X1 _0787_ (.A1(_0282_),
    .A2(_0284_),
    .B1(_0285_),
    .B2(_0248_),
    .ZN(_0018_));
 NOR2_X1 _0788_ (.A1(_0278_),
    .A2(_0279_),
    .ZN(_0286_));
 NAND3_X1 _0789_ (.A1(_0176_),
    .A2(_0274_),
    .A3(_0286_),
    .ZN(_0287_));
 AND2_X1 _0790_ (.A1(_0095_),
    .A2(_0287_),
    .ZN(_0288_));
 NOR3_X1 _0791_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0288_),
    .ZN(_0289_));
 NAND2_X1 _0792_ (.A1(net44),
    .A2(_0283_),
    .ZN(_0290_));
 OR3_X1 _0793_ (.A1(net44),
    .A2(_0057_),
    .A3(_0287_),
    .ZN(_0291_));
 OAI22_X1 _0794_ (.A1(_0289_),
    .A2(_0290_),
    .B1(_0291_),
    .B2(_0248_),
    .ZN(_0019_));
 CLKBUF_X3 _0795_ (.A(_0263_),
    .Z(_0292_));
 NAND2_X2 _0796_ (.A1(_0176_),
    .A2(net44),
    .ZN(_0293_));
 NOR2_X1 _0797_ (.A1(_0280_),
    .A2(_0293_),
    .ZN(_0294_));
 NOR2_X1 _0798_ (.A1(_0292_),
    .A2(_0294_),
    .ZN(_0295_));
 NOR3_X1 _0799_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0295_),
    .ZN(_0296_));
 NAND2_X1 _0800_ (.A1(net45),
    .A2(_0283_),
    .ZN(_0297_));
 INV_X1 _0801_ (.A(net45),
    .ZN(_0298_));
 NAND3_X1 _0802_ (.A1(_0298_),
    .A2(_0259_),
    .A3(_0294_),
    .ZN(_0299_));
 OAI22_X1 _0803_ (.A1(_0296_),
    .A2(_0297_),
    .B1(_0299_),
    .B2(_0248_),
    .ZN(_0020_));
 NOR2_X1 _0804_ (.A1(_0298_),
    .A2(_0293_),
    .ZN(_0300_));
 AND3_X1 _0805_ (.A1(_0274_),
    .A2(_0286_),
    .A3(_0300_),
    .ZN(_0301_));
 NOR2_X1 _0806_ (.A1(_0292_),
    .A2(_0301_),
    .ZN(_0302_));
 NOR3_X1 _0807_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0302_),
    .ZN(_0303_));
 NAND2_X1 _0808_ (.A1(net46),
    .A2(_0283_),
    .ZN(_0304_));
 INV_X1 _0809_ (.A(net46),
    .ZN(_0305_));
 CLKBUF_X3 _0810_ (.A(_0055_),
    .Z(_0306_));
 NAND3_X1 _0811_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0301_),
    .ZN(_0307_));
 OAI22_X1 _0812_ (.A1(_0303_),
    .A2(_0304_),
    .B1(_0307_),
    .B2(_0248_),
    .ZN(_0021_));
 NAND2_X1 _0813_ (.A1(net45),
    .A2(net46),
    .ZN(_0308_));
 NOR3_X1 _0814_ (.A1(_0280_),
    .A2(_0293_),
    .A3(_0308_),
    .ZN(_0309_));
 NOR2_X1 _0815_ (.A1(_0292_),
    .A2(_0309_),
    .ZN(_0310_));
 NOR3_X1 _0816_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0310_),
    .ZN(_0311_));
 NAND2_X1 _0817_ (.A1(net47),
    .A2(_0283_),
    .ZN(_0312_));
 INV_X1 _0818_ (.A(net47),
    .ZN(_0313_));
 NAND3_X1 _0819_ (.A1(_0313_),
    .A2(_0306_),
    .A3(_0309_),
    .ZN(_0314_));
 OAI22_X1 _0820_ (.A1(_0311_),
    .A2(_0312_),
    .B1(_0314_),
    .B2(_0248_),
    .ZN(_0022_));
 NOR2_X1 _0821_ (.A1(_0235_),
    .A2(_0242_),
    .ZN(_0315_));
 NOR2_X1 _0822_ (.A1(_0305_),
    .A2(_0313_),
    .ZN(_0316_));
 AND4_X1 _0823_ (.A1(_0274_),
    .A2(_0286_),
    .A3(_0300_),
    .A4(_0316_),
    .ZN(_0317_));
 BUF_X2 _0824_ (.A(_0317_),
    .Z(_0318_));
 OAI21_X1 _0825_ (.A(_0177_),
    .B1(_0186_),
    .B2(_0318_),
    .ZN(_0319_));
 INV_X1 _0826_ (.A(_0319_),
    .ZN(_0320_));
 NAND2_X1 _0827_ (.A1(_0301_),
    .A2(_0316_),
    .ZN(_0321_));
 OR4_X1 _0828_ (.A1(_0186_),
    .A2(_0208_),
    .A3(_0241_),
    .A4(_0321_),
    .ZN(_0322_));
 INV_X1 _0829_ (.A(_0177_),
    .ZN(_0323_));
 AOI221_X1 _0830_ (.A(_0057_),
    .B1(_0315_),
    .B2(_0320_),
    .C1(_0322_),
    .C2(_0323_),
    .ZN(_0023_));
 INV_X1 _0831_ (.A(net49),
    .ZN(_0324_));
 NOR4_X4 _0832_ (.A1(_0313_),
    .A2(_0280_),
    .A3(_0293_),
    .A4(_0308_),
    .ZN(_0325_));
 NAND4_X1 _0833_ (.A1(_0177_),
    .A2(_0324_),
    .A3(_0055_),
    .A4(_0325_),
    .ZN(_0326_));
 OR4_X1 _0834_ (.A1(_0292_),
    .A2(_0235_),
    .A3(_0242_),
    .A4(_0326_),
    .ZN(_0327_));
 NAND2_X1 _0835_ (.A1(net49),
    .A2(_0283_),
    .ZN(_0328_));
 AOI21_X1 _0836_ (.A(_0263_),
    .B1(_0325_),
    .B2(_0177_),
    .ZN(_0329_));
 NOR3_X1 _0837_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0329_),
    .ZN(_0330_));
 OAI21_X1 _0838_ (.A(_0327_),
    .B1(_0328_),
    .B2(_0330_),
    .ZN(_0024_));
 NOR2_X1 _0839_ (.A1(_0323_),
    .A2(_0324_),
    .ZN(_0331_));
 NOR2_X1 _0840_ (.A1(_0160_),
    .A2(_0057_),
    .ZN(_0332_));
 NAND3_X1 _0841_ (.A1(_0318_),
    .A2(_0331_),
    .A3(_0332_),
    .ZN(_0333_));
 OR4_X1 _0842_ (.A1(_0292_),
    .A2(_0235_),
    .A3(_0242_),
    .A4(_0333_),
    .ZN(_0334_));
 NAND2_X1 _0843_ (.A1(_0160_),
    .A2(_0283_),
    .ZN(_0335_));
 AOI21_X1 _0844_ (.A(_0263_),
    .B1(_0318_),
    .B2(_0331_),
    .ZN(_0336_));
 NOR3_X1 _0845_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0336_),
    .ZN(_0337_));
 OAI21_X1 _0846_ (.A(_0334_),
    .B1(_0335_),
    .B2(_0337_),
    .ZN(_0025_));
 OAI21_X1 _0847_ (.A(net51),
    .B1(_0236_),
    .B2(_0243_),
    .ZN(_0338_));
 NAND2_X1 _0848_ (.A1(_0522_),
    .A2(_0095_),
    .ZN(_0339_));
 OR3_X1 _0849_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0339_),
    .ZN(_0340_));
 AOI21_X1 _0850_ (.A(_0058_),
    .B1(_0338_),
    .B2(_0340_),
    .ZN(_0026_));
 AND2_X1 _0851_ (.A1(_0160_),
    .A2(_0331_),
    .ZN(_0341_));
 NOR2_X1 _0852_ (.A1(net52),
    .A2(_0056_),
    .ZN(_0342_));
 NAND3_X1 _0853_ (.A1(_0325_),
    .A2(_0341_),
    .A3(_0342_),
    .ZN(_0343_));
 OR4_X1 _0854_ (.A1(_0292_),
    .A2(_0235_),
    .A3(_0242_),
    .A4(_0343_),
    .ZN(_0344_));
 NAND2_X1 _0855_ (.A1(net52),
    .A2(_0283_),
    .ZN(_0345_));
 AOI21_X1 _0856_ (.A(_0263_),
    .B1(_0325_),
    .B2(_0341_),
    .ZN(_0346_));
 NOR3_X1 _0857_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0346_),
    .ZN(_0347_));
 OAI21_X1 _0858_ (.A(_0344_),
    .B1(_0345_),
    .B2(_0347_),
    .ZN(_0027_));
 AND2_X1 _0859_ (.A1(_0161_),
    .A2(_0268_),
    .ZN(_0348_));
 NOR2_X1 _0860_ (.A1(_0161_),
    .A2(_0234_),
    .ZN(_0349_));
 AND4_X1 _0861_ (.A1(_0177_),
    .A2(net49),
    .A3(_0160_),
    .A4(net52),
    .ZN(_0350_));
 NAND2_X1 _0862_ (.A1(_0318_),
    .A2(_0350_),
    .ZN(_0351_));
 NOR3_X1 _0863_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0351_),
    .ZN(_0352_));
 MUX2_X1 _0864_ (.A(_0348_),
    .B(_0349_),
    .S(_0352_),
    .Z(_0028_));
 AND2_X1 _0865_ (.A1(net54),
    .A2(_0268_),
    .ZN(_0353_));
 NOR2_X1 _0866_ (.A1(net54),
    .A2(_0234_),
    .ZN(_0354_));
 NAND3_X1 _0867_ (.A1(_0161_),
    .A2(_0325_),
    .A3(_0350_),
    .ZN(_0355_));
 NOR3_X1 _0868_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0355_),
    .ZN(_0356_));
 MUX2_X1 _0869_ (.A(_0353_),
    .B(_0354_),
    .S(_0356_),
    .Z(_0029_));
 AND2_X1 _0870_ (.A1(net55),
    .A2(_0268_),
    .ZN(_0357_));
 NOR2_X1 _0871_ (.A1(net55),
    .A2(_0234_),
    .ZN(_0358_));
 AND3_X1 _0872_ (.A1(_0161_),
    .A2(net54),
    .A3(_0350_),
    .ZN(_0359_));
 NAND2_X1 _0873_ (.A1(_0318_),
    .A2(_0359_),
    .ZN(_0360_));
 NOR3_X1 _0874_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0360_),
    .ZN(_0361_));
 MUX2_X1 _0875_ (.A(_0357_),
    .B(_0358_),
    .S(_0361_),
    .Z(_0030_));
 AND2_X1 _0876_ (.A1(_0157_),
    .A2(_0268_),
    .ZN(_0362_));
 NOR2_X1 _0877_ (.A1(_0157_),
    .A2(_0234_),
    .ZN(_0363_));
 AND2_X1 _0878_ (.A1(net55),
    .A2(_0359_),
    .ZN(_0364_));
 BUF_X2 _0879_ (.A(_0364_),
    .Z(_0365_));
 NAND2_X1 _0880_ (.A1(_0325_),
    .A2(_0365_),
    .ZN(_0366_));
 NOR3_X1 _0881_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0366_),
    .ZN(_0367_));
 MUX2_X1 _0882_ (.A(_0362_),
    .B(_0363_),
    .S(_0367_),
    .Z(_0031_));
 AND2_X1 _0883_ (.A1(_0158_),
    .A2(_0268_),
    .ZN(_0368_));
 NOR2_X1 _0884_ (.A1(_0158_),
    .A2(_0234_),
    .ZN(_0369_));
 NAND3_X1 _0885_ (.A1(_0157_),
    .A2(_0318_),
    .A3(_0365_),
    .ZN(_0370_));
 NOR3_X1 _0886_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0370_),
    .ZN(_0371_));
 MUX2_X1 _0887_ (.A(_0368_),
    .B(_0369_),
    .S(_0371_),
    .Z(_0032_));
 AND2_X1 _0888_ (.A1(net58),
    .A2(_0268_),
    .ZN(_0372_));
 NOR2_X1 _0889_ (.A1(net58),
    .A2(_0234_),
    .ZN(_0373_));
 NAND4_X1 _0890_ (.A1(_0157_),
    .A2(_0158_),
    .A3(_0325_),
    .A4(_0365_),
    .ZN(_0374_));
 NOR3_X1 _0891_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0374_),
    .ZN(_0375_));
 MUX2_X1 _0892_ (.A(_0372_),
    .B(_0373_),
    .S(_0375_),
    .Z(_0033_));
 AND2_X1 _0893_ (.A1(net59),
    .A2(_0268_),
    .ZN(_0376_));
 NOR2_X1 _0894_ (.A1(net59),
    .A2(_0234_),
    .ZN(_0377_));
 AND3_X1 _0895_ (.A1(_0157_),
    .A2(_0158_),
    .A3(net58),
    .ZN(_0378_));
 NAND3_X1 _0896_ (.A1(_0318_),
    .A2(_0365_),
    .A3(_0378_),
    .ZN(_0379_));
 NOR3_X1 _0897_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0379_),
    .ZN(_0380_));
 MUX2_X1 _0898_ (.A(_0376_),
    .B(_0377_),
    .S(_0380_),
    .Z(_0034_));
 AND2_X1 _0899_ (.A1(_0155_),
    .A2(_0268_),
    .ZN(_0381_));
 NOR2_X1 _0900_ (.A1(_0155_),
    .A2(_0234_),
    .ZN(_0382_));
 AND2_X1 _0901_ (.A1(net59),
    .A2(_0378_),
    .ZN(_0383_));
 NAND3_X1 _0902_ (.A1(_0325_),
    .A2(_0365_),
    .A3(_0383_),
    .ZN(_0384_));
 NOR3_X1 _0903_ (.A1(_0271_),
    .A2(_0245_),
    .A3(_0384_),
    .ZN(_0385_));
 MUX2_X1 _0904_ (.A(_0381_),
    .B(_0382_),
    .S(_0385_),
    .Z(_0035_));
 AND2_X1 _0905_ (.A1(net61),
    .A2(_0268_),
    .ZN(_0386_));
 NOR2_X1 _0906_ (.A1(net61),
    .A2(_0233_),
    .ZN(_0387_));
 NAND4_X1 _0907_ (.A1(_0155_),
    .A2(_0318_),
    .A3(_0365_),
    .A4(_0383_),
    .ZN(_0388_));
 NOR3_X1 _0908_ (.A1(_0271_),
    .A2(_0242_),
    .A3(_0388_),
    .ZN(_0389_));
 MUX2_X1 _0909_ (.A(_0386_),
    .B(_0387_),
    .S(_0389_),
    .Z(_0036_));
 NOR2_X1 _0910_ (.A1(_0523_),
    .A2(_0263_),
    .ZN(_0390_));
 NOR3_X1 _0911_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0390_),
    .ZN(_0391_));
 NAND2_X1 _0912_ (.A1(_0169_),
    .A2(_0259_),
    .ZN(_0392_));
 INV_X1 _0913_ (.A(_0169_),
    .ZN(_0393_));
 NAND3_X1 _0914_ (.A1(_0523_),
    .A2(_0393_),
    .A3(_0306_),
    .ZN(_0394_));
 OAI22_X1 _0915_ (.A1(_0391_),
    .A2(_0392_),
    .B1(_0394_),
    .B2(_0248_),
    .ZN(_0037_));
 AND2_X1 _0916_ (.A1(net63),
    .A2(_0267_),
    .ZN(_0395_));
 NOR2_X1 _0917_ (.A1(net63),
    .A2(_0233_),
    .ZN(_0396_));
 AND3_X1 _0918_ (.A1(_0155_),
    .A2(net61),
    .A3(_0383_),
    .ZN(_0397_));
 NAND3_X1 _0919_ (.A1(_0325_),
    .A2(_0365_),
    .A3(_0397_),
    .ZN(_0398_));
 NOR3_X1 _0920_ (.A1(_0235_),
    .A2(_0242_),
    .A3(_0398_),
    .ZN(_0399_));
 MUX2_X1 _0921_ (.A(_0395_),
    .B(_0396_),
    .S(_0399_),
    .Z(_0038_));
 AND2_X1 _0922_ (.A1(net64),
    .A2(_0267_),
    .ZN(_0400_));
 NOR2_X1 _0923_ (.A1(net64),
    .A2(_0233_),
    .ZN(_0401_));
 AND4_X1 _0924_ (.A1(_0155_),
    .A2(net61),
    .A3(net63),
    .A4(_0383_),
    .ZN(_0402_));
 NAND3_X1 _0925_ (.A1(_0318_),
    .A2(_0365_),
    .A3(_0402_),
    .ZN(_0403_));
 NOR3_X1 _0926_ (.A1(_0235_),
    .A2(_0242_),
    .A3(_0403_),
    .ZN(_0404_));
 MUX2_X1 _0927_ (.A(_0400_),
    .B(_0401_),
    .S(_0404_),
    .Z(_0039_));
 NOR2_X1 _0928_ (.A1(_0393_),
    .A2(_0272_),
    .ZN(_0405_));
 NOR2_X1 _0929_ (.A1(_0292_),
    .A2(_0405_),
    .ZN(_0406_));
 NOR3_X1 _0930_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0406_),
    .ZN(_0407_));
 NAND2_X1 _0931_ (.A1(_0170_),
    .A2(_0259_),
    .ZN(_0408_));
 INV_X1 _0932_ (.A(_0170_),
    .ZN(_0409_));
 NAND3_X1 _0933_ (.A1(_0409_),
    .A2(_0306_),
    .A3(_0405_),
    .ZN(_0410_));
 OAI22_X1 _0934_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0410_),
    .B2(_0248_),
    .ZN(_0040_));
 AND3_X1 _0935_ (.A1(_0523_),
    .A2(_0169_),
    .A3(_0170_),
    .ZN(_0411_));
 NOR2_X1 _0936_ (.A1(_0292_),
    .A2(_0411_),
    .ZN(_0412_));
 NOR3_X1 _0937_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0412_),
    .ZN(_0413_));
 NAND2_X1 _0938_ (.A1(_0171_),
    .A2(_0259_),
    .ZN(_0414_));
 INV_X1 _0939_ (.A(_0171_),
    .ZN(_0415_));
 NAND3_X1 _0940_ (.A1(_0415_),
    .A2(_0306_),
    .A3(_0411_),
    .ZN(_0416_));
 OAI22_X1 _0941_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0416_),
    .B2(_0248_),
    .ZN(_0041_));
 NOR4_X2 _0942_ (.A1(_0393_),
    .A2(_0409_),
    .A3(_0415_),
    .A4(_0272_),
    .ZN(_0417_));
 NOR2_X1 _0943_ (.A1(_0292_),
    .A2(_0417_),
    .ZN(_0418_));
 NOR3_X1 _0944_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0418_),
    .ZN(_0419_));
 NAND2_X1 _0945_ (.A1(_0172_),
    .A2(_0259_),
    .ZN(_0420_));
 INV_X1 _0946_ (.A(_0172_),
    .ZN(_0421_));
 NAND3_X1 _0947_ (.A1(_0421_),
    .A2(_0306_),
    .A3(_0417_),
    .ZN(_0422_));
 OAI22_X1 _0948_ (.A1(_0419_),
    .A2(_0420_),
    .B1(_0422_),
    .B2(_0248_),
    .ZN(_0042_));
 NOR2_X1 _0949_ (.A1(_0251_),
    .A2(_0252_),
    .ZN(_0423_));
 NOR2_X1 _0950_ (.A1(_0292_),
    .A2(_0423_),
    .ZN(_0424_));
 NOR3_X1 _0951_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0424_),
    .ZN(_0425_));
 NAND2_X1 _0952_ (.A1(_0164_),
    .A2(_0259_),
    .ZN(_0426_));
 NAND3_X1 _0953_ (.A1(_0249_),
    .A2(_0306_),
    .A3(_0423_),
    .ZN(_0427_));
 OAI22_X1 _0954_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0427_),
    .B2(_0247_),
    .ZN(_0043_));
 NOR3_X1 _0955_ (.A1(_0249_),
    .A2(_0272_),
    .A3(_0273_),
    .ZN(_0428_));
 NOR2_X1 _0956_ (.A1(_0263_),
    .A2(_0428_),
    .ZN(_0429_));
 NOR3_X1 _0957_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0429_),
    .ZN(_0430_));
 NAND2_X1 _0958_ (.A1(_0165_),
    .A2(_0259_),
    .ZN(_0431_));
 NAND3_X1 _0959_ (.A1(_0250_),
    .A2(_0306_),
    .A3(_0428_),
    .ZN(_0432_));
 OAI22_X1 _0960_ (.A1(_0430_),
    .A2(_0431_),
    .B1(_0432_),
    .B2(_0247_),
    .ZN(_0044_));
 NOR2_X1 _0961_ (.A1(_0263_),
    .A2(_0253_),
    .ZN(_0433_));
 NOR3_X1 _0962_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0433_),
    .ZN(_0434_));
 NAND2_X1 _0963_ (.A1(_0166_),
    .A2(_0259_),
    .ZN(_0435_));
 NAND3_X1 _0964_ (.A1(_0254_),
    .A2(_0306_),
    .A3(_0253_),
    .ZN(_0436_));
 OAI22_X1 _0965_ (.A1(_0434_),
    .A2(_0435_),
    .B1(_0436_),
    .B2(_0247_),
    .ZN(_0045_));
 NOR2_X1 _0966_ (.A1(_0263_),
    .A2(_0275_),
    .ZN(_0437_));
 NOR3_X1 _0967_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0437_),
    .ZN(_0438_));
 NAND2_X1 _0968_ (.A1(_0167_),
    .A2(_0259_),
    .ZN(_0439_));
 NAND3_X1 _0969_ (.A1(_0255_),
    .A2(_0306_),
    .A3(_0275_),
    .ZN(_0440_));
 OAI22_X1 _0970_ (.A1(_0438_),
    .A2(_0439_),
    .B1(_0440_),
    .B2(_0247_),
    .ZN(_0046_));
 AOI21_X1 _0971_ (.A(_0076_),
    .B1(_0091_),
    .B2(_0066_),
    .ZN(_0441_));
 MUX2_X1 _0972_ (.A(_0077_),
    .B(_0441_),
    .S(_0187_),
    .Z(_0442_));
 OAI21_X1 _0973_ (.A(_0083_),
    .B1(_0263_),
    .B2(_0442_),
    .ZN(_0443_));
 NAND3_X1 _0974_ (.A1(_0086_),
    .A2(_0090_),
    .A3(_0097_),
    .ZN(_0444_));
 MUX2_X1 _0975_ (.A(_0070_),
    .B(_0091_),
    .S(_0074_),
    .Z(_0445_));
 OAI21_X1 _0976_ (.A(_0444_),
    .B1(_0445_),
    .B2(_0097_),
    .ZN(_0446_));
 NOR2_X1 _0977_ (.A1(_0061_),
    .A2(_0075_),
    .ZN(_0447_));
 AOI22_X1 _0978_ (.A1(_0063_),
    .A2(_0446_),
    .B1(_0447_),
    .B2(_0116_),
    .ZN(_0448_));
 OR2_X1 _0979_ (.A1(_0443_),
    .A2(_0448_),
    .ZN(_0449_));
 NAND2_X1 _0980_ (.A1(_0075_),
    .A2(_0443_),
    .ZN(_0450_));
 AOI21_X1 _0981_ (.A(_0058_),
    .B1(_0449_),
    .B2(_0450_),
    .ZN(_0047_));
 INV_X1 _0982_ (.A(_0061_),
    .ZN(_0451_));
 AOI21_X1 _0983_ (.A(_0073_),
    .B1(_0238_),
    .B2(_0451_),
    .ZN(_0452_));
 OR2_X1 _0984_ (.A1(_0209_),
    .A2(_0452_),
    .ZN(_0453_));
 AOI21_X1 _0985_ (.A(_0058_),
    .B1(_0192_),
    .B2(_0453_),
    .ZN(_0048_));
 OAI22_X2 _0986_ (.A1(_0066_),
    .A2(_0117_),
    .B1(_0089_),
    .B2(_0116_),
    .ZN(_0454_));
 NAND3_X1 _0987_ (.A1(_0073_),
    .A2(_0081_),
    .A3(_0149_),
    .ZN(_0455_));
 NOR2_X1 _0988_ (.A1(_0067_),
    .A2(_0088_),
    .ZN(_0456_));
 OAI21_X1 _0989_ (.A(_0063_),
    .B1(_0082_),
    .B2(_0456_),
    .ZN(_0457_));
 NAND4_X2 _0990_ (.A1(_0115_),
    .A2(_0454_),
    .A3(_0455_),
    .A4(_0457_),
    .ZN(_0458_));
 MUX2_X1 _0991_ (.A(_0205_),
    .B(_0061_),
    .S(_0458_),
    .Z(_0459_));
 AND2_X1 _0992_ (.A1(_0283_),
    .A2(_0459_),
    .ZN(_0049_));
 OAI21_X1 _0993_ (.A(_0069_),
    .B1(_0205_),
    .B2(_0458_),
    .ZN(_0460_));
 OR3_X1 _0994_ (.A1(_0069_),
    .A2(_0064_),
    .A3(_0458_),
    .ZN(_0461_));
 AOI21_X1 _0995_ (.A(_0058_),
    .B1(_0460_),
    .B2(_0461_),
    .ZN(_0050_));
 NAND3_X1 _0996_ (.A1(_0063_),
    .A2(_0074_),
    .A3(_0189_),
    .ZN(_0462_));
 MUX2_X1 _0997_ (.A(_0462_),
    .B(_0074_),
    .S(_0458_),
    .Z(_0463_));
 NAND3_X1 _0998_ (.A1(_0063_),
    .A2(_0086_),
    .A3(_0097_),
    .ZN(_0464_));
 AOI21_X1 _0999_ (.A(_0057_),
    .B1(_0463_),
    .B2(_0464_),
    .ZN(_0051_));
 OR3_X1 _1000_ (.A1(_0073_),
    .A2(_0187_),
    .A3(_0458_),
    .ZN(_0465_));
 AOI21_X1 _1001_ (.A(_0057_),
    .B1(_0455_),
    .B2(_0465_),
    .ZN(_0052_));
 MUX2_X1 _1002_ (.A(_0084_),
    .B(_0189_),
    .S(_0074_),
    .Z(_0466_));
 NAND2_X1 _1003_ (.A1(_0071_),
    .A2(_0466_),
    .ZN(_0467_));
 NOR2_X1 _1004_ (.A1(_0074_),
    .A2(_0070_),
    .ZN(_0468_));
 NOR3_X1 _1005_ (.A1(_0084_),
    .A2(_0086_),
    .A3(_0075_),
    .ZN(_0469_));
 OAI21_X1 _1006_ (.A(_0451_),
    .B1(_0468_),
    .B2(_0469_),
    .ZN(_0470_));
 AOI21_X1 _1007_ (.A(_0073_),
    .B1(_0467_),
    .B2(_0470_),
    .ZN(_0471_));
 NAND2_X1 _1008_ (.A1(_0189_),
    .A2(_0204_),
    .ZN(_0472_));
 OAI21_X1 _1009_ (.A(_0086_),
    .B1(_0189_),
    .B2(_0204_),
    .ZN(_0473_));
 NAND3_X1 _1010_ (.A1(_0083_),
    .A2(_0472_),
    .A3(_0473_),
    .ZN(_0474_));
 MUX2_X1 _1011_ (.A(_0471_),
    .B(_0090_),
    .S(_0474_),
    .Z(_0475_));
 AND2_X1 _1012_ (.A1(_0283_),
    .A2(_0475_),
    .ZN(_0053_));
 OAI21_X1 _1013_ (.A(_0109_),
    .B1(_0063_),
    .B2(_0451_),
    .ZN(net77));
 OAI21_X4 _1014_ (.A(_0205_),
    .B1(_0086_),
    .B2(_0069_),
    .ZN(net102));
 HA_X1 _1015_ (.A(_0519_),
    .B(_0520_),
    .CO(_0521_),
    .S(_0522_));
 HA_X1 _1016_ (.A(net40),
    .B(net51),
    .CO(_0523_),
    .S(_0524_));
 HA_X1 _1017_ (.A(_0525_),
    .B(_0526_),
    .CO(_0527_),
    .S(_0528_));
 HA_X1 _1018_ (.A(net72),
    .B(net73),
    .CO(_0529_),
    .S(_0530_));
 HA_X1 _1019_ (.A(_0531_),
    .B(_0532_),
    .CO(_0533_),
    .S(_0534_));
 HA_X1 _1020_ (.A(net76),
    .B(_0535_),
    .CO(_0536_),
    .S(_0537_));
 BUF_X1 _1021_ (.A(net102),
    .Z(net78));
 BUF_X1 _1022_ (.A(net102),
    .Z(net89));
 BUF_X1 _1023_ (.A(net102),
    .Z(net100));
 BUF_X1 _1024_ (.A(net102),
    .Z(net103));
 BUF_X1 _1025_ (.A(net102),
    .Z(net104));
 BUF_X1 _1026_ (.A(net102),
    .Z(net105));
 BUF_X1 _1027_ (.A(net102),
    .Z(net106));
 BUF_X1 _1028_ (.A(net102),
    .Z(net107));
 BUF_X1 _1029_ (.A(net102),
    .Z(net108));
 BUF_X1 _1030_ (.A(net102),
    .Z(net109));
 BUF_X1 _1031_ (.A(net102),
    .Z(net79));
 BUF_X1 _1032_ (.A(net102),
    .Z(net80));
 BUF_X1 _1033_ (.A(net102),
    .Z(net81));
 BUF_X1 _1034_ (.A(net102),
    .Z(net82));
 BUF_X1 _1035_ (.A(net102),
    .Z(net83));
 BUF_X1 _1036_ (.A(net102),
    .Z(net84));
 BUF_X1 _1037_ (.A(net102),
    .Z(net85));
 BUF_X1 _1038_ (.A(net102),
    .Z(net86));
 BUF_X1 _1039_ (.A(net102),
    .Z(net87));
 BUF_X1 _1040_ (.A(net102),
    .Z(net88));
 BUF_X1 _1041_ (.A(net102),
    .Z(net90));
 BUF_X1 _1042_ (.A(net102),
    .Z(net91));
 BUF_X1 _1043_ (.A(net102),
    .Z(net92));
 BUF_X1 _1044_ (.A(net102),
    .Z(net93));
 BUF_X1 _1045_ (.A(net102),
    .Z(net94));
 BUF_X1 _1046_ (.A(net102),
    .Z(net95));
 BUF_X1 _1047_ (.A(net102),
    .Z(net96));
 BUF_X1 _1048_ (.A(net102),
    .Z(net97));
 BUF_X1 _1049_ (.A(net102),
    .Z(net98));
 BUF_X1 _1050_ (.A(net102),
    .Z(net99));
 BUF_X1 _1051_ (.A(net102),
    .Z(net101));
 DFF_X1 \addr_counter[0]$_SDFFE_PN0P_  (.D(_0003_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net72),
    .QN(_0525_));
 DFF_X2 \addr_counter[1]$_SDFFE_PN0P_  (.D(_0004_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net73),
    .QN(_0526_));
 DFF_X1 \addr_counter[2]$_SDFFE_PN0P_  (.D(_0005_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net74),
    .QN(_0518_));
 DFF_X2 \addr_counter[3]$_SDFFE_PN0P_  (.D(_0006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net75),
    .QN(_0002_));
 DFF_X2 \addr_counter[4]$_SDFFE_PN0P_  (.D(_0007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net76),
    .QN(_0531_));
 DFF_X1 \bist_done$_SDFFE_PN0P_  (.D(_0008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net33),
    .QN(_0517_));
 DFF_X1 \bist_pass$_SDFFE_PN0P_  (.D(_0009_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net34),
    .QN(_0516_));
 DFF_X1 \error_addr[0]$_SDFFE_PN0P_  (.D(_0010_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net35),
    .QN(_0515_));
 DFF_X1 \error_addr[1]$_SDFFE_PN0P_  (.D(_0011_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net36),
    .QN(_0514_));
 DFF_X1 \error_addr[2]$_SDFFE_PN0P_  (.D(_0012_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net37),
    .QN(_0513_));
 DFF_X1 \error_addr[3]$_SDFFE_PN0P_  (.D(_0013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net38),
    .QN(_0512_));
 DFF_X1 \error_addr[4]$_SDFFE_PN0P_  (.D(_0014_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net39),
    .QN(_0511_));
 DFF_X2 \error_count[0]$_SDFFE_PN0P_  (.D(_0015_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net40),
    .QN(_0519_));
 DFF_X1 \error_count[10]$_SDFFE_PN0P_  (.D(_0016_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net41),
    .QN(_0510_));
 DFF_X2 \error_count[11]$_SDFFE_PN0P_  (.D(_0017_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net42),
    .QN(_0509_));
 DFF_X1 \error_count[12]$_SDFFE_PN0P_  (.D(_0018_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net43),
    .QN(_0508_));
 DFF_X2 \error_count[13]$_SDFFE_PN0P_  (.D(_0019_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net44),
    .QN(_0507_));
 DFF_X1 \error_count[14]$_SDFFE_PN0P_  (.D(_0020_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net45),
    .QN(_0506_));
 DFF_X2 \error_count[15]$_SDFFE_PN0P_  (.D(_0021_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net46),
    .QN(_0505_));
 DFF_X1 \error_count[16]$_SDFFE_PN0P_  (.D(_0022_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net47),
    .QN(_0504_));
 DFF_X1 \error_count[17]$_SDFFE_PN0P_  (.D(_0023_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net48),
    .QN(_0503_));
 DFF_X2 \error_count[18]$_SDFFE_PN0P_  (.D(_0024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net49),
    .QN(_0502_));
 DFF_X1 \error_count[19]$_SDFFE_PN0P_  (.D(_0025_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net50),
    .QN(_0501_));
 DFF_X2 \error_count[1]$_SDFFE_PN0P_  (.D(_0026_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net51),
    .QN(_0520_));
 DFF_X1 \error_count[20]$_SDFFE_PN0P_  (.D(_0027_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net52),
    .QN(_0500_));
 DFF_X1 \error_count[21]$_SDFFE_PN0P_  (.D(_0028_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net53),
    .QN(_0499_));
 DFF_X1 \error_count[22]$_SDFFE_PN0P_  (.D(_0029_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net54),
    .QN(_0498_));
 DFF_X1 \error_count[23]$_SDFFE_PN0P_  (.D(_0030_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net55),
    .QN(_0497_));
 DFF_X1 \error_count[24]$_SDFFE_PN0P_  (.D(_0031_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net56),
    .QN(_0496_));
 DFF_X1 \error_count[25]$_SDFFE_PN0P_  (.D(_0032_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net57),
    .QN(_0495_));
 DFF_X1 \error_count[26]$_SDFFE_PN0P_  (.D(_0033_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net58),
    .QN(_0494_));
 DFF_X1 \error_count[27]$_SDFFE_PN0P_  (.D(_0034_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net59),
    .QN(_0493_));
 DFF_X1 \error_count[28]$_SDFFE_PN0P_  (.D(_0035_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net60),
    .QN(_0492_));
 DFF_X1 \error_count[29]$_SDFFE_PN0P_  (.D(_0036_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net61),
    .QN(_0491_));
 DFF_X1 \error_count[2]$_SDFFE_PN0P_  (.D(_0037_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net62),
    .QN(_0490_));
 DFF_X1 \error_count[30]$_SDFFE_PN0P_  (.D(_0038_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net63),
    .QN(_0489_));
 DFF_X1 \error_count[31]$_SDFFE_PN0P_  (.D(_0039_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net64),
    .QN(_0488_));
 DFF_X1 \error_count[3]$_SDFFE_PN0P_  (.D(_0040_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net65),
    .QN(_0487_));
 DFF_X1 \error_count[4]$_SDFFE_PN0P_  (.D(_0041_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net66),
    .QN(_0486_));
 DFF_X1 \error_count[5]$_SDFFE_PN0P_  (.D(_0042_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net67),
    .QN(_0485_));
 DFF_X1 \error_count[6]$_SDFFE_PN0P_  (.D(_0043_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net68),
    .QN(_0484_));
 DFF_X1 \error_count[7]$_SDFFE_PN0P_  (.D(_0044_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net69),
    .QN(_0483_));
 DFF_X1 \error_count[8]$_SDFFE_PN0P_  (.D(_0045_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net70),
    .QN(_0482_));
 DFF_X1 \error_count[9]$_SDFFE_PN0P_  (.D(_0046_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net71),
    .QN(_0481_));
 DFF_X1 \phase_complete$_SDFFE_PN0P_  (.D(_0047_),
    .CK(clknet_2_0__leaf_clk),
    .Q(phase_complete),
    .QN(_0001_));
 DFF_X1 \read_phase$_SDFFE_PN0P_  (.D(_0048_),
    .CK(clknet_2_1__leaf_clk),
    .Q(read_phase),
    .QN(_0000_));
 DFF_X1 \state[0]$_SDFFE_PN0P_  (.D(_0049_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[0] ),
    .QN(_0480_));
 DFF_X1 \state[1]$_SDFFE_PN0P_  (.D(_0050_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[1] ),
    .QN(_0479_));
 DFF_X1 \state[2]$_SDFFE_PN0P_  (.D(_0051_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[2] ),
    .QN(_0478_));
 DFF_X1 \state[3]$_SDFFE_PN0P_  (.D(_0052_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[3] ),
    .QN(_0477_));
 DFF_X1 \write_phase$_SDFFE_PN0P_  (.D(_0053_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net110),
    .QN(_0476_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_55 ();
 BUF_X1 input1 (.A(mem_rdata[0]),
    .Z(net1));
 BUF_X1 input2 (.A(mem_rdata[10]),
    .Z(net2));
 BUF_X1 input3 (.A(mem_rdata[11]),
    .Z(net3));
 BUF_X1 input4 (.A(mem_rdata[12]),
    .Z(net4));
 BUF_X1 input5 (.A(mem_rdata[13]),
    .Z(net5));
 BUF_X1 input6 (.A(mem_rdata[14]),
    .Z(net6));
 BUF_X1 input7 (.A(mem_rdata[15]),
    .Z(net7));
 BUF_X1 input8 (.A(mem_rdata[16]),
    .Z(net8));
 BUF_X1 input9 (.A(mem_rdata[17]),
    .Z(net9));
 BUF_X1 input10 (.A(mem_rdata[18]),
    .Z(net10));
 BUF_X1 input11 (.A(mem_rdata[19]),
    .Z(net11));
 BUF_X1 input12 (.A(mem_rdata[1]),
    .Z(net12));
 BUF_X1 input13 (.A(mem_rdata[20]),
    .Z(net13));
 BUF_X1 input14 (.A(mem_rdata[21]),
    .Z(net14));
 BUF_X1 input15 (.A(mem_rdata[22]),
    .Z(net15));
 BUF_X1 input16 (.A(mem_rdata[23]),
    .Z(net16));
 BUF_X1 input17 (.A(mem_rdata[24]),
    .Z(net17));
 BUF_X1 input18 (.A(mem_rdata[25]),
    .Z(net18));
 BUF_X1 input19 (.A(mem_rdata[26]),
    .Z(net19));
 BUF_X1 input20 (.A(mem_rdata[27]),
    .Z(net20));
 BUF_X1 input21 (.A(mem_rdata[28]),
    .Z(net21));
 BUF_X1 input22 (.A(mem_rdata[29]),
    .Z(net22));
 BUF_X1 input23 (.A(mem_rdata[2]),
    .Z(net23));
 BUF_X1 input24 (.A(mem_rdata[30]),
    .Z(net24));
 BUF_X1 input25 (.A(mem_rdata[31]),
    .Z(net25));
 BUF_X1 input26 (.A(mem_rdata[3]),
    .Z(net26));
 BUF_X1 input27 (.A(mem_rdata[4]),
    .Z(net27));
 BUF_X1 input28 (.A(mem_rdata[5]),
    .Z(net28));
 BUF_X1 input29 (.A(mem_rdata[6]),
    .Z(net29));
 BUF_X1 input30 (.A(mem_rdata[7]),
    .Z(net30));
 BUF_X1 input31 (.A(mem_rdata[8]),
    .Z(net31));
 BUF_X1 input32 (.A(mem_rdata[9]),
    .Z(net32));
 BUF_X1 output33 (.A(net33),
    .Z(bist_done));
 BUF_X1 output34 (.A(net34),
    .Z(bist_pass));
 BUF_X1 output35 (.A(net35),
    .Z(error_addr[0]));
 BUF_X1 output36 (.A(net36),
    .Z(error_addr[1]));
 BUF_X1 output37 (.A(net37),
    .Z(error_addr[2]));
 BUF_X1 output38 (.A(net38),
    .Z(error_addr[3]));
 BUF_X1 output39 (.A(net39),
    .Z(error_addr[4]));
 BUF_X1 output40 (.A(net40),
    .Z(error_count[0]));
 BUF_X1 output41 (.A(net41),
    .Z(error_count[10]));
 BUF_X1 output42 (.A(net42),
    .Z(error_count[11]));
 BUF_X1 output43 (.A(net43),
    .Z(error_count[12]));
 BUF_X1 output44 (.A(net44),
    .Z(error_count[13]));
 BUF_X1 output45 (.A(net45),
    .Z(error_count[14]));
 BUF_X1 output46 (.A(net46),
    .Z(error_count[15]));
 BUF_X1 output47 (.A(net47),
    .Z(error_count[16]));
 BUF_X1 output48 (.A(net48),
    .Z(error_count[17]));
 BUF_X1 output49 (.A(net49),
    .Z(error_count[18]));
 BUF_X1 output50 (.A(net50),
    .Z(error_count[19]));
 BUF_X1 output51 (.A(net51),
    .Z(error_count[1]));
 BUF_X1 output52 (.A(net52),
    .Z(error_count[20]));
 BUF_X1 output53 (.A(net53),
    .Z(error_count[21]));
 BUF_X1 output54 (.A(net54),
    .Z(error_count[22]));
 BUF_X1 output55 (.A(net55),
    .Z(error_count[23]));
 BUF_X1 output56 (.A(net56),
    .Z(error_count[24]));
 BUF_X1 output57 (.A(net57),
    .Z(error_count[25]));
 BUF_X1 output58 (.A(net58),
    .Z(error_count[26]));
 BUF_X1 output59 (.A(net59),
    .Z(error_count[27]));
 BUF_X1 output60 (.A(net60),
    .Z(error_count[28]));
 BUF_X1 output61 (.A(net61),
    .Z(error_count[29]));
 BUF_X1 output62 (.A(net62),
    .Z(error_count[2]));
 BUF_X1 output63 (.A(net63),
    .Z(error_count[30]));
 BUF_X1 output64 (.A(net64),
    .Z(error_count[31]));
 BUF_X1 output65 (.A(net65),
    .Z(error_count[3]));
 BUF_X1 output66 (.A(net66),
    .Z(error_count[4]));
 BUF_X1 output67 (.A(net67),
    .Z(error_count[5]));
 BUF_X1 output68 (.A(net68),
    .Z(error_count[6]));
 BUF_X1 output69 (.A(net69),
    .Z(error_count[7]));
 BUF_X1 output70 (.A(net70),
    .Z(error_count[8]));
 BUF_X1 output71 (.A(net71),
    .Z(error_count[9]));
 BUF_X1 output72 (.A(net72),
    .Z(mem_addr[0]));
 BUF_X1 output73 (.A(net73),
    .Z(mem_addr[1]));
 BUF_X1 output74 (.A(net74),
    .Z(mem_addr[2]));
 BUF_X1 output75 (.A(net75),
    .Z(mem_addr[3]));
 BUF_X1 output76 (.A(net76),
    .Z(mem_addr[4]));
 BUF_X1 output77 (.A(net77),
    .Z(mem_enable));
 BUF_X1 output78 (.A(net78),
    .Z(mem_wdata[0]));
 BUF_X1 output79 (.A(net79),
    .Z(mem_wdata[10]));
 BUF_X1 output80 (.A(net80),
    .Z(mem_wdata[11]));
 BUF_X1 output81 (.A(net81),
    .Z(mem_wdata[12]));
 BUF_X1 output82 (.A(net82),
    .Z(mem_wdata[13]));
 BUF_X1 output83 (.A(net83),
    .Z(mem_wdata[14]));
 BUF_X1 output84 (.A(net84),
    .Z(mem_wdata[15]));
 BUF_X1 output85 (.A(net85),
    .Z(mem_wdata[16]));
 BUF_X1 output86 (.A(net86),
    .Z(mem_wdata[17]));
 BUF_X1 output87 (.A(net87),
    .Z(mem_wdata[18]));
 BUF_X1 output88 (.A(net88),
    .Z(mem_wdata[19]));
 BUF_X1 output89 (.A(net89),
    .Z(mem_wdata[1]));
 BUF_X1 output90 (.A(net90),
    .Z(mem_wdata[20]));
 BUF_X1 output91 (.A(net91),
    .Z(mem_wdata[21]));
 BUF_X1 output92 (.A(net92),
    .Z(mem_wdata[22]));
 BUF_X1 output93 (.A(net93),
    .Z(mem_wdata[23]));
 BUF_X1 output94 (.A(net94),
    .Z(mem_wdata[24]));
 BUF_X1 output95 (.A(net95),
    .Z(mem_wdata[25]));
 BUF_X1 output96 (.A(net96),
    .Z(mem_wdata[26]));
 BUF_X1 output97 (.A(net97),
    .Z(mem_wdata[27]));
 BUF_X1 output98 (.A(net98),
    .Z(mem_wdata[28]));
 BUF_X1 output99 (.A(net99),
    .Z(mem_wdata[29]));
 BUF_X1 output100 (.A(net100),
    .Z(mem_wdata[2]));
 BUF_X1 output101 (.A(net101),
    .Z(mem_wdata[30]));
 BUF_X1 output102 (.A(net102),
    .Z(mem_wdata[31]));
 BUF_X1 output103 (.A(net103),
    .Z(mem_wdata[3]));
 BUF_X1 output104 (.A(net104),
    .Z(mem_wdata[4]));
 BUF_X1 output105 (.A(net105),
    .Z(mem_wdata[5]));
 BUF_X1 output106 (.A(net106),
    .Z(mem_wdata[6]));
 BUF_X1 output107 (.A(net107),
    .Z(mem_wdata[7]));
 BUF_X1 output108 (.A(net108),
    .Z(mem_wdata[8]));
 BUF_X1 output109 (.A(net109),
    .Z(mem_wdata[9]));
 BUF_X1 output110 (.A(net110),
    .Z(mem_write));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X4 clkload1 (.A(clknet_2_1__leaf_clk));
 INV_X1 clkload2 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_17 ();
 FILLCELL_X2 FILLER_0_25 ();
 FILLCELL_X16 FILLER_0_30 ();
 FILLCELL_X2 FILLER_0_46 ();
 FILLCELL_X2 FILLER_0_51 ();
 FILLCELL_X1 FILLER_0_53 ();
 FILLCELL_X2 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_139 ();
 FILLCELL_X2 FILLER_0_143 ();
 FILLCELL_X1 FILLER_0_145 ();
 FILLCELL_X4 FILLER_0_149 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X32 FILLER_0_157 ();
 FILLCELL_X16 FILLER_0_189 ();
 FILLCELL_X2 FILLER_0_205 ();
 FILLCELL_X1 FILLER_0_207 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X4 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_40 ();
 FILLCELL_X2 FILLER_1_77 ();
 FILLCELL_X2 FILLER_1_117 ();
 FILLCELL_X8 FILLER_1_139 ();
 FILLCELL_X2 FILLER_1_147 ();
 FILLCELL_X1 FILLER_1_149 ();
 FILLCELL_X32 FILLER_1_167 ();
 FILLCELL_X8 FILLER_1_199 ();
 FILLCELL_X1 FILLER_1_207 ();
 FILLCELL_X16 FILLER_2_1 ();
 FILLCELL_X8 FILLER_2_17 ();
 FILLCELL_X2 FILLER_2_47 ();
 FILLCELL_X1 FILLER_2_49 ();
 FILLCELL_X4 FILLER_2_58 ();
 FILLCELL_X2 FILLER_2_62 ();
 FILLCELL_X1 FILLER_2_64 ();
 FILLCELL_X1 FILLER_2_67 ();
 FILLCELL_X4 FILLER_2_73 ();
 FILLCELL_X4 FILLER_2_81 ();
 FILLCELL_X2 FILLER_2_85 ();
 FILLCELL_X1 FILLER_2_87 ();
 FILLCELL_X4 FILLER_2_92 ();
 FILLCELL_X2 FILLER_2_96 ();
 FILLCELL_X8 FILLER_2_104 ();
 FILLCELL_X2 FILLER_2_112 ();
 FILLCELL_X1 FILLER_2_114 ();
 FILLCELL_X8 FILLER_2_123 ();
 FILLCELL_X4 FILLER_2_131 ();
 FILLCELL_X1 FILLER_2_135 ();
 FILLCELL_X4 FILLER_2_156 ();
 FILLCELL_X2 FILLER_2_164 ();
 FILLCELL_X1 FILLER_2_166 ();
 FILLCELL_X2 FILLER_2_195 ();
 FILLCELL_X1 FILLER_2_197 ();
 FILLCELL_X4 FILLER_2_201 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X8 FILLER_3_17 ();
 FILLCELL_X2 FILLER_3_25 ();
 FILLCELL_X4 FILLER_3_29 ();
 FILLCELL_X1 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_42 ();
 FILLCELL_X1 FILLER_3_50 ();
 FILLCELL_X8 FILLER_3_76 ();
 FILLCELL_X1 FILLER_3_84 ();
 FILLCELL_X4 FILLER_3_89 ();
 FILLCELL_X2 FILLER_3_93 ();
 FILLCELL_X16 FILLER_3_116 ();
 FILLCELL_X4 FILLER_3_132 ();
 FILLCELL_X1 FILLER_3_136 ();
 FILLCELL_X4 FILLER_3_151 ();
 FILLCELL_X2 FILLER_3_155 ();
 FILLCELL_X2 FILLER_3_167 ();
 FILLCELL_X1 FILLER_3_179 ();
 FILLCELL_X1 FILLER_3_207 ();
 FILLCELL_X2 FILLER_4_20 ();
 FILLCELL_X1 FILLER_4_22 ();
 FILLCELL_X4 FILLER_4_27 ();
 FILLCELL_X2 FILLER_4_31 ();
 FILLCELL_X1 FILLER_4_59 ();
 FILLCELL_X8 FILLER_4_78 ();
 FILLCELL_X2 FILLER_4_86 ();
 FILLCELL_X1 FILLER_4_95 ();
 FILLCELL_X8 FILLER_4_107 ();
 FILLCELL_X4 FILLER_4_115 ();
 FILLCELL_X1 FILLER_4_119 ();
 FILLCELL_X8 FILLER_4_124 ();
 FILLCELL_X4 FILLER_4_132 ();
 FILLCELL_X2 FILLER_4_136 ();
 FILLCELL_X8 FILLER_4_146 ();
 FILLCELL_X4 FILLER_4_154 ();
 FILLCELL_X2 FILLER_4_162 ();
 FILLCELL_X4 FILLER_4_173 ();
 FILLCELL_X16 FILLER_4_188 ();
 FILLCELL_X4 FILLER_4_204 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X1 FILLER_5_46 ();
 FILLCELL_X2 FILLER_5_86 ();
 FILLCELL_X2 FILLER_5_105 ();
 FILLCELL_X1 FILLER_5_107 ();
 FILLCELL_X4 FILLER_5_115 ();
 FILLCELL_X2 FILLER_5_119 ();
 FILLCELL_X1 FILLER_5_121 ();
 FILLCELL_X2 FILLER_5_139 ();
 FILLCELL_X2 FILLER_5_152 ();
 FILLCELL_X4 FILLER_5_162 ();
 FILLCELL_X2 FILLER_5_166 ();
 FILLCELL_X1 FILLER_5_173 ();
 FILLCELL_X1 FILLER_5_182 ();
 FILLCELL_X2 FILLER_5_193 ();
 FILLCELL_X4 FILLER_5_198 ();
 FILLCELL_X2 FILLER_5_202 ();
 FILLCELL_X1 FILLER_5_207 ();
 FILLCELL_X16 FILLER_6_1 ();
 FILLCELL_X2 FILLER_6_17 ();
 FILLCELL_X1 FILLER_6_49 ();
 FILLCELL_X32 FILLER_6_59 ();
 FILLCELL_X32 FILLER_6_95 ();
 FILLCELL_X4 FILLER_6_127 ();
 FILLCELL_X2 FILLER_6_131 ();
 FILLCELL_X1 FILLER_6_133 ();
 FILLCELL_X4 FILLER_6_141 ();
 FILLCELL_X2 FILLER_6_154 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X4 FILLER_6_177 ();
 FILLCELL_X1 FILLER_6_181 ();
 FILLCELL_X4 FILLER_6_202 ();
 FILLCELL_X2 FILLER_6_206 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_17 ();
 FILLCELL_X2 FILLER_7_21 ();
 FILLCELL_X1 FILLER_7_23 ();
 FILLCELL_X1 FILLER_7_31 ();
 FILLCELL_X1 FILLER_7_42 ();
 FILLCELL_X1 FILLER_7_47 ();
 FILLCELL_X4 FILLER_7_54 ();
 FILLCELL_X1 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_69 ();
 FILLCELL_X2 FILLER_7_73 ();
 FILLCELL_X4 FILLER_7_82 ();
 FILLCELL_X1 FILLER_7_86 ();
 FILLCELL_X1 FILLER_7_104 ();
 FILLCELL_X16 FILLER_7_117 ();
 FILLCELL_X16 FILLER_7_152 ();
 FILLCELL_X4 FILLER_7_168 ();
 FILLCELL_X1 FILLER_7_172 ();
 FILLCELL_X1 FILLER_7_186 ();
 FILLCELL_X8 FILLER_7_190 ();
 FILLCELL_X4 FILLER_7_198 ();
 FILLCELL_X2 FILLER_7_202 ();
 FILLCELL_X1 FILLER_7_204 ();
 FILLCELL_X4 FILLER_8_33 ();
 FILLCELL_X2 FILLER_8_37 ();
 FILLCELL_X1 FILLER_8_83 ();
 FILLCELL_X4 FILLER_8_95 ();
 FILLCELL_X1 FILLER_8_144 ();
 FILLCELL_X1 FILLER_8_149 ();
 FILLCELL_X1 FILLER_8_153 ();
 FILLCELL_X1 FILLER_8_159 ();
 FILLCELL_X4 FILLER_8_165 ();
 FILLCELL_X2 FILLER_8_169 ();
 FILLCELL_X1 FILLER_8_171 ();
 FILLCELL_X1 FILLER_8_179 ();
 FILLCELL_X4 FILLER_9_10 ();
 FILLCELL_X2 FILLER_9_30 ();
 FILLCELL_X1 FILLER_9_32 ();
 FILLCELL_X1 FILLER_9_36 ();
 FILLCELL_X1 FILLER_9_61 ();
 FILLCELL_X1 FILLER_9_66 ();
 FILLCELL_X1 FILLER_9_76 ();
 FILLCELL_X1 FILLER_9_84 ();
 FILLCELL_X4 FILLER_9_89 ();
 FILLCELL_X2 FILLER_9_93 ();
 FILLCELL_X8 FILLER_9_105 ();
 FILLCELL_X4 FILLER_9_117 ();
 FILLCELL_X1 FILLER_9_121 ();
 FILLCELL_X1 FILLER_9_146 ();
 FILLCELL_X8 FILLER_9_171 ();
 FILLCELL_X2 FILLER_9_179 ();
 FILLCELL_X8 FILLER_9_192 ();
 FILLCELL_X2 FILLER_9_200 ();
 FILLCELL_X2 FILLER_10_13 ();
 FILLCELL_X1 FILLER_10_15 ();
 FILLCELL_X8 FILLER_10_19 ();
 FILLCELL_X1 FILLER_10_27 ();
 FILLCELL_X1 FILLER_10_31 ();
 FILLCELL_X2 FILLER_10_50 ();
 FILLCELL_X1 FILLER_10_52 ();
 FILLCELL_X1 FILLER_10_63 ();
 FILLCELL_X1 FILLER_10_71 ();
 FILLCELL_X8 FILLER_10_107 ();
 FILLCELL_X4 FILLER_10_115 ();
 FILLCELL_X2 FILLER_10_119 ();
 FILLCELL_X1 FILLER_10_121 ();
 FILLCELL_X8 FILLER_10_125 ();
 FILLCELL_X2 FILLER_10_133 ();
 FILLCELL_X2 FILLER_10_140 ();
 FILLCELL_X1 FILLER_10_142 ();
 FILLCELL_X16 FILLER_10_146 ();
 FILLCELL_X8 FILLER_10_162 ();
 FILLCELL_X4 FILLER_10_170 ();
 FILLCELL_X1 FILLER_10_174 ();
 FILLCELL_X4 FILLER_11_43 ();
 FILLCELL_X1 FILLER_11_47 ();
 FILLCELL_X1 FILLER_11_52 ();
 FILLCELL_X2 FILLER_11_57 ();
 FILLCELL_X2 FILLER_11_63 ();
 FILLCELL_X1 FILLER_11_80 ();
 FILLCELL_X2 FILLER_11_84 ();
 FILLCELL_X1 FILLER_11_86 ();
 FILLCELL_X16 FILLER_11_109 ();
 FILLCELL_X4 FILLER_11_125 ();
 FILLCELL_X2 FILLER_11_129 ();
 FILLCELL_X2 FILLER_11_143 ();
 FILLCELL_X1 FILLER_11_145 ();
 FILLCELL_X4 FILLER_11_163 ();
 FILLCELL_X1 FILLER_11_167 ();
 FILLCELL_X1 FILLER_11_181 ();
 FILLCELL_X4 FILLER_11_186 ();
 FILLCELL_X2 FILLER_11_190 ();
 FILLCELL_X8 FILLER_11_195 ();
 FILLCELL_X4 FILLER_11_203 ();
 FILLCELL_X1 FILLER_11_207 ();
 FILLCELL_X1 FILLER_12_14 ();
 FILLCELL_X1 FILLER_12_18 ();
 FILLCELL_X2 FILLER_12_26 ();
 FILLCELL_X1 FILLER_12_28 ();
 FILLCELL_X2 FILLER_12_41 ();
 FILLCELL_X1 FILLER_12_43 ();
 FILLCELL_X4 FILLER_12_48 ();
 FILLCELL_X2 FILLER_12_52 ();
 FILLCELL_X4 FILLER_12_89 ();
 FILLCELL_X8 FILLER_12_98 ();
 FILLCELL_X4 FILLER_12_106 ();
 FILLCELL_X2 FILLER_12_110 ();
 FILLCELL_X1 FILLER_12_112 ();
 FILLCELL_X16 FILLER_12_116 ();
 FILLCELL_X4 FILLER_12_132 ();
 FILLCELL_X2 FILLER_12_136 ();
 FILLCELL_X1 FILLER_12_138 ();
 FILLCELL_X2 FILLER_12_174 ();
 FILLCELL_X1 FILLER_12_176 ();
 FILLCELL_X2 FILLER_12_191 ();
 FILLCELL_X8 FILLER_12_196 ();
 FILLCELL_X4 FILLER_12_204 ();
 FILLCELL_X2 FILLER_13_4 ();
 FILLCELL_X1 FILLER_13_6 ();
 FILLCELL_X4 FILLER_13_20 ();
 FILLCELL_X2 FILLER_13_24 ();
 FILLCELL_X4 FILLER_13_28 ();
 FILLCELL_X2 FILLER_13_32 ();
 FILLCELL_X4 FILLER_13_46 ();
 FILLCELL_X1 FILLER_13_57 ();
 FILLCELL_X4 FILLER_13_61 ();
 FILLCELL_X1 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_76 ();
 FILLCELL_X16 FILLER_13_84 ();
 FILLCELL_X8 FILLER_13_100 ();
 FILLCELL_X2 FILLER_13_108 ();
 FILLCELL_X1 FILLER_13_110 ();
 FILLCELL_X1 FILLER_13_119 ();
 FILLCELL_X4 FILLER_13_164 ();
 FILLCELL_X1 FILLER_14_10 ();
 FILLCELL_X2 FILLER_14_19 ();
 FILLCELL_X4 FILLER_14_84 ();
 FILLCELL_X8 FILLER_14_95 ();
 FILLCELL_X1 FILLER_14_103 ();
 FILLCELL_X16 FILLER_14_124 ();
 FILLCELL_X1 FILLER_14_140 ();
 FILLCELL_X1 FILLER_14_146 ();
 FILLCELL_X1 FILLER_14_160 ();
 FILLCELL_X8 FILLER_14_169 ();
 FILLCELL_X8 FILLER_14_184 ();
 FILLCELL_X2 FILLER_14_192 ();
 FILLCELL_X8 FILLER_14_197 ();
 FILLCELL_X2 FILLER_14_205 ();
 FILLCELL_X1 FILLER_14_207 ();
 FILLCELL_X4 FILLER_15_19 ();
 FILLCELL_X1 FILLER_15_39 ();
 FILLCELL_X1 FILLER_15_47 ();
 FILLCELL_X1 FILLER_15_54 ();
 FILLCELL_X1 FILLER_15_84 ();
 FILLCELL_X8 FILLER_15_90 ();
 FILLCELL_X4 FILLER_15_98 ();
 FILLCELL_X1 FILLER_15_102 ();
 FILLCELL_X4 FILLER_15_135 ();
 FILLCELL_X2 FILLER_15_139 ();
 FILLCELL_X1 FILLER_15_141 ();
 FILLCELL_X4 FILLER_15_155 ();
 FILLCELL_X1 FILLER_15_159 ();
 FILLCELL_X8 FILLER_15_164 ();
 FILLCELL_X2 FILLER_15_176 ();
 FILLCELL_X1 FILLER_15_178 ();
 FILLCELL_X8 FILLER_15_192 ();
 FILLCELL_X4 FILLER_15_200 ();
 FILLCELL_X1 FILLER_15_204 ();
 FILLCELL_X16 FILLER_16_19 ();
 FILLCELL_X2 FILLER_16_35 ();
 FILLCELL_X2 FILLER_16_41 ();
 FILLCELL_X2 FILLER_16_56 ();
 FILLCELL_X1 FILLER_16_71 ();
 FILLCELL_X1 FILLER_16_84 ();
 FILLCELL_X8 FILLER_16_94 ();
 FILLCELL_X4 FILLER_16_102 ();
 FILLCELL_X2 FILLER_16_106 ();
 FILLCELL_X1 FILLER_16_108 ();
 FILLCELL_X2 FILLER_16_120 ();
 FILLCELL_X8 FILLER_16_141 ();
 FILLCELL_X2 FILLER_16_205 ();
 FILLCELL_X1 FILLER_16_207 ();
 FILLCELL_X2 FILLER_17_13 ();
 FILLCELL_X16 FILLER_17_21 ();
 FILLCELL_X1 FILLER_17_37 ();
 FILLCELL_X1 FILLER_17_42 ();
 FILLCELL_X2 FILLER_17_56 ();
 FILLCELL_X4 FILLER_17_62 ();
 FILLCELL_X2 FILLER_17_66 ();
 FILLCELL_X8 FILLER_17_90 ();
 FILLCELL_X2 FILLER_17_98 ();
 FILLCELL_X1 FILLER_17_108 ();
 FILLCELL_X4 FILLER_17_113 ();
 FILLCELL_X1 FILLER_17_117 ();
 FILLCELL_X1 FILLER_17_126 ();
 FILLCELL_X32 FILLER_17_149 ();
 FILLCELL_X16 FILLER_17_181 ();
 FILLCELL_X8 FILLER_17_197 ();
 FILLCELL_X2 FILLER_17_205 ();
 FILLCELL_X1 FILLER_17_207 ();
 FILLCELL_X8 FILLER_18_20 ();
 FILLCELL_X2 FILLER_18_28 ();
 FILLCELL_X16 FILLER_18_47 ();
 FILLCELL_X16 FILLER_18_68 ();
 FILLCELL_X2 FILLER_18_84 ();
 FILLCELL_X4 FILLER_18_89 ();
 FILLCELL_X1 FILLER_18_93 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X1 FILLER_18_117 ();
 FILLCELL_X8 FILLER_18_137 ();
 FILLCELL_X4 FILLER_18_145 ();
 FILLCELL_X1 FILLER_18_149 ();
 FILLCELL_X4 FILLER_18_157 ();
 FILLCELL_X4 FILLER_18_194 ();
 FILLCELL_X2 FILLER_18_198 ();
 FILLCELL_X2 FILLER_18_206 ();
 FILLCELL_X1 FILLER_19_1 ();
 FILLCELL_X16 FILLER_19_25 ();
 FILLCELL_X4 FILLER_19_41 ();
 FILLCELL_X2 FILLER_19_45 ();
 FILLCELL_X1 FILLER_19_47 ();
 FILLCELL_X8 FILLER_19_65 ();
 FILLCELL_X4 FILLER_19_73 ();
 FILLCELL_X2 FILLER_19_77 ();
 FILLCELL_X4 FILLER_19_97 ();
 FILLCELL_X16 FILLER_19_110 ();
 FILLCELL_X8 FILLER_19_126 ();
 FILLCELL_X2 FILLER_19_139 ();
 FILLCELL_X1 FILLER_19_149 ();
 FILLCELL_X2 FILLER_19_182 ();
 FILLCELL_X1 FILLER_20_20 ();
 FILLCELL_X32 FILLER_20_26 ();
 FILLCELL_X16 FILLER_20_58 ();
 FILLCELL_X4 FILLER_20_74 ();
 FILLCELL_X2 FILLER_20_98 ();
 FILLCELL_X1 FILLER_20_100 ();
 FILLCELL_X4 FILLER_20_110 ();
 FILLCELL_X8 FILLER_20_119 ();
 FILLCELL_X1 FILLER_20_127 ();
 FILLCELL_X1 FILLER_20_141 ();
 FILLCELL_X4 FILLER_20_147 ();
 FILLCELL_X2 FILLER_20_164 ();
 FILLCELL_X1 FILLER_20_170 ();
 FILLCELL_X2 FILLER_20_179 ();
 FILLCELL_X4 FILLER_20_201 ();
 FILLCELL_X1 FILLER_21_13 ();
 FILLCELL_X32 FILLER_21_17 ();
 FILLCELL_X16 FILLER_21_49 ();
 FILLCELL_X8 FILLER_21_65 ();
 FILLCELL_X4 FILLER_21_73 ();
 FILLCELL_X1 FILLER_21_77 ();
 FILLCELL_X1 FILLER_21_99 ();
 FILLCELL_X1 FILLER_21_103 ();
 FILLCELL_X1 FILLER_21_115 ();
 FILLCELL_X8 FILLER_21_121 ();
 FILLCELL_X2 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_149 ();
 FILLCELL_X2 FILLER_21_166 ();
 FILLCELL_X1 FILLER_21_179 ();
 FILLCELL_X16 FILLER_21_189 ();
 FILLCELL_X2 FILLER_21_205 ();
 FILLCELL_X1 FILLER_21_207 ();
 FILLCELL_X1 FILLER_22_4 ();
 FILLCELL_X1 FILLER_22_11 ();
 FILLCELL_X32 FILLER_22_15 ();
 FILLCELL_X16 FILLER_22_47 ();
 FILLCELL_X8 FILLER_22_63 ();
 FILLCELL_X2 FILLER_22_71 ();
 FILLCELL_X1 FILLER_22_73 ();
 FILLCELL_X2 FILLER_22_94 ();
 FILLCELL_X1 FILLER_22_104 ();
 FILLCELL_X16 FILLER_22_108 ();
 FILLCELL_X4 FILLER_22_124 ();
 FILLCELL_X1 FILLER_22_140 ();
 FILLCELL_X4 FILLER_22_176 ();
 FILLCELL_X2 FILLER_22_180 ();
 FILLCELL_X16 FILLER_22_189 ();
 FILLCELL_X2 FILLER_22_205 ();
 FILLCELL_X1 FILLER_22_207 ();
 FILLCELL_X4 FILLER_23_7 ();
 FILLCELL_X32 FILLER_23_20 ();
 FILLCELL_X8 FILLER_23_52 ();
 FILLCELL_X2 FILLER_23_60 ();
 FILLCELL_X1 FILLER_23_94 ();
 FILLCELL_X2 FILLER_23_99 ();
 FILLCELL_X16 FILLER_23_103 ();
 FILLCELL_X1 FILLER_23_128 ();
 FILLCELL_X1 FILLER_23_138 ();
 FILLCELL_X8 FILLER_23_144 ();
 FILLCELL_X1 FILLER_23_167 ();
 FILLCELL_X4 FILLER_23_177 ();
 FILLCELL_X1 FILLER_23_181 ();
 FILLCELL_X4 FILLER_23_202 ();
 FILLCELL_X2 FILLER_23_206 ();
 FILLCELL_X1 FILLER_24_7 ();
 FILLCELL_X1 FILLER_24_17 ();
 FILLCELL_X32 FILLER_24_21 ();
 FILLCELL_X16 FILLER_24_53 ();
 FILLCELL_X8 FILLER_24_69 ();
 FILLCELL_X1 FILLER_24_77 ();
 FILLCELL_X1 FILLER_24_85 ();
 FILLCELL_X1 FILLER_24_90 ();
 FILLCELL_X1 FILLER_24_94 ();
 FILLCELL_X1 FILLER_24_98 ();
 FILLCELL_X1 FILLER_24_103 ();
 FILLCELL_X2 FILLER_24_108 ();
 FILLCELL_X1 FILLER_24_113 ();
 FILLCELL_X2 FILLER_24_127 ();
 FILLCELL_X1 FILLER_24_129 ();
 FILLCELL_X2 FILLER_24_157 ();
 FILLCELL_X1 FILLER_24_159 ();
 FILLCELL_X1 FILLER_24_168 ();
 FILLCELL_X8 FILLER_24_171 ();
 FILLCELL_X16 FILLER_24_183 ();
 FILLCELL_X8 FILLER_24_199 ();
 FILLCELL_X1 FILLER_24_207 ();
 FILLCELL_X2 FILLER_25_10 ();
 FILLCELL_X4 FILLER_25_21 ();
 FILLCELL_X2 FILLER_25_25 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_65 ();
 FILLCELL_X2 FILLER_25_73 ();
 FILLCELL_X1 FILLER_25_75 ();
 FILLCELL_X4 FILLER_25_81 ();
 FILLCELL_X2 FILLER_25_85 ();
 FILLCELL_X1 FILLER_25_87 ();
 FILLCELL_X8 FILLER_25_93 ();
 FILLCELL_X2 FILLER_25_101 ();
 FILLCELL_X1 FILLER_25_103 ();
 FILLCELL_X1 FILLER_25_112 ();
 FILLCELL_X1 FILLER_25_117 ();
 FILLCELL_X8 FILLER_25_126 ();
 FILLCELL_X1 FILLER_25_139 ();
 FILLCELL_X1 FILLER_25_143 ();
 FILLCELL_X1 FILLER_25_152 ();
 FILLCELL_X2 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_180 ();
 FILLCELL_X8 FILLER_25_196 ();
 FILLCELL_X4 FILLER_25_204 ();
 FILLCELL_X1 FILLER_26_13 ();
 FILLCELL_X1 FILLER_26_79 ();
 FILLCELL_X1 FILLER_26_97 ();
 FILLCELL_X1 FILLER_26_115 ();
 FILLCELL_X1 FILLER_26_133 ();
 FILLCELL_X1 FILLER_26_151 ();
 FILLCELL_X32 FILLER_26_173 ();
 FILLCELL_X2 FILLER_26_205 ();
 FILLCELL_X1 FILLER_26_207 ();
 FILLCELL_X1 FILLER_27_13 ();
 FILLCELL_X8 FILLER_27_68 ();
 FILLCELL_X1 FILLER_27_76 ();
 FILLCELL_X8 FILLER_27_80 ();
 FILLCELL_X4 FILLER_27_88 ();
 FILLCELL_X8 FILLER_27_101 ();
 FILLCELL_X8 FILLER_27_115 ();
 FILLCELL_X4 FILLER_27_123 ();
 FILLCELL_X1 FILLER_27_133 ();
 FILLCELL_X4 FILLER_27_138 ();
 FILLCELL_X2 FILLER_27_142 ();
 FILLCELL_X1 FILLER_27_144 ();
 FILLCELL_X16 FILLER_27_148 ();
 FILLCELL_X2 FILLER_27_164 ();
 FILLCELL_X8 FILLER_27_169 ();
 FILLCELL_X2 FILLER_27_177 ();
 FILLCELL_X1 FILLER_27_179 ();
 FILLCELL_X16 FILLER_27_183 ();
 FILLCELL_X8 FILLER_27_199 ();
 FILLCELL_X1 FILLER_27_207 ();
endmodule
