module parameterized_fft (busy,
    clk,
    data_ready,
    data_valid_in,
    data_valid_out,
    rst_n,
    start,
    data_in_imag,
    data_in_real,
    data_out_imag,
    data_out_real);
 output busy;
 input clk;
 output data_ready;
 input data_valid_in;
 output data_valid_out;
 input rst_n;
 input start;
 input [15:0] data_in_imag;
 input [15:0] data_in_real;
 output [127:0] data_out_imag;
 output [127:0] data_out_real;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire net31;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire net40;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire clknet_leaf_0_clk;
 wire net369;
 wire \bit_rev_idx[0] ;
 wire \bit_rev_idx[1] ;
 wire \bit_rev_idx[2] ;
 wire \butterfly_count[0] ;
 wire \butterfly_count[1] ;
 wire \butterfly_count[2] ;
 wire \butterfly_in_group[0] ;
 wire \butterfly_in_group[1] ;
 wire \butterfly_in_group[2] ;
 wire \group[0] ;
 wire \group[1] ;
 wire \group[2] ;
 wire \idx1[0] ;
 wire \idx1[1] ;
 wire \idx1[2] ;
 wire \idx2[0] ;
 wire \idx2[1] ;
 wire \idx2[2] ;
 wire \sample_count[0] ;
 wire \sample_count[1] ;
 wire \sample_count[2] ;
 wire \samples_imag[0][0] ;
 wire \samples_imag[0][10] ;
 wire \samples_imag[0][11] ;
 wire \samples_imag[0][12] ;
 wire \samples_imag[0][13] ;
 wire \samples_imag[0][14] ;
 wire \samples_imag[0][15] ;
 wire \samples_imag[0][1] ;
 wire \samples_imag[0][2] ;
 wire \samples_imag[0][3] ;
 wire \samples_imag[0][4] ;
 wire \samples_imag[0][5] ;
 wire \samples_imag[0][6] ;
 wire \samples_imag[0][7] ;
 wire \samples_imag[0][8] ;
 wire \samples_imag[0][9] ;
 wire \samples_imag[1][0] ;
 wire \samples_imag[1][10] ;
 wire \samples_imag[1][11] ;
 wire \samples_imag[1][12] ;
 wire \samples_imag[1][13] ;
 wire \samples_imag[1][14] ;
 wire \samples_imag[1][15] ;
 wire \samples_imag[1][1] ;
 wire \samples_imag[1][2] ;
 wire \samples_imag[1][3] ;
 wire \samples_imag[1][4] ;
 wire \samples_imag[1][5] ;
 wire \samples_imag[1][6] ;
 wire \samples_imag[1][7] ;
 wire \samples_imag[1][8] ;
 wire \samples_imag[1][9] ;
 wire \samples_imag[2][0] ;
 wire \samples_imag[2][10] ;
 wire \samples_imag[2][11] ;
 wire \samples_imag[2][12] ;
 wire \samples_imag[2][13] ;
 wire \samples_imag[2][14] ;
 wire \samples_imag[2][15] ;
 wire \samples_imag[2][1] ;
 wire \samples_imag[2][2] ;
 wire \samples_imag[2][3] ;
 wire \samples_imag[2][4] ;
 wire \samples_imag[2][5] ;
 wire \samples_imag[2][6] ;
 wire \samples_imag[2][7] ;
 wire \samples_imag[2][8] ;
 wire \samples_imag[2][9] ;
 wire \samples_imag[3][0] ;
 wire \samples_imag[3][10] ;
 wire \samples_imag[3][11] ;
 wire \samples_imag[3][12] ;
 wire \samples_imag[3][13] ;
 wire \samples_imag[3][14] ;
 wire \samples_imag[3][15] ;
 wire \samples_imag[3][1] ;
 wire \samples_imag[3][2] ;
 wire \samples_imag[3][3] ;
 wire \samples_imag[3][4] ;
 wire \samples_imag[3][5] ;
 wire \samples_imag[3][6] ;
 wire \samples_imag[3][7] ;
 wire \samples_imag[3][8] ;
 wire \samples_imag[3][9] ;
 wire \samples_imag[4][0] ;
 wire \samples_imag[4][10] ;
 wire \samples_imag[4][11] ;
 wire \samples_imag[4][12] ;
 wire \samples_imag[4][13] ;
 wire \samples_imag[4][14] ;
 wire \samples_imag[4][15] ;
 wire \samples_imag[4][1] ;
 wire \samples_imag[4][2] ;
 wire \samples_imag[4][3] ;
 wire \samples_imag[4][4] ;
 wire \samples_imag[4][5] ;
 wire \samples_imag[4][6] ;
 wire \samples_imag[4][7] ;
 wire \samples_imag[4][8] ;
 wire \samples_imag[4][9] ;
 wire \samples_imag[5][0] ;
 wire \samples_imag[5][10] ;
 wire \samples_imag[5][11] ;
 wire \samples_imag[5][12] ;
 wire \samples_imag[5][13] ;
 wire \samples_imag[5][14] ;
 wire \samples_imag[5][15] ;
 wire \samples_imag[5][1] ;
 wire \samples_imag[5][2] ;
 wire \samples_imag[5][3] ;
 wire \samples_imag[5][4] ;
 wire \samples_imag[5][5] ;
 wire \samples_imag[5][6] ;
 wire \samples_imag[5][7] ;
 wire \samples_imag[5][8] ;
 wire \samples_imag[5][9] ;
 wire \samples_imag[6][0] ;
 wire \samples_imag[6][10] ;
 wire \samples_imag[6][11] ;
 wire \samples_imag[6][12] ;
 wire \samples_imag[6][13] ;
 wire \samples_imag[6][14] ;
 wire \samples_imag[6][15] ;
 wire \samples_imag[6][1] ;
 wire \samples_imag[6][2] ;
 wire \samples_imag[6][3] ;
 wire \samples_imag[6][4] ;
 wire \samples_imag[6][5] ;
 wire \samples_imag[6][6] ;
 wire \samples_imag[6][7] ;
 wire \samples_imag[6][8] ;
 wire \samples_imag[6][9] ;
 wire \samples_imag[7][0] ;
 wire \samples_imag[7][10] ;
 wire \samples_imag[7][11] ;
 wire \samples_imag[7][12] ;
 wire \samples_imag[7][13] ;
 wire \samples_imag[7][14] ;
 wire \samples_imag[7][15] ;
 wire \samples_imag[7][1] ;
 wire \samples_imag[7][2] ;
 wire \samples_imag[7][3] ;
 wire \samples_imag[7][4] ;
 wire \samples_imag[7][5] ;
 wire \samples_imag[7][6] ;
 wire \samples_imag[7][7] ;
 wire \samples_imag[7][8] ;
 wire \samples_imag[7][9] ;
 wire \samples_real[0][0] ;
 wire \samples_real[0][10] ;
 wire \samples_real[0][11] ;
 wire \samples_real[0][12] ;
 wire \samples_real[0][13] ;
 wire \samples_real[0][14] ;
 wire \samples_real[0][15] ;
 wire \samples_real[0][1] ;
 wire \samples_real[0][2] ;
 wire \samples_real[0][3] ;
 wire \samples_real[0][4] ;
 wire \samples_real[0][5] ;
 wire \samples_real[0][6] ;
 wire \samples_real[0][7] ;
 wire \samples_real[0][8] ;
 wire \samples_real[0][9] ;
 wire \samples_real[1][0] ;
 wire \samples_real[1][10] ;
 wire \samples_real[1][11] ;
 wire \samples_real[1][12] ;
 wire \samples_real[1][13] ;
 wire \samples_real[1][14] ;
 wire \samples_real[1][15] ;
 wire \samples_real[1][1] ;
 wire \samples_real[1][2] ;
 wire \samples_real[1][3] ;
 wire \samples_real[1][4] ;
 wire \samples_real[1][5] ;
 wire \samples_real[1][6] ;
 wire \samples_real[1][7] ;
 wire \samples_real[1][8] ;
 wire \samples_real[1][9] ;
 wire \samples_real[2][0] ;
 wire \samples_real[2][10] ;
 wire \samples_real[2][11] ;
 wire \samples_real[2][12] ;
 wire \samples_real[2][13] ;
 wire \samples_real[2][14] ;
 wire \samples_real[2][15] ;
 wire \samples_real[2][1] ;
 wire \samples_real[2][2] ;
 wire \samples_real[2][3] ;
 wire \samples_real[2][4] ;
 wire \samples_real[2][5] ;
 wire \samples_real[2][6] ;
 wire \samples_real[2][7] ;
 wire \samples_real[2][8] ;
 wire \samples_real[2][9] ;
 wire \samples_real[3][0] ;
 wire \samples_real[3][10] ;
 wire \samples_real[3][11] ;
 wire \samples_real[3][12] ;
 wire \samples_real[3][13] ;
 wire \samples_real[3][14] ;
 wire \samples_real[3][15] ;
 wire \samples_real[3][1] ;
 wire \samples_real[3][2] ;
 wire \samples_real[3][3] ;
 wire \samples_real[3][4] ;
 wire \samples_real[3][5] ;
 wire \samples_real[3][6] ;
 wire \samples_real[3][7] ;
 wire \samples_real[3][8] ;
 wire \samples_real[3][9] ;
 wire \samples_real[4][0] ;
 wire \samples_real[4][10] ;
 wire \samples_real[4][11] ;
 wire \samples_real[4][12] ;
 wire \samples_real[4][13] ;
 wire \samples_real[4][14] ;
 wire \samples_real[4][15] ;
 wire \samples_real[4][1] ;
 wire \samples_real[4][2] ;
 wire \samples_real[4][3] ;
 wire \samples_real[4][4] ;
 wire \samples_real[4][5] ;
 wire \samples_real[4][6] ;
 wire \samples_real[4][7] ;
 wire \samples_real[4][8] ;
 wire \samples_real[4][9] ;
 wire \samples_real[5][0] ;
 wire \samples_real[5][10] ;
 wire \samples_real[5][11] ;
 wire \samples_real[5][12] ;
 wire \samples_real[5][13] ;
 wire \samples_real[5][14] ;
 wire \samples_real[5][15] ;
 wire \samples_real[5][1] ;
 wire \samples_real[5][2] ;
 wire \samples_real[5][3] ;
 wire \samples_real[5][4] ;
 wire \samples_real[5][5] ;
 wire \samples_real[5][6] ;
 wire \samples_real[5][7] ;
 wire \samples_real[5][8] ;
 wire \samples_real[5][9] ;
 wire \samples_real[6][0] ;
 wire \samples_real[6][10] ;
 wire \samples_real[6][11] ;
 wire \samples_real[6][12] ;
 wire \samples_real[6][13] ;
 wire \samples_real[6][14] ;
 wire \samples_real[6][15] ;
 wire \samples_real[6][1] ;
 wire \samples_real[6][2] ;
 wire \samples_real[6][3] ;
 wire \samples_real[6][4] ;
 wire \samples_real[6][5] ;
 wire \samples_real[6][6] ;
 wire \samples_real[6][7] ;
 wire \samples_real[6][8] ;
 wire \samples_real[6][9] ;
 wire \samples_real[7][0] ;
 wire \samples_real[7][10] ;
 wire \samples_real[7][11] ;
 wire \samples_real[7][12] ;
 wire \samples_real[7][13] ;
 wire \samples_real[7][14] ;
 wire \samples_real[7][15] ;
 wire \samples_real[7][1] ;
 wire \samples_real[7][2] ;
 wire \samples_real[7][3] ;
 wire \samples_real[7][4] ;
 wire \samples_real[7][5] ;
 wire \samples_real[7][6] ;
 wire \samples_real[7][7] ;
 wire \samples_real[7][8] ;
 wire \samples_real[7][9] ;
 wire \stage[0] ;
 wire \stage[1] ;
 wire \stage[2] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \temp_imag[0] ;
 wire \temp_real[0] ;
 wire \twiddle_idx[0] ;
 wire \twiddle_idx[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net394;
 wire net395;
 wire net396;
 wire net385;
 wire net391;
 wire net392;
 wire net393;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;

 gf180mcu_fd_sc_mcu9t5v0__buf_12 _08311_ (.I(\state[3] ),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08312_ (.I(_00563_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _08313_ (.I(net82),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08314_ (.A1(\state[0] ),
    .A2(_00565_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08315_ (.A1(_00564_),
    .A2(_00566_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _08316_ (.I(\stage[2] ),
    .ZN(_07787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08317_ (.A1(_07775_),
    .A2(_07787_),
    .ZN(_07076_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08318_ (.I(\stage[2] ),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08319_ (.A1(_00567_),
    .A2(_07779_),
    .ZN(_07136_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _08320_ (.I(_07136_),
    .ZN(_07664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08321_ (.A1(_00567_),
    .A2(_07781_),
    .ZN(_07123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08322_ (.I(_07123_),
    .ZN(_07668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08323_ (.A1(_00567_),
    .A2(_07775_),
    .ZN(_07103_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _08324_ (.I(_07103_),
    .ZN(_07672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08325_ (.A1(_07787_),
    .A2(_07779_),
    .Z(_07680_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08326_ (.A1(_07787_),
    .A2(_07781_),
    .Z(_05877_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08327_ (.I(_07794_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08328_ (.I(_00568_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08329_ (.I(_00569_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08330_ (.I(_00570_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08331_ (.I(_00571_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08332_ (.I(_00572_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08333_ (.I(_00573_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08334_ (.I(_00574_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08335_ (.I(_00575_),
    .Z(_07177_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08336_ (.A1(_07775_),
    .A2(_07781_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _08337_ (.I(_07794_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08338_ (.A1(_07779_),
    .A2(_07791_),
    .A3(_00577_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08339_ (.A1(_00567_),
    .A2(_00576_),
    .B(_00578_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08340_ (.I(_00579_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _08341_ (.I(\butterfly_count[2] ),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _08342_ (.I(_07660_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _08343_ (.I(_00582_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08344_ (.A1(_07779_),
    .A2(_07781_),
    .B(\stage[2] ),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08345_ (.A1(_00581_),
    .A2(_00584_),
    .A3(_07769_),
    .A4(_00583_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08346_ (.A1(_07672_),
    .A2(_07676_),
    .A3(_07680_),
    .A4(_00585_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08347_ (.A1(_07775_),
    .A2(_07781_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08348_ (.A1(_00567_),
    .A2(_00587_),
    .B(_07078_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08349_ (.A1(_00586_),
    .A2(_00580_),
    .B(_00588_),
    .ZN(_07079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08350_ (.I(net1),
    .ZN(_07637_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _08351_ (.I(_07080_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08352_ (.I(_07775_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08353_ (.A1(_00567_),
    .A2(_00589_),
    .A3(_00590_),
    .A4(_00578_),
    .ZN(_07086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08354_ (.A1(_00581_),
    .A2(_07769_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08355_ (.A1(_07260_),
    .A2(_07252_),
    .A3(_07255_),
    .A4(_07258_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08356_ (.A1(_07243_),
    .A2(_07246_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08357_ (.A1(_07249_),
    .A2(_00591_),
    .A3(_00592_),
    .A4(_00593_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08358_ (.I(_07158_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08359_ (.A1(_07162_),
    .A2(_07164_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08360_ (.A1(_07161_),
    .A2(_00596_),
    .B(_07159_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08361_ (.A1(_00597_),
    .A2(_00595_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08362_ (.A1(_07176_),
    .A2(_07175_),
    .B(_07174_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08363_ (.A1(_07170_),
    .A2(_07173_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08364_ (.A1(_07170_),
    .A2(_07171_),
    .B(_07168_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08365_ (.A1(_00599_),
    .A2(_00600_),
    .B(_00601_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08366_ (.A1(_07162_),
    .A2(_07159_),
    .A3(_07165_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08367_ (.A1(_00602_),
    .A2(_07167_),
    .B(_00603_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08368_ (.A1(_00604_),
    .A2(_00598_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08369_ (.A1(_00581_),
    .A2(_00582_),
    .A3(_07769_),
    .A4(_00584_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08370_ (.A1(_07117_),
    .A2(_07106_),
    .A3(_07109_),
    .A4(_07112_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08371_ (.A1(_07115_),
    .A2(_00607_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08372_ (.I(_07108_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08373_ (.A1(_07112_),
    .A2(_07111_),
    .B(_07109_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08374_ (.A1(_07117_),
    .A2(_07116_),
    .B(_07115_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08375_ (.A1(_07108_),
    .A2(_07111_),
    .A3(_07114_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08376_ (.A1(_00609_),
    .A2(_00610_),
    .B1(_00611_),
    .B2(_00612_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08377_ (.A1(_07106_),
    .A2(_00568_),
    .A3(_00584_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08378_ (.A1(_07105_),
    .A2(_00569_),
    .A3(_00584_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08379_ (.A1(_00608_),
    .A2(_00606_),
    .B1(_00613_),
    .B2(_00614_),
    .C(_00615_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08380_ (.A1(_07122_),
    .A2(_07121_),
    .B(_07135_),
    .C(_07120_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08381_ (.A1(_07135_),
    .A2(_07119_),
    .B(_07134_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08382_ (.A1(_00617_),
    .A2(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08383_ (.A1(\stage[2] ),
    .A2(_07779_),
    .B(_07794_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08384_ (.A1(_07126_),
    .A2(_07129_),
    .A3(_07132_),
    .A4(_00620_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08385_ (.A1(_07126_),
    .A2(_07131_),
    .A3(_07129_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08386_ (.A1(_00620_),
    .A2(_00622_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08387_ (.A1(_07126_),
    .A2(_07128_),
    .B(_07125_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08388_ (.A1(_00577_),
    .A2(_07664_),
    .A3(_00624_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08389_ (.A1(_00619_),
    .A2(_00621_),
    .B(_00625_),
    .C(_00623_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08390_ (.A1(net26),
    .A2(_07779_),
    .A3(_07781_),
    .A4(_00577_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08391_ (.A1(_00567_),
    .A2(_00577_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08392_ (.A1(_07090_),
    .A2(_07089_),
    .B(_07085_),
    .C(_07088_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08393_ (.A1(_07085_),
    .A2(_07087_),
    .B(_07084_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08394_ (.A1(_07676_),
    .A2(_07090_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08395_ (.A1(_00627_),
    .A2(_00628_),
    .B1(_00629_),
    .B2(_00630_),
    .C(_00631_),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08396_ (.A1(_07775_),
    .A2(_07779_),
    .A3(_07781_),
    .B(\stage[2] ),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08397_ (.A1(_07102_),
    .A2(_07101_),
    .B(_07100_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08398_ (.A1(_07102_),
    .A2(_07100_),
    .A3(_07101_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08399_ (.A1(_00569_),
    .A2(_00632_),
    .A3(_00633_),
    .A4(_00634_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08400_ (.A1(_07093_),
    .A2(_07096_),
    .A3(_07099_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08401_ (.A1(_07093_),
    .A2(_07097_),
    .A3(_07096_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08402_ (.A1(_07093_),
    .A2(_07094_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08403_ (.A1(_00633_),
    .A2(_00636_),
    .B(_00638_),
    .C(_00637_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08404_ (.I0(_07098_),
    .I1(_00635_),
    .S(_00639_),
    .Z(_07110_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08405_ (.A1(net5),
    .A2(_07110_),
    .A3(_00626_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08406_ (.A1(_00617_),
    .A2(_00618_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08407_ (.A1(_07126_),
    .A2(_07129_),
    .A3(_07132_),
    .A4(_00620_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08408_ (.A1(_07126_),
    .A2(_07128_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08409_ (.A1(_07125_),
    .A2(_00643_),
    .A3(_00622_),
    .B(_00620_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08410_ (.A1(_00641_),
    .A2(_00642_),
    .B(_00644_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08411_ (.I(_07114_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08412_ (.A1(_00646_),
    .A2(_00611_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08413_ (.A1(_07112_),
    .A2(_00647_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08414_ (.A1(net5),
    .A2(_00645_),
    .A3(_00648_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _08415_ (.I(_07138_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08416_ (.A1(_07142_),
    .A2(_07145_),
    .A3(_07148_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08417_ (.A1(_07156_),
    .A2(_07139_),
    .A3(_07151_),
    .A4(_07154_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08418_ (.A1(_00581_),
    .A2(_00583_),
    .A3(_07769_),
    .A4(_00652_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08419_ (.A1(_00650_),
    .A2(net36),
    .B1(_00651_),
    .B2(_00653_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08420_ (.I(_07139_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08421_ (.A1(_07142_),
    .A2(_07147_),
    .A3(_07145_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08422_ (.A1(_07142_),
    .A2(_07144_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08423_ (.A1(_07141_),
    .A2(_00656_),
    .A3(_00657_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08424_ (.A1(_00577_),
    .A2(_00651_),
    .A3(_00655_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08425_ (.A1(_07156_),
    .A2(_07155_),
    .B(_07154_),
    .C(_07151_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08426_ (.A1(_07151_),
    .A2(_07153_),
    .B(_07150_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08427_ (.A1(_00660_),
    .A2(_00661_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _08428_ (.A1(_00658_),
    .A2(net36),
    .A3(_00655_),
    .B1(_00659_),
    .B2(_00662_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08429_ (.I(_07132_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08430_ (.A1(_00617_),
    .A2(_00618_),
    .B(_00664_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08431_ (.A1(_00664_),
    .A2(_00617_),
    .A3(_00618_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08432_ (.A1(_00665_),
    .A2(_00644_),
    .A3(_00666_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08433_ (.A1(_00654_),
    .A2(_00663_),
    .A3(_00667_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08434_ (.A1(_00640_),
    .A2(_00649_),
    .A3(_00668_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08435_ (.A1(_00663_),
    .A2(_00654_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08436_ (.I(_07148_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08437_ (.A1(_00660_),
    .A2(_00661_),
    .B(_00671_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08438_ (.A1(_07147_),
    .A2(_00672_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08439_ (.A1(_07145_),
    .A2(_00673_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08440_ (.A1(_00674_),
    .A2(_00670_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08441_ (.A1(_00669_),
    .A2(_00675_),
    .ZN(_07160_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08442_ (.A1(_00660_),
    .A2(_00661_),
    .B(_00651_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08443_ (.A1(_07141_),
    .A2(_00656_),
    .A3(_00657_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08444_ (.A1(_00676_),
    .A2(_00677_),
    .B(_07139_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08445_ (.A1(_07122_),
    .A2(_07121_),
    .B(_07120_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08446_ (.A1(_07119_),
    .A2(_07134_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08447_ (.A1(_07135_),
    .A2(_07134_),
    .B(_07129_),
    .C(_07132_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08448_ (.A1(_00679_),
    .A2(_00680_),
    .B(_00681_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08449_ (.A1(_07129_),
    .A2(_07131_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08450_ (.A1(_07128_),
    .A2(_00683_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08451_ (.A1(_07126_),
    .A2(_00682_),
    .A3(_00684_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08452_ (.A1(_00682_),
    .A2(_00684_),
    .B(_07126_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08453_ (.A1(_07125_),
    .A2(_00620_),
    .A3(_00685_),
    .A4(_00686_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08454_ (.A1(_00651_),
    .A2(_00653_),
    .B(_00650_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08455_ (.A1(_07139_),
    .A2(_00676_),
    .A3(_00677_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08456_ (.A1(_00689_),
    .A2(_00688_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08457_ (.A1(_00687_),
    .A2(_00688_),
    .B(_00690_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08458_ (.A1(_00570_),
    .A2(_00678_),
    .A3(_00691_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _08459_ (.I(_00616_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08460_ (.A1(_00569_),
    .A2(_00632_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08461_ (.A1(_00639_),
    .A2(_00694_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08462_ (.A1(_00567_),
    .A2(_07080_),
    .A3(_00590_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08463_ (.A1(_00579_),
    .A2(_00696_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _08464_ (.I(_07081_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08465_ (.A1(_00698_),
    .A2(_00589_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08466_ (.A1(_07077_),
    .A2(_07080_),
    .A3(_00698_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08467_ (.A1(_07077_),
    .A2(_00698_),
    .B1(_00588_),
    .B2(_00699_),
    .C(_00700_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08468_ (.A1(_00588_),
    .A2(_00579_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08469_ (.A1(_07676_),
    .A2(_07672_),
    .A3(_07680_),
    .A4(_00585_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _08470_ (.I(_07676_),
    .ZN(_07091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08471_ (.A1(_00569_),
    .A2(_00632_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08472_ (.A1(_00630_),
    .A2(_00629_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08473_ (.A1(_07088_),
    .A2(_07085_),
    .A3(_07090_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08474_ (.A1(_07103_),
    .A2(_00706_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08475_ (.A1(_00705_),
    .A2(_00704_),
    .B1(_00585_),
    .B2(_00707_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _08476_ (.A1(_00697_),
    .A2(_00701_),
    .B1(_00702_),
    .B2(_00703_),
    .C1(_07091_),
    .C2(_00708_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08477_ (.A1(_07090_),
    .A2(_07089_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08478_ (.A1(_07088_),
    .A2(_00710_),
    .B(_07087_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08479_ (.A1(_07085_),
    .A2(_00711_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08480_ (.A1(_07091_),
    .A2(_00708_),
    .A3(_00712_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08481_ (.I(_07099_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08482_ (.I(_07097_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08483_ (.A1(_00714_),
    .A2(_00633_),
    .B(_00715_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08484_ (.A1(_07096_),
    .A2(_00716_),
    .B(_07094_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08485_ (.A1(_07094_),
    .A2(_07096_),
    .A3(_00716_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08486_ (.A1(_07093_),
    .A2(_00694_),
    .A3(_00717_),
    .A4(_00718_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08487_ (.A1(_00713_),
    .A2(_00709_),
    .A3(_00695_),
    .B(_00719_),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08488_ (.A1(_00569_),
    .A2(_00678_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08489_ (.A1(_07106_),
    .A2(_00613_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08490_ (.A1(net5),
    .A2(_00721_),
    .B(_00626_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08491_ (.A1(_00688_),
    .A2(_00720_),
    .A3(_00722_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08492_ (.A1(_00693_),
    .A2(_07104_),
    .B(_00723_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08493_ (.A1(_00605_),
    .A2(_07160_),
    .A3(_00692_),
    .A4(_00724_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08494_ (.I(_07164_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08495_ (.A1(_00602_),
    .A2(_07167_),
    .B(_07165_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08496_ (.I(_07162_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08497_ (.A1(_00727_),
    .A2(_00726_),
    .B(_00728_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08498_ (.A1(_00727_),
    .A2(_00726_),
    .A3(_00728_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08499_ (.A1(_00729_),
    .A2(_00730_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08500_ (.A1(net36),
    .A2(_00731_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08501_ (.A1(_07159_),
    .A2(_07161_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08502_ (.A1(_07158_),
    .A2(_00733_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08503_ (.A1(_00729_),
    .A2(_00730_),
    .A3(_07660_),
    .A4(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08504_ (.A1(_00654_),
    .A2(_00663_),
    .A3(_00645_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08505_ (.A1(_00693_),
    .A2(_00736_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08506_ (.A1(_07106_),
    .A2(_00613_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08507_ (.A1(net5),
    .A2(_00738_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08508_ (.A1(_00569_),
    .A2(_00678_),
    .A3(_00689_),
    .A4(_00688_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08509_ (.A1(_00670_),
    .A2(_00687_),
    .B1(_00739_),
    .B2(_00736_),
    .C(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08510_ (.A1(_07104_),
    .A2(_00737_),
    .B(_00741_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08511_ (.I0(_00732_),
    .I1(_00735_),
    .S(_00742_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08512_ (.I(_07182_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08513_ (.I(_07186_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08514_ (.A1(_07191_),
    .A2(_07189_),
    .B(_07188_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08515_ (.I(_07185_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08516_ (.A1(_00746_),
    .A2(_00745_),
    .B(_00747_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08517_ (.A1(_07183_),
    .A2(_00748_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08518_ (.I(_07197_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08519_ (.A1(_07200_),
    .A2(_07199_),
    .B(_07198_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08520_ (.I(_07195_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08521_ (.A1(_00750_),
    .A2(_00751_),
    .B(_00752_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08522_ (.A1(_07183_),
    .A2(_07186_),
    .A3(_07189_),
    .A4(_07192_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08523_ (.A1(_07194_),
    .A2(_00753_),
    .B(_00754_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08524_ (.A1(_00744_),
    .A2(_00749_),
    .A3(_00755_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08525_ (.A1(_07180_),
    .A2(_00756_),
    .B(_07179_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08526_ (.A1(net18),
    .A2(_00569_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08527_ (.A1(_00598_),
    .A2(_00604_),
    .A3(_00758_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08528_ (.A1(_00598_),
    .A2(_00604_),
    .B(net18),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08529_ (.A1(_00759_),
    .A2(_00760_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08530_ (.A1(_00757_),
    .A2(_00761_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08531_ (.A1(_07186_),
    .A2(_07189_),
    .A3(_07192_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08532_ (.A1(_07194_),
    .A2(_00753_),
    .B(_00763_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08533_ (.A1(_00748_),
    .A2(_07182_),
    .A3(_07179_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08534_ (.A1(_07179_),
    .A2(_07183_),
    .A3(_07182_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08535_ (.A1(_07179_),
    .A2(_07180_),
    .B(_00766_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08536_ (.A1(_00765_),
    .A2(_00764_),
    .B(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08537_ (.A1(_00569_),
    .A2(_00678_),
    .A3(_00689_),
    .A4(_00688_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08538_ (.A1(_00769_),
    .A2(_00768_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08539_ (.A1(_00670_),
    .A2(_00687_),
    .B1(_00739_),
    .B2(_00736_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08540_ (.A1(_07104_),
    .A2(_00737_),
    .B(_00771_),
    .C(_00770_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08541_ (.A1(_00762_),
    .A2(_00772_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08542_ (.I(_07660_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08543_ (.A1(_00725_),
    .A2(_00743_),
    .B(_00773_),
    .C(_00774_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08544_ (.A1(_07183_),
    .A2(_00748_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08545_ (.A1(_00764_),
    .A2(_00776_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08546_ (.A1(_00749_),
    .A2(_00755_),
    .A3(_00777_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08547_ (.I(_07211_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08548_ (.I(_07217_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08549_ (.A1(_07220_),
    .A2(_07219_),
    .B(_07218_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _08550_ (.I(_07215_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08551_ (.A1(_00780_),
    .A2(_00781_),
    .B(_00782_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08552_ (.A1(_07214_),
    .A2(_00783_),
    .B(_07212_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08553_ (.A1(_07209_),
    .A2(_07206_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08554_ (.A1(_00779_),
    .A2(_00784_),
    .B(_00785_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08555_ (.A1(_07206_),
    .A2(_07208_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08556_ (.A1(_07205_),
    .A2(_00786_),
    .A3(_07202_),
    .A4(_00787_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08557_ (.I(_07203_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08558_ (.I(_07202_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08559_ (.A1(_00789_),
    .A2(_00790_),
    .B(_00569_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08560_ (.A1(_00791_),
    .A2(_00788_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _08561_ (.I(_00583_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08562_ (.A1(_00757_),
    .A2(_00778_),
    .B1(_00792_),
    .B2(_00793_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08563_ (.A1(net18),
    .A2(_00734_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08564_ (.A1(_00729_),
    .A2(_00730_),
    .A3(_00795_),
    .B1(_00760_),
    .B2(_00759_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08565_ (.A1(_00778_),
    .A2(_00761_),
    .B1(_00796_),
    .B2(_00768_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08566_ (.A1(_00640_),
    .A2(_00649_),
    .A3(_00668_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08567_ (.A1(_00670_),
    .A2(_00674_),
    .B(net18),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08568_ (.A1(_00798_),
    .A2(_00799_),
    .B(_00768_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08569_ (.I0(_00797_),
    .I1(_00800_),
    .S(_00742_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08570_ (.A1(_00762_),
    .A2(_00772_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08571_ (.I(_00778_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08572_ (.A1(_07205_),
    .A2(_00786_),
    .A3(_00787_),
    .B(_07203_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08573_ (.I(net36),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08574_ (.A1(_00790_),
    .A2(_00804_),
    .B(_00805_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08575_ (.A1(_00803_),
    .A2(_00806_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08576_ (.A1(_00794_),
    .A2(_00801_),
    .B1(net33),
    .B2(_00807_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08577_ (.A1(_00605_),
    .A2(_07160_),
    .A3(_00692_),
    .A4(_00724_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08578_ (.A1(net36),
    .A2(_00731_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08579_ (.A1(_00583_),
    .A2(_00669_),
    .A3(_00675_),
    .B(_00735_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _08580_ (.I0(_00810_),
    .I1(_00811_),
    .S(_00742_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08581_ (.A1(_00742_),
    .A2(_00731_),
    .A3(_00795_),
    .B(_00806_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08582_ (.A1(_00813_),
    .A2(_00773_),
    .A3(_00812_),
    .A4(_00809_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08583_ (.A1(_00775_),
    .A2(_00808_),
    .A3(_00814_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08584_ (.I(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08585_ (.A1(_07161_),
    .A2(_00729_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08586_ (.A1(_07159_),
    .A2(_00805_),
    .A3(_00742_),
    .A4(_00817_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08587_ (.A1(_00629_),
    .A2(_00630_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08588_ (.A1(_07103_),
    .A2(_00706_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08589_ (.A1(_00694_),
    .A2(_00819_),
    .B1(_00606_),
    .B2(_00820_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08590_ (.A1(_07088_),
    .A2(_00710_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08591_ (.A1(_07091_),
    .A2(_07103_),
    .A3(_00706_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08592_ (.A1(_00585_),
    .A2(_00823_),
    .B(_07086_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08593_ (.A1(_07091_),
    .A2(_00694_),
    .A3(_00819_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _08594_ (.A1(_00821_),
    .A2(_07676_),
    .A3(_00822_),
    .B1(_00824_),
    .B2(_00825_),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08595_ (.A1(_00694_),
    .A2(_00639_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08596_ (.A1(_00616_),
    .A2(_00826_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08597_ (.A1(_07111_),
    .A2(_07114_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08598_ (.A1(_07112_),
    .A2(_07111_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08599_ (.A1(_00611_),
    .A2(_00828_),
    .B(_00829_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08600_ (.A1(_07109_),
    .A2(_00830_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08601_ (.A1(_07094_),
    .A2(_07096_),
    .B(_07093_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08602_ (.A1(_00715_),
    .A2(_00714_),
    .A3(_00633_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _08603_ (.A1(_00704_),
    .A2(_00716_),
    .A3(_00832_),
    .A4(_00833_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08604_ (.I0(_00831_),
    .I1(_00834_),
    .S(_00616_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08605_ (.A1(_07095_),
    .A2(_00827_),
    .B(_00835_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08606_ (.A1(_07129_),
    .A2(_07131_),
    .A3(_00665_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08607_ (.A1(_07131_),
    .A2(_00665_),
    .B(_07129_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08608_ (.A1(_00625_),
    .A2(_00837_),
    .A3(_00838_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08609_ (.I(_07142_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08610_ (.A1(_00840_),
    .A2(_07144_),
    .A3(_07147_),
    .A4(_00672_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08611_ (.A1(_00840_),
    .A2(_07145_),
    .A3(_00672_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08612_ (.A1(_00840_),
    .A2(_07145_),
    .A3(_07147_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08613_ (.A1(_00840_),
    .A2(_07145_),
    .A3(_07144_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08614_ (.A1(_00840_),
    .A2(_07144_),
    .B(_00843_),
    .C(_00844_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08615_ (.A1(_00841_),
    .A2(_00842_),
    .A3(_00845_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08616_ (.I0(_00839_),
    .I1(_00846_),
    .S(_00670_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08617_ (.A1(_00736_),
    .A2(_00836_),
    .B(_00847_),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08618_ (.A1(_07159_),
    .A2(_07162_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08619_ (.A1(_00726_),
    .A2(_00727_),
    .B(_00848_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08620_ (.A1(_00733_),
    .A2(_00849_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08621_ (.I(_00742_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08622_ (.A1(_07158_),
    .A2(_07157_),
    .A3(_00850_),
    .B1(_00805_),
    .B2(_00851_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08623_ (.A1(_07159_),
    .A2(_00817_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08624_ (.A1(_00805_),
    .A2(_00742_),
    .A3(_00853_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08625_ (.A1(_00818_),
    .A2(_00852_),
    .A3(_00854_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08626_ (.A1(_07159_),
    .A2(_00595_),
    .A3(_07161_),
    .A4(_00729_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08627_ (.A1(_00850_),
    .A2(_00856_),
    .B(_00774_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08628_ (.A1(_00850_),
    .A2(_00856_),
    .B(_00583_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08629_ (.I0(_00857_),
    .I1(_00858_),
    .S(_00851_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08630_ (.A1(_00793_),
    .A2(_00805_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08631_ (.A1(_00736_),
    .A2(_00836_),
    .B(_00847_),
    .C(_07660_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08632_ (.I0(_00860_),
    .I1(_00861_),
    .S(_00742_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08633_ (.A1(net33),
    .A2(_00859_),
    .A3(_00862_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08634_ (.A1(_07180_),
    .A2(_00756_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08635_ (.A1(_00762_),
    .A2(net34),
    .A3(_00864_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08636_ (.A1(_00855_),
    .A2(_00863_),
    .B(_00865_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08637_ (.A1(_00851_),
    .A2(_00761_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08638_ (.A1(_00816_),
    .A2(_00866_),
    .B(_00768_),
    .C(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08639_ (.I(_00868_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08640_ (.A1(_00757_),
    .A2(_00851_),
    .A3(_00761_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08641_ (.A1(_07212_),
    .A2(_07218_),
    .A3(_07206_),
    .A4(_07209_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08642_ (.A1(_07203_),
    .A2(_07215_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08643_ (.A1(_07220_),
    .A2(_00591_),
    .A3(_00871_),
    .A4(_00872_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08644_ (.A1(_00570_),
    .A2(_00873_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08645_ (.A1(_00805_),
    .A2(_00873_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08646_ (.I0(_00874_),
    .I1(_00875_),
    .S(_00778_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08647_ (.A1(_00762_),
    .A2(net34),
    .A3(_00876_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08648_ (.A1(_00865_),
    .A2(_00870_),
    .A3(_00877_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08649_ (.A1(_00855_),
    .A2(_00863_),
    .B(_00878_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08650_ (.I(_00879_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08651_ (.A1(_07237_),
    .A2(_07236_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08652_ (.A1(_07235_),
    .A2(_00881_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08653_ (.A1(_00882_),
    .A2(_07234_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08654_ (.A1(_00883_),
    .A2(_07232_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08655_ (.A1(_00782_),
    .A2(_00780_),
    .A3(_00781_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08656_ (.A1(_00783_),
    .A2(_00885_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08657_ (.A1(_07791_),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08658_ (.A1(_00816_),
    .A2(_00880_),
    .B(_00884_),
    .C(_00887_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08659_ (.A1(_00818_),
    .A2(_00852_),
    .A3(_00854_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08660_ (.A1(net33),
    .A2(_00859_),
    .A3(_00862_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08661_ (.A1(_00889_),
    .A2(_00890_),
    .B(_00775_),
    .C(_00808_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08662_ (.A1(_07198_),
    .A2(_07200_),
    .A3(_07199_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08663_ (.A1(_00751_),
    .A2(_00892_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08664_ (.A1(_07176_),
    .A2(_00768_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08665_ (.A1(net18),
    .A2(_00805_),
    .A3(_00605_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _08666_ (.A1(_00772_),
    .A2(_00893_),
    .A3(_00762_),
    .B1(_00894_),
    .B2(_00895_),
    .B3(_00851_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08667_ (.I(_07176_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08668_ (.A1(_00897_),
    .A2(_00757_),
    .A3(_00759_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08669_ (.A1(_07660_),
    .A2(_00605_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08670_ (.A1(_00894_),
    .A2(_00899_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08671_ (.I0(_00898_),
    .I1(_00900_),
    .S(_00851_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08672_ (.A1(_00896_),
    .A2(_00901_),
    .B(_07791_),
    .C(_00884_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _08673_ (.I(_00884_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08674_ (.A1(_07791_),
    .A2(_00903_),
    .A3(_00896_),
    .A4(_00901_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08675_ (.A1(_00865_),
    .A2(_00870_),
    .A3(_00877_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08676_ (.A1(_00904_),
    .A2(_00902_),
    .B(_00814_),
    .C(_00905_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08677_ (.A1(_07226_),
    .A2(_07228_),
    .B(_07225_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08678_ (.A1(_07240_),
    .A2(_07231_),
    .B(_07239_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08679_ (.A1(_00907_),
    .A2(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08680_ (.A1(_00891_),
    .A2(_00906_),
    .B(_00909_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08681_ (.A1(_07226_),
    .A2(_07229_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08682_ (.A1(_00907_),
    .A2(_00911_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08683_ (.A1(_00910_),
    .A2(_00888_),
    .B(_00912_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _08684_ (.I(_07223_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08685_ (.A1(_00896_),
    .A2(_00901_),
    .Z(_07213_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08686_ (.A1(_07791_),
    .A2(_07213_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08687_ (.I(_00805_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08688_ (.I(_07191_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08689_ (.A1(_07194_),
    .A2(_00753_),
    .B(_07192_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08690_ (.I(_07189_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08691_ (.A1(_00917_),
    .A2(_00918_),
    .B(_00919_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08692_ (.A1(_07188_),
    .A2(_00920_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08693_ (.A1(_00745_),
    .A2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08694_ (.A1(_00762_),
    .A2(_00772_),
    .A3(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08695_ (.A1(_07117_),
    .A2(_07115_),
    .A3(_07116_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08696_ (.A1(_00611_),
    .A2(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08697_ (.I(_07102_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08698_ (.A1(_00926_),
    .A2(_00694_),
    .A3(_00639_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08699_ (.I0(_00925_),
    .I1(_00927_),
    .S(_00616_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08700_ (.I(_07119_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08701_ (.A1(_00929_),
    .A2(_00679_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08702_ (.A1(_07135_),
    .A2(_00930_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08703_ (.A1(_00645_),
    .A2(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08704_ (.A1(_07148_),
    .A2(_00662_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08705_ (.A1(_00654_),
    .A2(_00663_),
    .B(_00933_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08706_ (.A1(_00736_),
    .A2(_00928_),
    .B1(_00932_),
    .B2(_00670_),
    .C(_00934_),
    .ZN(_07163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08707_ (.A1(_00899_),
    .A2(_07163_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08708_ (.A1(_07165_),
    .A2(_07167_),
    .A3(_00602_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08709_ (.A1(_00727_),
    .A2(_00936_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08710_ (.A1(_00899_),
    .A2(_00937_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08711_ (.A1(_00935_),
    .A2(_00938_),
    .B(_00851_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08712_ (.A1(_00916_),
    .A2(_00923_),
    .A3(_00939_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08713_ (.A1(_00570_),
    .A2(_00762_),
    .A3(net34),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08714_ (.I0(_00570_),
    .I1(_00941_),
    .S(_00923_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08715_ (.A1(_00805_),
    .A2(_00851_),
    .A3(_00937_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08716_ (.A1(_00939_),
    .A2(_00943_),
    .B(_00916_),
    .C(_00773_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08717_ (.A1(_00940_),
    .A2(_00942_),
    .A3(_00944_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08718_ (.A1(_00581_),
    .A2(_07769_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08719_ (.A1(_07235_),
    .A2(_07237_),
    .A3(_07223_),
    .A4(_07232_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08720_ (.A1(_00947_),
    .A2(_00911_),
    .A3(_00946_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08721_ (.A1(_00915_),
    .A2(_00945_),
    .A3(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08722_ (.A1(net33),
    .A2(_00864_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08723_ (.A1(_00778_),
    .A2(_00762_),
    .A3(net34),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08724_ (.A1(_00809_),
    .A2(_00773_),
    .A3(_00812_),
    .B(_00951_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08725_ (.A1(_00889_),
    .A2(_00890_),
    .B(_00950_),
    .C(_00952_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08726_ (.A1(_00790_),
    .A2(_00570_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08727_ (.A1(_00788_),
    .A2(_00791_),
    .B1(_00954_),
    .B2(_00804_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08728_ (.A1(_00768_),
    .A2(_00955_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08729_ (.A1(_00768_),
    .A2(_00955_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08730_ (.A1(_00867_),
    .A2(_00956_),
    .B(_00957_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08731_ (.A1(_00809_),
    .A2(_00812_),
    .B(_00955_),
    .C(net33),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08732_ (.A1(_00803_),
    .A2(_00958_),
    .B(_00959_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08733_ (.A1(_00815_),
    .A2(_00879_),
    .A3(_00953_),
    .A4(_00960_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08734_ (.A1(_00952_),
    .A2(_00955_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08735_ (.I(_00887_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08736_ (.A1(_07203_),
    .A2(_07205_),
    .A3(_00786_),
    .A4(_00787_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08737_ (.A1(_00804_),
    .A2(_00964_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08738_ (.A1(_00805_),
    .A2(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08739_ (.I(_00966_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08740_ (.A1(_00948_),
    .A2(_00967_),
    .A3(_00963_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08741_ (.A1(_00870_),
    .A2(_00968_),
    .A3(_00962_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08742_ (.A1(_00815_),
    .A2(_00866_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08743_ (.A1(_00949_),
    .A2(_00961_),
    .B1(_00970_),
    .B2(_00969_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08744_ (.A1(_00571_),
    .A2(_00965_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08745_ (.A1(_00816_),
    .A2(_00880_),
    .B(_00972_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08746_ (.A1(_00939_),
    .A2(_00943_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08747_ (.A1(_00773_),
    .A2(_00974_),
    .B(_00923_),
    .ZN(_07201_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08748_ (.A1(_00570_),
    .A2(_00816_),
    .A3(_00880_),
    .A4(_07201_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08749_ (.A1(_07223_),
    .A2(_00973_),
    .A3(_00975_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08750_ (.A1(_00774_),
    .A2(_00570_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08751_ (.A1(_00816_),
    .A2(_00880_),
    .B(_00977_),
    .C(_00965_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08752_ (.A1(_00814_),
    .A2(_00808_),
    .A3(_00775_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08753_ (.A1(_00889_),
    .A2(_00890_),
    .B(_00905_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08754_ (.A1(_00979_),
    .A2(_00980_),
    .A3(_00977_),
    .A4(_07201_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08755_ (.A1(_00978_),
    .A2(_00981_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08756_ (.A1(_00914_),
    .A2(_00971_),
    .B1(_00976_),
    .B2(_00982_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08757_ (.A1(_00816_),
    .A2(_00880_),
    .B(_00966_),
    .C(_07222_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08758_ (.I(_07222_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08759_ (.A1(_00985_),
    .A2(_00815_),
    .A3(_00879_),
    .A4(_00945_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08760_ (.A1(_00984_),
    .A2(_00986_),
    .Z(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08761_ (.A1(_00815_),
    .A2(_00880_),
    .B(_00965_),
    .C(_00793_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08762_ (.A1(_00793_),
    .A2(_00979_),
    .A3(_00980_),
    .A4(_07201_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08763_ (.A1(_00988_),
    .A2(_00989_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08764_ (.A1(_00919_),
    .A2(_00917_),
    .A3(_00918_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08765_ (.I(_07173_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08766_ (.A1(_00992_),
    .A2(_00599_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08767_ (.A1(_07171_),
    .A2(_00993_),
    .B(_07170_),
    .C(_07168_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08768_ (.A1(_00602_),
    .A2(_00994_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08769_ (.A1(_07117_),
    .A2(net5),
    .ZN(_07118_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08770_ (.A1(_07120_),
    .A2(_07122_),
    .A3(_07121_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08771_ (.A1(_00679_),
    .A2(_00996_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08772_ (.I0(_07118_),
    .I1(_00997_),
    .S(_00645_),
    .Z(_07149_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08773_ (.A1(_07156_),
    .A2(_07155_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08774_ (.A1(_07154_),
    .A2(_00998_),
    .B(_07153_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08775_ (.A1(_07151_),
    .A2(_00999_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08776_ (.I0(_07149_),
    .I1(_01000_),
    .S(_00670_),
    .Z(_07166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _08777_ (.I0(_00916_),
    .I1(_00899_),
    .S(_00851_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08778_ (.I0(_00995_),
    .I1(_07166_),
    .S(_01001_),
    .Z(_07187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08779_ (.A1(_00802_),
    .A2(_07187_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08780_ (.A1(_00802_),
    .A2(_00920_),
    .A3(_00991_),
    .B(_01002_),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08781_ (.A1(_00779_),
    .A2(_00784_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08782_ (.A1(_07209_),
    .A2(_01003_),
    .B(_07208_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08783_ (.A1(_07206_),
    .A2(_01004_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08784_ (.A1(_00980_),
    .A2(_00979_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08785_ (.I0(_07204_),
    .I1(_01005_),
    .S(_01006_),
    .Z(_07221_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08786_ (.A1(_00971_),
    .A2(_00987_),
    .A3(_00990_),
    .A4(_07221_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08787_ (.A1(_00915_),
    .A2(_00945_),
    .A3(_00948_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08788_ (.A1(_00815_),
    .A2(_00880_),
    .A3(_00953_),
    .A4(_00960_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08789_ (.A1(_00870_),
    .A2(_00962_),
    .A3(_00968_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08790_ (.A1(_00979_),
    .A2(_00866_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08791_ (.A1(_01008_),
    .A2(_01009_),
    .B1(_01010_),
    .B2(_01011_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08792_ (.A1(_00984_),
    .A2(_00986_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08793_ (.A1(_00988_),
    .A2(_00989_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _08794_ (.A1(_01012_),
    .A2(_01013_),
    .A3(_01014_),
    .B1(_00913_),
    .B2(net21),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08795_ (.A1(_00913_),
    .A2(_00983_),
    .B1(_01007_),
    .B2(_01015_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08796_ (.A1(_00571_),
    .A2(_00594_),
    .B(_00869_),
    .C(_01016_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08797_ (.I(_00916_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08798_ (.I(_07251_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08799_ (.I(_07257_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08800_ (.A1(_07260_),
    .A2(_07259_),
    .B(_07258_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08801_ (.A1(_01021_),
    .A2(_01020_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08802_ (.A1(_01022_),
    .A2(_07255_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08803_ (.A1(_01023_),
    .A2(_07254_),
    .B(_07252_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08804_ (.A1(_01019_),
    .A2(_01024_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08805_ (.A1(_01025_),
    .A2(_07249_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08806_ (.A1(_01026_),
    .A2(_07248_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08807_ (.A1(_07246_),
    .A2(_01027_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08808_ (.A1(_01028_),
    .A2(_07245_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08809_ (.A1(_01029_),
    .A2(_07243_),
    .B(_07242_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08810_ (.A1(_01018_),
    .A2(_01030_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08811_ (.A1(_00571_),
    .A2(_01030_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08812_ (.A1(_00571_),
    .A2(_01030_),
    .B(_00774_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08813_ (.A1(_01032_),
    .A2(_01033_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08814_ (.I0(_01031_),
    .I1(_01034_),
    .S(_01016_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08815_ (.A1(_01017_),
    .A2(_01035_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08816_ (.A1(_00980_),
    .A2(_00979_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08817_ (.A1(_00816_),
    .A2(_00880_),
    .A3(_00945_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08818_ (.A1(_01037_),
    .A2(_00967_),
    .B(_01038_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08819_ (.A1(_07223_),
    .A2(_01039_),
    .A3(_00913_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08820_ (.A1(_01037_),
    .A2(_00955_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _08821_ (.A1(_00952_),
    .A2(_01041_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08822_ (.A1(_00916_),
    .A2(_00778_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08823_ (.A1(_01043_),
    .A2(_00873_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08824_ (.A1(_00870_),
    .A2(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08825_ (.A1(_00809_),
    .A2(_00812_),
    .B(_00570_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08826_ (.A1(_07104_),
    .A2(_00737_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08827_ (.A1(_00741_),
    .A2(_01047_),
    .A3(_00735_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08828_ (.A1(_00851_),
    .A2(_00761_),
    .B(_00570_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08829_ (.A1(_00757_),
    .A2(_00873_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08830_ (.A1(_01048_),
    .A2(_01049_),
    .B(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08831_ (.A1(_00773_),
    .A2(_01045_),
    .B1(_01046_),
    .B2(_01051_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08832_ (.A1(_00866_),
    .A2(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08833_ (.A1(_00816_),
    .A2(_00866_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08834_ (.A1(_00979_),
    .A2(_01053_),
    .B(_01054_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08835_ (.A1(_01012_),
    .A2(_00987_),
    .A3(_00990_),
    .A4(_01055_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08836_ (.A1(net6),
    .A2(_01042_),
    .A3(_01056_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08837_ (.A1(_00868_),
    .A2(_01057_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08838_ (.A1(_01018_),
    .A2(_01030_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08839_ (.I(_01033_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _08840_ (.I0(_01059_),
    .I1(_01060_),
    .S(_01016_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08841_ (.A1(_07223_),
    .A2(_00913_),
    .A3(_01039_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08842_ (.A1(_00952_),
    .A2(_01041_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08843_ (.A1(_01063_),
    .A2(_01056_),
    .B(_00971_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08844_ (.I0(_00866_),
    .I1(_01053_),
    .S(_00979_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08845_ (.A1(_07229_),
    .A2(_07239_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08846_ (.A1(_07228_),
    .A2(_01066_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08847_ (.A1(_07226_),
    .A2(_01067_),
    .B(_07225_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08848_ (.A1(_07231_),
    .A2(_00884_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08849_ (.A1(_07229_),
    .A2(_07228_),
    .B(_01069_),
    .C(_07226_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08850_ (.A1(_00816_),
    .A2(_00880_),
    .A3(_00915_),
    .A4(_01070_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08851_ (.I(_01070_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08852_ (.A1(_00816_),
    .A2(_00880_),
    .B(_00887_),
    .C(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08853_ (.A1(_01068_),
    .A2(_01071_),
    .A3(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08854_ (.A1(_01065_),
    .A2(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08855_ (.A1(_00987_),
    .A2(_00990_),
    .A3(_01065_),
    .A4(_01074_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08856_ (.A1(_01075_),
    .A2(_01076_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08857_ (.A1(_01062_),
    .A2(_01042_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08858_ (.A1(_00987_),
    .A2(_00990_),
    .B(_01065_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08859_ (.A1(_01042_),
    .A2(_01079_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08860_ (.A1(_01062_),
    .A2(_01064_),
    .B1(_01077_),
    .B2(_01078_),
    .C(_01080_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08861_ (.I0(_07201_),
    .I1(_00965_),
    .S(_01006_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08862_ (.A1(_00990_),
    .A2(_00971_),
    .A3(_00987_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08863_ (.A1(_00985_),
    .A2(_00916_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08864_ (.A1(_01068_),
    .A2(_01071_),
    .A3(_01073_),
    .A4(_01084_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08865_ (.A1(_01071_),
    .A2(_01073_),
    .B(_00914_),
    .C(_00916_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08866_ (.A1(_00914_),
    .A2(_00916_),
    .A3(_01068_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08867_ (.A1(_00914_),
    .A2(_00985_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08868_ (.I0(_07222_),
    .I1(_01088_),
    .S(_00916_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08869_ (.A1(_01085_),
    .A2(_01086_),
    .A3(_01087_),
    .A4(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08870_ (.A1(_01040_),
    .A2(_01083_),
    .B(_01090_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _08871_ (.A1(_01082_),
    .A2(_01091_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08872_ (.A1(_01058_),
    .A2(_01061_),
    .B(_01081_),
    .C(_01092_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08873_ (.A1(_00987_),
    .A2(_00990_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08874_ (.A1(_01042_),
    .A2(_01094_),
    .A3(_01065_),
    .B(_01012_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08875_ (.A1(_01075_),
    .A2(_01076_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08876_ (.A1(_01062_),
    .A2(_01042_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08877_ (.A1(_01042_),
    .A2(_01079_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _08878_ (.A1(_01040_),
    .A2(_01095_),
    .B1(_01096_),
    .B2(_01097_),
    .C(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08879_ (.A1(_00868_),
    .A2(_01057_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08880_ (.A1(_01018_),
    .A2(_01030_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08881_ (.A1(_00977_),
    .A2(_01030_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08882_ (.I0(_01101_),
    .I1(_01102_),
    .S(_01016_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08883_ (.A1(_01099_),
    .A2(_01092_),
    .A3(_01100_),
    .A4(_01103_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08884_ (.A1(_01036_),
    .A2(_01093_),
    .B(_01104_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08885_ (.A1(_01082_),
    .A2(_01091_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _08886_ (.I(_01106_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _08887_ (.I0(_01031_),
    .I1(_01033_),
    .S(_01016_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 clone31 (.I0(_01031_),
    .I1(_01033_),
    .S(_01016_),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08889_ (.A1(_00888_),
    .A2(_00910_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08890_ (.A1(_01110_),
    .A2(_00912_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08891_ (.A1(net21),
    .A2(_00973_),
    .A3(_00975_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08892_ (.A1(_00978_),
    .A2(_00981_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08893_ (.A1(net21),
    .A2(_01012_),
    .B1(_01112_),
    .B2(_01113_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08894_ (.A1(_01111_),
    .A2(_01114_),
    .B(_00594_),
    .C(_01018_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08895_ (.A1(_00571_),
    .A2(_00594_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08896_ (.A1(_01007_),
    .A2(_01015_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08897_ (.A1(_01007_),
    .A2(_01115_),
    .B1(_01116_),
    .B2(_01117_),
    .C(_00868_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08898_ (.A1(_07266_),
    .A2(_07263_),
    .A3(_07272_),
    .A4(_07280_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08899_ (.A1(_07277_),
    .A2(_07274_),
    .A3(_07269_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08900_ (.A1(_00591_),
    .A2(_01119_),
    .A3(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08901_ (.A1(_07243_),
    .A2(_01029_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08902_ (.A1(_01018_),
    .A2(_01121_),
    .A3(_01122_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08903_ (.A1(_00571_),
    .A2(_01121_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08904_ (.A1(_01122_),
    .A2(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08905_ (.A1(_01107_),
    .A2(net31),
    .A3(_01118_),
    .B1(_01123_),
    .B2(_01125_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08906_ (.A1(_07239_),
    .A2(_01069_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08907_ (.A1(_07229_),
    .A2(_01127_),
    .B(_07228_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08908_ (.I0(_01067_),
    .I1(_01128_),
    .S(_07226_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08909_ (.I(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08910_ (.I(_07226_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08911_ (.A1(_01131_),
    .A2(_07229_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08912_ (.A1(_01069_),
    .A2(_01132_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08913_ (.A1(_07228_),
    .A2(_07239_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08914_ (.A1(_07226_),
    .A2(_01134_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08915_ (.I0(_00915_),
    .I1(_00963_),
    .S(_01006_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08916_ (.I0(_01133_),
    .I1(_01135_),
    .S(_01136_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08917_ (.A1(net6),
    .A2(_01083_),
    .B1(_01130_),
    .B2(_01137_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08918_ (.A1(_07171_),
    .A2(_00993_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08919_ (.A1(_07122_),
    .A2(_00626_),
    .ZN(_07152_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08920_ (.A1(_07154_),
    .A2(_00998_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08921_ (.I0(_07152_),
    .I1(_01140_),
    .S(_00670_),
    .Z(_07169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08922_ (.I0(_01139_),
    .I1(_07169_),
    .S(_01001_),
    .Z(_07190_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08923_ (.A1(_07192_),
    .A2(_07194_),
    .A3(_00753_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08924_ (.A1(_00918_),
    .A2(_01141_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08925_ (.I0(_07190_),
    .I1(_01142_),
    .S(_00773_),
    .Z(_07207_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08926_ (.A1(_07209_),
    .A2(_01003_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08927_ (.I0(_07207_),
    .I1(_01143_),
    .S(_01006_),
    .Z(_07224_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08928_ (.A1(net6),
    .A2(_01083_),
    .A3(_07224_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08929_ (.A1(_01138_),
    .A2(_01144_),
    .B(_01124_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08930_ (.A1(_01107_),
    .A2(_01108_),
    .A3(_01118_),
    .A4(_01145_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08931_ (.A1(_01018_),
    .A2(_01121_),
    .A3(_01138_),
    .A4(_01144_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08932_ (.A1(_01107_),
    .A2(_01108_),
    .A3(_01118_),
    .A4(_01147_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08933_ (.A1(_01126_),
    .A2(_01146_),
    .A3(_01148_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08934_ (.A1(_01111_),
    .A2(_01114_),
    .B(_01117_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08935_ (.A1(_01092_),
    .A2(_01061_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08936_ (.A1(_01069_),
    .A2(_01132_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08937_ (.A1(_07226_),
    .A2(_01134_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08938_ (.I0(_01152_),
    .I1(_01153_),
    .S(_01136_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _08939_ (.A1(_01062_),
    .A2(_01012_),
    .A3(_01094_),
    .B1(_01129_),
    .B2(_01154_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08940_ (.A1(_01040_),
    .A2(_01083_),
    .A3(_07224_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08941_ (.I(_07265_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08942_ (.A1(_07274_),
    .A2(_07273_),
    .B(_07266_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08943_ (.A1(_01157_),
    .A2(_01158_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08944_ (.A1(_01159_),
    .A2(_07263_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08945_ (.A1(_07262_),
    .A2(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08946_ (.A1(_07272_),
    .A2(_01161_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08947_ (.A1(_07271_),
    .A2(_01162_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08948_ (.A1(_07269_),
    .A2(_01163_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08949_ (.A1(_01164_),
    .A2(_07268_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08950_ (.A1(_07280_),
    .A2(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08951_ (.A1(_01166_),
    .A2(_07279_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08952_ (.A1(_07277_),
    .A2(_01167_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08953_ (.A1(_01168_),
    .A2(_07276_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08954_ (.A1(_01155_),
    .A2(_01156_),
    .B(_01169_),
    .C(_00571_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08955_ (.A1(_01168_),
    .A2(_07276_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08956_ (.A1(_01171_),
    .A2(_01155_),
    .A3(_01156_),
    .A4(_00571_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08957_ (.A1(_01155_),
    .A2(_01156_),
    .B(_00774_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08958_ (.A1(_01170_),
    .A2(_01173_),
    .A3(_01172_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08959_ (.A1(_00571_),
    .A2(_00913_),
    .A3(_00594_),
    .A4(_00983_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08960_ (.A1(_01018_),
    .A2(_00913_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08961_ (.A1(_00914_),
    .A2(_01176_),
    .B(_01115_),
    .C(_01083_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08962_ (.A1(_01099_),
    .A2(_01118_),
    .A3(_01175_),
    .A4(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08963_ (.A1(_01150_),
    .A2(_01151_),
    .A3(_01174_),
    .A4(_01178_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08964_ (.A1(_07243_),
    .A2(_01029_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08965_ (.A1(_01018_),
    .A2(_01122_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08966_ (.A1(_01171_),
    .A2(_01181_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08967_ (.A1(_00774_),
    .A2(_01180_),
    .B(_01182_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08968_ (.A1(_01016_),
    .A2(_01032_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08969_ (.A1(_01183_),
    .A2(_01184_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08970_ (.A1(_01106_),
    .A2(_01099_),
    .A3(_01108_),
    .A4(_01118_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _08971_ (.I(_01186_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08972_ (.A1(_01185_),
    .A2(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08973_ (.A1(_01105_),
    .A2(_01149_),
    .B1(_01179_),
    .B2(_01188_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08974_ (.A1(_01183_),
    .A2(_01184_),
    .A3(_01187_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08975_ (.A1(_01150_),
    .A2(_01174_),
    .A3(net28),
    .B(_01190_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08976_ (.A1(_01189_),
    .A2(_01191_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08977_ (.A1(_01189_),
    .A2(_01191_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08978_ (.A1(_01099_),
    .A2(_01118_),
    .A3(_01175_),
    .A4(_01177_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08979_ (.A1(_01151_),
    .A2(_01194_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08980_ (.A1(_01107_),
    .A2(net31),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08981_ (.A1(_01195_),
    .A2(_01196_),
    .B(_01185_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08982_ (.A1(_01099_),
    .A2(_01106_),
    .A3(_01108_),
    .A4(_01118_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _08983_ (.A1(_01099_),
    .A2(_01170_),
    .A3(_01172_),
    .A4(_01173_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08984_ (.A1(_01107_),
    .A2(net31),
    .A3(_01118_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08985_ (.A1(_00572_),
    .A2(_01169_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08986_ (.A1(_01183_),
    .A2(_01198_),
    .B1(_01199_),
    .B2(_01200_),
    .C(_01201_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08987_ (.A1(_01036_),
    .A2(_01093_),
    .B(_01201_),
    .C(_01104_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08988_ (.A1(_01155_),
    .A2(_01156_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08989_ (.I(_01204_),
    .ZN(_07241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08990_ (.I0(_07241_),
    .I1(_01122_),
    .S(_01186_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08991_ (.A1(_01202_),
    .A2(_01203_),
    .A3(_01205_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08992_ (.A1(_01202_),
    .A2(_01203_),
    .B(_01205_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08993_ (.A1(_01197_),
    .A2(_01206_),
    .A3(_01207_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08994_ (.A1(_01193_),
    .A2(_01208_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08995_ (.A1(_01017_),
    .A2(_01035_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08996_ (.A1(_01100_),
    .A2(net31),
    .B(_01099_),
    .C(_01107_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _08997_ (.A1(_01099_),
    .A2(_01092_),
    .A3(_01100_),
    .A4(_01103_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08998_ (.A1(_01210_),
    .A2(_01211_),
    .B(_01212_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08999_ (.A1(_00793_),
    .A2(_01122_),
    .B1(_01171_),
    .B2(_01181_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09000_ (.A1(_01099_),
    .A2(_01170_),
    .A3(_01172_),
    .A4(_01173_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09001_ (.A1(_01106_),
    .A2(_01108_),
    .A3(_01118_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09002_ (.A1(_01214_),
    .A2(_01186_),
    .B1(_01215_),
    .B2(_01216_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _09003_ (.A1(_07277_),
    .A2(_01167_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _09004_ (.I(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09005_ (.A1(_00572_),
    .A2(_01219_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09006_ (.I(_01018_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09007_ (.A1(_01221_),
    .A2(_01218_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _09008_ (.A1(_01213_),
    .A2(_01217_),
    .B1(_01220_),
    .B2(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09009_ (.A1(_00752_),
    .A2(_00750_),
    .A3(_00751_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09010_ (.A1(_07176_),
    .A2(_07174_),
    .A3(_07175_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09011_ (.A1(_00599_),
    .A2(_01225_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09012_ (.A1(_00650_),
    .A2(_00678_),
    .B(_00916_),
    .C(_07156_),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09013_ (.I0(_01226_),
    .I1(_07172_),
    .S(_01001_),
    .Z(_07193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09014_ (.A1(_00802_),
    .A2(_07193_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09015_ (.A1(_00753_),
    .A2(_00802_),
    .A3(_01224_),
    .B(_01227_),
    .ZN(_07210_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09016_ (.A1(_07212_),
    .A2(_07214_),
    .A3(_00783_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09017_ (.A1(_00784_),
    .A2(_01228_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09018_ (.I0(_07210_),
    .I1(_01229_),
    .S(_01006_),
    .Z(_07227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09019_ (.A1(_00891_),
    .A2(_00906_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09020_ (.A1(_00908_),
    .A2(_00888_),
    .A3(_01230_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09021_ (.A1(_07229_),
    .A2(_01231_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09022_ (.A1(_01083_),
    .A2(_01040_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09023_ (.I0(_07227_),
    .I1(_01232_),
    .S(_01233_),
    .Z(_07244_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09024_ (.I(_07244_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09025_ (.A1(_07246_),
    .A2(_01027_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09026_ (.I(_01235_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09027_ (.I0(_01234_),
    .I1(_01236_),
    .S(_01186_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09028_ (.A1(_00572_),
    .A2(_01213_),
    .A3(_01217_),
    .A4(_01237_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09029_ (.A1(_07300_),
    .A2(_07292_),
    .A3(_07295_),
    .A4(_07298_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09030_ (.A1(_07283_),
    .A2(_07286_),
    .A3(_07289_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09031_ (.A1(_00591_),
    .A2(_01239_),
    .A3(_01240_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09032_ (.A1(_01223_),
    .A2(_01238_),
    .B(_01241_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09033_ (.A1(_01105_),
    .A2(_01149_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09034_ (.A1(_01062_),
    .A2(_00971_),
    .A3(_01094_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09035_ (.A1(_01042_),
    .A2(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09036_ (.A1(_01092_),
    .A2(_01061_),
    .A3(_01245_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09037_ (.A1(_01092_),
    .A2(_01061_),
    .B(_01245_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09038_ (.A1(_01194_),
    .A2(_01246_),
    .B(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09039_ (.A1(_01107_),
    .A2(_01103_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09040_ (.A1(_01035_),
    .A2(_01107_),
    .B(_01214_),
    .C(_01249_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09041_ (.A1(_01179_),
    .A2(_01248_),
    .A3(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09042_ (.A1(_01179_),
    .A2(_01250_),
    .B(_01248_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09043_ (.A1(_01243_),
    .A2(_01251_),
    .A3(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09044_ (.A1(net21),
    .A2(_01039_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09045_ (.A1(_00987_),
    .A2(_00990_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09046_ (.A1(_01254_),
    .A2(_01074_),
    .B(_01255_),
    .C(_01042_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09047_ (.A1(net6),
    .A2(_00971_),
    .B(_01256_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09048_ (.I0(_01256_),
    .I1(_01257_),
    .S(_01055_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09049_ (.A1(_01246_),
    .A2(_01258_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09050_ (.A1(_01100_),
    .A2(_01259_),
    .B(net28),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _09051_ (.I(_01237_),
    .ZN(_07275_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09052_ (.A1(_01017_),
    .A2(_01035_),
    .A3(_01107_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09053_ (.A1(_01107_),
    .A2(_01103_),
    .B(_01099_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09054_ (.A1(_01261_),
    .A2(_01262_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09055_ (.I(_01241_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09056_ (.A1(_00572_),
    .A2(_01264_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09057_ (.A1(_01217_),
    .A2(_07275_),
    .A3(_01263_),
    .A4(_01265_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09058_ (.A1(_01092_),
    .A2(_01061_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09059_ (.A1(_01063_),
    .A2(_01244_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09060_ (.A1(_01267_),
    .A2(_01268_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09061_ (.A1(_01081_),
    .A2(_01061_),
    .B(_01058_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _09062_ (.A1(_01100_),
    .A2(_01262_),
    .B1(_01270_),
    .B2(_01261_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09063_ (.A1(_01269_),
    .A2(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09064_ (.A1(_01179_),
    .A2(_01250_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09065_ (.A1(_01260_),
    .A2(_01266_),
    .B1(_01272_),
    .B2(_01273_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09066_ (.A1(_01242_),
    .A2(_01253_),
    .A3(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09067_ (.I0(_01174_),
    .I1(_01214_),
    .S(_01186_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09068_ (.I(_01276_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09069_ (.A1(_01105_),
    .A2(net42),
    .A3(_07275_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09070_ (.I(_01105_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09071_ (.A1(_01279_),
    .A2(net42),
    .B(_01219_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09072_ (.I(_00774_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09073_ (.I(_07297_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09074_ (.A1(_07300_),
    .A2(_07299_),
    .B(_07298_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09075_ (.A1(_01282_),
    .A2(_01283_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09076_ (.A1(_01284_),
    .A2(_07295_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09077_ (.A1(_07294_),
    .A2(_01285_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09078_ (.A1(_07292_),
    .A2(_01286_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09079_ (.A1(_01287_),
    .A2(_07291_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09080_ (.A1(_07289_),
    .A2(_01288_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09081_ (.A1(_01289_),
    .A2(_07288_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09082_ (.A1(_07286_),
    .A2(_01290_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09083_ (.A1(_07285_),
    .A2(_01291_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09084_ (.A1(_07283_),
    .A2(_01292_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09085_ (.A1(_01293_),
    .A2(_07282_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09086_ (.I(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09087_ (.A1(_01295_),
    .A2(_01221_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09088_ (.A1(_01281_),
    .A2(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09089_ (.A1(_01278_),
    .A2(_01280_),
    .B(_01297_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09090_ (.A1(_07282_),
    .A2(_01293_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09091_ (.A1(_01221_),
    .A2(_01278_),
    .A3(_01280_),
    .A4(_01299_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09092_ (.A1(_01298_),
    .A2(_01300_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09093_ (.A1(_01189_),
    .A2(_01191_),
    .A3(_01206_),
    .A4(_01207_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09094_ (.A1(_01018_),
    .A2(_01169_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _09095_ (.A1(_01214_),
    .A2(net28),
    .B1(_01215_),
    .B2(_01216_),
    .C(_01303_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09096_ (.A1(_01210_),
    .A2(_01211_),
    .B(_01303_),
    .C(_01212_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09097_ (.I0(_01204_),
    .I1(_01180_),
    .S(net28),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09098_ (.A1(_01304_),
    .A2(_01305_),
    .A3(_01306_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09099_ (.A1(_01304_),
    .A2(_01305_),
    .B(_01306_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09100_ (.A1(_01307_),
    .A2(_01308_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _09101_ (.A1(_01192_),
    .A2(_01309_),
    .A3(_01298_),
    .A4(_01300_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09102_ (.A1(_01209_),
    .A2(_01275_),
    .B1(_01301_),
    .B2(_01302_),
    .C(_01310_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09103_ (.A1(_01213_),
    .A2(_01217_),
    .A3(_01237_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09104_ (.A1(_01213_),
    .A2(_01217_),
    .B(_01218_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09105_ (.A1(_01312_),
    .A2(_01313_),
    .B1(_00774_),
    .B2(_01296_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _09106_ (.A1(_00572_),
    .A2(_01295_),
    .A3(_01313_),
    .A4(_01312_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09107_ (.A1(_01193_),
    .A2(_01208_),
    .A3(_01314_),
    .A4(_01315_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09108_ (.A1(_01279_),
    .A2(_01149_),
    .B1(_01179_),
    .B2(_01250_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09109_ (.A1(_01197_),
    .A2(_01317_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09110_ (.A1(_01081_),
    .A2(_01092_),
    .A3(_01061_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09111_ (.A1(_01058_),
    .A2(_01319_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09112_ (.A1(_01183_),
    .A2(_01263_),
    .B(_01320_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09113_ (.A1(_01118_),
    .A2(_01175_),
    .A3(_01177_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09114_ (.A1(_01322_),
    .A2(_01319_),
    .B1(_01268_),
    .B2(_01258_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09115_ (.A1(_01267_),
    .A2(_01258_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09116_ (.A1(_01323_),
    .A2(_01324_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09117_ (.A1(_01318_),
    .A2(_01321_),
    .A3(_01325_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09118_ (.A1(_01253_),
    .A2(_01316_),
    .B(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09119_ (.A1(_01311_),
    .A2(_01327_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09120_ (.A1(_00572_),
    .A2(_01219_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09121_ (.A1(_01221_),
    .A2(_01218_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09122_ (.A1(_01279_),
    .A2(net42),
    .B1(_01329_),
    .B2(_01330_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09123_ (.A1(_01221_),
    .A2(_01279_),
    .A3(_01277_),
    .A4(_07275_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09124_ (.A1(_01331_),
    .A2(_01332_),
    .B(_01264_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09125_ (.A1(_01243_),
    .A2(_01251_),
    .A3(_01252_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09126_ (.A1(_01246_),
    .A2(_01258_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09127_ (.A1(_01058_),
    .A2(_01335_),
    .B(_01198_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09128_ (.A1(_01217_),
    .A2(_07275_),
    .A3(_01263_),
    .A4(_01265_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09129_ (.A1(_01269_),
    .A2(_01271_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09130_ (.A1(_01179_),
    .A2(_01250_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _09131_ (.A1(_01336_),
    .A2(_01337_),
    .B1(_01338_),
    .B2(_01339_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09132_ (.A1(_01333_),
    .A2(_01334_),
    .A3(_01340_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09133_ (.I(_01341_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09134_ (.A1(_01314_),
    .A2(_01208_),
    .A3(_01193_),
    .A4(_01315_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09135_ (.I(_01343_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09136_ (.A1(_07283_),
    .A2(_01292_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09137_ (.A1(_01221_),
    .A2(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09138_ (.A1(_01342_),
    .A2(net38),
    .B(_01346_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09139_ (.A1(_07280_),
    .A2(_01165_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09140_ (.A1(_01279_),
    .A2(_01277_),
    .B(_01348_),
    .C(_01166_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09141_ (.I0(_07213_),
    .I1(_00886_),
    .S(_01006_),
    .Z(_07238_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09142_ (.A1(_07240_),
    .A2(_01069_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09143_ (.I0(_07238_),
    .I1(_01350_),
    .S(_01233_),
    .Z(_07247_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09144_ (.A1(_07249_),
    .A2(_01025_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09145_ (.I0(_07247_),
    .I1(_01351_),
    .S(_01186_),
    .Z(_07278_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09146_ (.A1(_01279_),
    .A2(_01277_),
    .A3(_07278_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09147_ (.A1(_01349_),
    .A2(_01352_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09148_ (.I(_01353_),
    .ZN(_07281_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09149_ (.A1(_00573_),
    .A2(_01341_),
    .A3(_01343_),
    .A4(_07281_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09150_ (.A1(_01312_),
    .A2(_01313_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09151_ (.A1(_00793_),
    .A2(_01219_),
    .A3(net32),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09152_ (.A1(_01279_),
    .A2(net42),
    .B(_01356_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09153_ (.A1(_00774_),
    .A2(_01299_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09154_ (.A1(_01279_),
    .A2(net42),
    .A3(_07275_),
    .A4(_01358_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09155_ (.A1(_01307_),
    .A2(_01308_),
    .B(_01357_),
    .C(_01359_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09156_ (.A1(_01122_),
    .A2(_01236_),
    .A3(_01299_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09157_ (.A1(_01180_),
    .A2(_01235_),
    .A3(_01295_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09158_ (.A1(_01198_),
    .A2(_01361_),
    .A3(_01362_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09159_ (.A1(_01204_),
    .A2(_07244_),
    .A3(net32),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09160_ (.A1(_01204_),
    .A2(_07244_),
    .A3(_01295_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09161_ (.A1(net28),
    .A2(_01364_),
    .A3(_01365_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09162_ (.A1(_01363_),
    .A2(_01366_),
    .B(_00572_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09163_ (.A1(_01219_),
    .A2(_01299_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09164_ (.A1(_01218_),
    .A2(_01294_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09165_ (.I(_01369_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09166_ (.A1(_01204_),
    .A2(_01169_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09167_ (.I0(_01368_),
    .I1(_01370_),
    .S(_01371_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09168_ (.A1(_01169_),
    .A2(_01218_),
    .A3(_01295_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09169_ (.A1(_01171_),
    .A2(_01219_),
    .A3(_01299_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09170_ (.A1(_01373_),
    .A2(_01374_),
    .B(_01180_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09171_ (.A1(_01198_),
    .A2(_01375_),
    .B(_01221_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09172_ (.A1(_01169_),
    .A2(_01369_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09173_ (.A1(_01169_),
    .A2(_01368_),
    .B(_01377_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09174_ (.A1(_01180_),
    .A2(_01198_),
    .A3(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09175_ (.A1(_01198_),
    .A2(_01372_),
    .B(_01376_),
    .C(_01379_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09176_ (.A1(_01277_),
    .A2(_01279_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09177_ (.I0(_01367_),
    .I1(_01380_),
    .S(_01381_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09178_ (.A1(_00573_),
    .A2(_01360_),
    .B(_01382_),
    .C(_01193_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09179_ (.I(_01221_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09180_ (.A1(_01312_),
    .A2(_01313_),
    .B(net32),
    .C(_01281_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09181_ (.A1(_01312_),
    .A2(_01313_),
    .A3(net32),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09182_ (.A1(_01384_),
    .A2(_01309_),
    .A3(_01385_),
    .A4(_01386_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09183_ (.A1(_01355_),
    .A2(_01343_),
    .B1(_01383_),
    .B2(_01387_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _09184_ (.A1(_01243_),
    .A2(_01251_),
    .A3(_01252_),
    .B1(_01349_),
    .B2(_01352_),
    .B3(_00573_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09185_ (.A1(_01242_),
    .A2(_01274_),
    .A3(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _09186_ (.A1(_01314_),
    .A2(_01315_),
    .A3(_01302_),
    .B1(_01317_),
    .B2(_01197_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09187_ (.I(_00591_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09188_ (.A1(_07303_),
    .A2(_07306_),
    .A3(_07309_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09189_ (.A1(_07320_),
    .A2(_07312_),
    .A3(_07315_),
    .A4(_07318_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09190_ (.A1(_01392_),
    .A2(_01393_),
    .A3(_01394_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09191_ (.A1(_01316_),
    .A2(_01390_),
    .B(_01391_),
    .C(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09192_ (.A1(_01347_),
    .A2(_01354_),
    .A3(_01388_),
    .A4(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09193_ (.I(_01309_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09194_ (.A1(_07283_),
    .A2(_01292_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09195_ (.A1(_07309_),
    .A2(_07311_),
    .B(_07308_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09196_ (.I(_07317_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09197_ (.A1(_07320_),
    .A2(_07319_),
    .B(_07318_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09198_ (.A1(_01401_),
    .A2(_01402_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09199_ (.A1(_01403_),
    .A2(_07315_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09200_ (.A1(_01404_),
    .A2(_07314_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09201_ (.A1(_07312_),
    .A2(_01405_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09202_ (.A1(_01406_),
    .A2(_07309_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09203_ (.A1(_01400_),
    .A2(_01407_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09204_ (.A1(_07306_),
    .A2(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09205_ (.A1(_01409_),
    .A2(_07305_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09206_ (.A1(_07303_),
    .A2(_01410_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09207_ (.A1(_01411_),
    .A2(_07302_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09208_ (.A1(_01412_),
    .A2(_01346_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09209_ (.A1(_00774_),
    .A2(_01399_),
    .B(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09210_ (.A1(_01221_),
    .A2(_01299_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09211_ (.A1(_01415_),
    .A2(_01414_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09212_ (.I(_01416_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09213_ (.A1(_00793_),
    .A2(_01345_),
    .B1(_01346_),
    .B2(_01412_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09214_ (.A1(_01418_),
    .A2(_01415_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09215_ (.I0(_01417_),
    .I1(_01419_),
    .S(_01355_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09216_ (.A1(_01398_),
    .A2(_01420_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09217_ (.A1(_01298_),
    .A2(_01300_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09218_ (.A1(_01193_),
    .A2(_01208_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09219_ (.A1(_01423_),
    .A2(_01342_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09220_ (.A1(_01312_),
    .A2(_01313_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09221_ (.A1(_07302_),
    .A2(_01411_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09222_ (.A1(_00572_),
    .A2(_01426_),
    .B(_01281_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09223_ (.A1(_00572_),
    .A2(_01412_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09224_ (.I0(_01427_),
    .I1(_01428_),
    .S(_01353_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09225_ (.A1(_01425_),
    .A2(_01429_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _09226_ (.A1(_01424_),
    .A2(_01422_),
    .A3(_01430_),
    .B1(_01420_),
    .B2(_01398_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _09227_ (.A1(_01328_),
    .A2(_01397_),
    .B1(_01421_),
    .B2(_01422_),
    .C(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09228_ (.A1(_01192_),
    .A2(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09229_ (.I(_01316_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09230_ (.A1(_01333_),
    .A2(_01340_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09231_ (.A1(_01253_),
    .A2(_01435_),
    .A3(_01316_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09232_ (.A1(_01253_),
    .A2(_01434_),
    .B(_01436_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09233_ (.I(_01275_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09234_ (.A1(_01425_),
    .A2(_01429_),
    .A3(_01316_),
    .A4(_01438_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09235_ (.A1(_01438_),
    .A2(_01434_),
    .B(_01420_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09236_ (.A1(_01192_),
    .A2(_01309_),
    .A3(_01298_),
    .A4(_01300_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09237_ (.A1(_01298_),
    .A2(_01300_),
    .B(_01302_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09238_ (.A1(_01423_),
    .A2(_01342_),
    .B(_01441_),
    .C(_01442_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09239_ (.A1(_01318_),
    .A2(_01321_),
    .A3(_01325_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09240_ (.A1(_01334_),
    .A2(_01344_),
    .B(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09241_ (.A1(_01440_),
    .A2(_01439_),
    .B(_01443_),
    .C(_01445_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09242_ (.A1(_01383_),
    .A2(_01387_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09243_ (.A1(_01312_),
    .A2(_01313_),
    .B(net32),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09244_ (.A1(_01448_),
    .A2(_01386_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09245_ (.A1(_00573_),
    .A2(_01399_),
    .A3(_01393_),
    .A4(_01406_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09246_ (.I(_01400_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09247_ (.A1(_07306_),
    .A2(_01451_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09248_ (.A1(_07305_),
    .A2(_01452_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09249_ (.A1(_07303_),
    .A2(_01453_),
    .B(_07302_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09250_ (.A1(_00573_),
    .A2(_01454_),
    .B(_01281_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09251_ (.A1(_01384_),
    .A2(_01454_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09252_ (.I0(_01455_),
    .I1(_01456_),
    .S(_01399_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _09253_ (.A1(_01384_),
    .A2(_01345_),
    .A3(_01393_),
    .A4(_01406_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09254_ (.A1(_01448_),
    .A2(_01386_),
    .A3(_01458_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09255_ (.A1(_01449_),
    .A2(_01450_),
    .B(_01457_),
    .C(_01459_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09256_ (.A1(_01429_),
    .A2(_01438_),
    .A3(_01316_),
    .A4(_01425_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09257_ (.A1(_01447_),
    .A2(_01460_),
    .B(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09258_ (.A1(_01446_),
    .A2(_01462_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09259_ (.A1(_01437_),
    .A2(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09260_ (.A1(_01342_),
    .A2(_01434_),
    .B(_01391_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09261_ (.A1(_01437_),
    .A2(_01463_),
    .A3(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _09262_ (.A1(_01433_),
    .A2(_01464_),
    .B1(_01465_),
    .B2(_01437_),
    .C(_01466_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09263_ (.A1(_01446_),
    .A2(_01462_),
    .A3(_01465_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09264_ (.A1(_01462_),
    .A2(_01465_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09265_ (.A1(_01468_),
    .A2(_01469_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09266_ (.A1(_01221_),
    .A2(_01426_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09267_ (.A1(_01399_),
    .A2(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09268_ (.A1(_01438_),
    .A2(_01434_),
    .B(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09269_ (.A1(_01438_),
    .A2(_01316_),
    .A3(_01353_),
    .A4(_01471_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09270_ (.A1(_01438_),
    .A2(_01434_),
    .B(_01399_),
    .C(_01471_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _09271_ (.A1(_01342_),
    .A2(_01344_),
    .A3(_01353_),
    .A4(_01471_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09272_ (.A1(_01473_),
    .A2(_01474_),
    .A3(_01475_),
    .A4(_01476_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09273_ (.A1(_01438_),
    .A2(_01316_),
    .A3(_01429_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09274_ (.A1(_01414_),
    .A2(_01415_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09275_ (.A1(_01438_),
    .A2(_01434_),
    .B(_01416_),
    .C(_01479_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09276_ (.A1(_01425_),
    .A2(_01478_),
    .A3(_01480_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09277_ (.A1(_01478_),
    .A2(_01480_),
    .B(_01425_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09278_ (.A1(_01355_),
    .A2(_01415_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09279_ (.A1(_01355_),
    .A2(_01415_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _09280_ (.A1(_01341_),
    .A2(_01344_),
    .B1(_01483_),
    .B2(_01484_),
    .C(_01414_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09281_ (.A1(_01485_),
    .A2(_01461_),
    .B(_01311_),
    .C(_01327_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09282_ (.I(_01486_),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09283_ (.A1(_01343_),
    .A2(_01341_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09284_ (.I0(_07281_),
    .I1(_01345_),
    .S(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _09285_ (.A1(_01477_),
    .A2(_01481_),
    .A3(_01482_),
    .B1(_01487_),
    .B2(_01489_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09286_ (.I(_01488_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _09287_ (.A1(_07286_),
    .A2(_01290_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09288_ (.A1(_07200_),
    .A2(_00802_),
    .ZN(_07216_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09289_ (.A1(_07218_),
    .A2(_07220_),
    .A3(_07219_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09290_ (.A1(_00781_),
    .A2(_01493_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09291_ (.I0(_07216_),
    .I1(_01494_),
    .S(_01006_),
    .Z(_07230_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09292_ (.A1(_07232_),
    .A2(_00883_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09293_ (.I0(_07230_),
    .I1(_01495_),
    .S(_01233_),
    .Z(_07250_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09294_ (.A1(_07252_),
    .A2(_07254_),
    .A3(_01023_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09295_ (.A1(_01024_),
    .A2(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09296_ (.I0(_07250_),
    .I1(_01497_),
    .S(_01187_),
    .Z(_07267_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09297_ (.I(_07267_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09298_ (.A1(_07269_),
    .A2(_01163_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09299_ (.I0(_01498_),
    .I1(_01499_),
    .S(_01381_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09300_ (.A1(_01342_),
    .A2(_01344_),
    .A3(_01500_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09301_ (.I(_07337_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09302_ (.A1(_07340_),
    .A2(_07339_),
    .B(_07338_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09303_ (.A1(_01503_),
    .A2(_01502_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09304_ (.A1(_07335_),
    .A2(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09305_ (.A1(_07334_),
    .A2(_01505_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09306_ (.A1(_07332_),
    .A2(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09307_ (.A1(_01507_),
    .A2(_07331_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09308_ (.A1(_07329_),
    .A2(_01508_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09309_ (.A1(_01509_),
    .A2(_07328_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09310_ (.A1(_07326_),
    .A2(_01510_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09311_ (.A1(_01511_),
    .A2(_07325_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09312_ (.A1(_01512_),
    .A2(_07323_),
    .B(_07322_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _09313_ (.I(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09314_ (.A1(_01384_),
    .A2(_01514_),
    .B(_00793_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09315_ (.A1(net13),
    .A2(_01492_),
    .B(_01501_),
    .C(_01515_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09316_ (.A1(_01514_),
    .A2(_00573_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09317_ (.A1(_01500_),
    .A2(_01517_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09318_ (.A1(_01492_),
    .A2(_01517_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09319_ (.I0(_01518_),
    .I1(_01519_),
    .S(net13),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09320_ (.A1(_01516_),
    .A2(_01520_),
    .B(_01446_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09321_ (.A1(_01311_),
    .A2(_01327_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09322_ (.I(_01517_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09323_ (.A1(_07303_),
    .A2(_01410_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09324_ (.I0(_01523_),
    .I1(_01515_),
    .S(_01524_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _09325_ (.I(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09326_ (.A1(_01526_),
    .A2(_01439_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09327_ (.A1(_01522_),
    .A2(_01526_),
    .B1(_01440_),
    .B2(_01527_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _09328_ (.A1(_01311_),
    .A2(_01490_),
    .A3(_01528_),
    .A4(_01521_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09329_ (.A1(_01437_),
    .A2(_01470_),
    .A3(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09330_ (.A1(_01467_),
    .A2(_01530_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09331_ (.A1(_01490_),
    .A2(_01521_),
    .A3(_01528_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09332_ (.A1(_01309_),
    .A2(_01422_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09333_ (.A1(_01424_),
    .A2(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09334_ (.A1(_01347_),
    .A2(_01354_),
    .A3(_01388_),
    .A4(_01396_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09335_ (.A1(_01439_),
    .A2(_01440_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09336_ (.A1(_01522_),
    .A2(_01535_),
    .B(_01536_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09337_ (.A1(_01534_),
    .A2(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09338_ (.A1(_01532_),
    .A2(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09339_ (.A1(_01425_),
    .A2(_01438_),
    .A3(_01434_),
    .B(_01484_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09340_ (.A1(_01342_),
    .A2(net38),
    .B(_01483_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09341_ (.A1(_01540_),
    .A2(_01541_),
    .B(_01311_),
    .C(_01327_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09342_ (.A1(_01438_),
    .A2(_01434_),
    .B(_01418_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09343_ (.A1(_01435_),
    .A2(_01434_),
    .B(_01391_),
    .C(_01334_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09344_ (.A1(_01478_),
    .A2(_01543_),
    .B(_01544_),
    .C(_01388_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09345_ (.A1(_01535_),
    .A2(_01542_),
    .B(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09346_ (.A1(_01217_),
    .A2(_01263_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09347_ (.A1(_01317_),
    .A2(_01324_),
    .B(_01323_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09348_ (.A1(_01547_),
    .A2(_01320_),
    .B(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09349_ (.A1(_01436_),
    .A2(_01549_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _09350_ (.A1(_01546_),
    .A2(_01550_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09351_ (.A1(_01437_),
    .A2(_01468_),
    .A3(_01469_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09352_ (.A1(_00573_),
    .A2(_01524_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09353_ (.A1(_07338_),
    .A2(_07329_),
    .A3(_07332_),
    .A4(_07335_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09354_ (.A1(_07340_),
    .A2(_07323_),
    .A3(_07326_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09355_ (.A1(_01392_),
    .A2(_01554_),
    .A3(_01555_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09356_ (.A1(_01553_),
    .A2(_01556_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09357_ (.A1(_01321_),
    .A2(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09358_ (.A1(_01334_),
    .A2(net38),
    .B(_01318_),
    .C(_01325_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09359_ (.A1(_01439_),
    .A2(_01440_),
    .B(_01443_),
    .C(_01559_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09360_ (.A1(_01253_),
    .A2(_01435_),
    .A3(_01434_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09361_ (.I(_01321_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09362_ (.A1(_01561_),
    .A2(_01548_),
    .B(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09363_ (.A1(_01558_),
    .A2(_01560_),
    .B1(_01563_),
    .B2(_01557_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09364_ (.A1(_01384_),
    .A2(_01492_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09365_ (.A1(_01384_),
    .A2(_01492_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09366_ (.A1(_01342_),
    .A2(net38),
    .B1(_01565_),
    .B2(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09367_ (.I(_01500_),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09368_ (.A1(_00573_),
    .A2(_07284_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09369_ (.A1(_01384_),
    .A2(_01500_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09370_ (.A1(_01568_),
    .A2(_01569_),
    .B(net13),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09371_ (.A1(net22),
    .A2(_01556_),
    .A3(_01567_),
    .A4(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09372_ (.A1(_01564_),
    .A2(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09373_ (.A1(_01551_),
    .A2(_01552_),
    .A3(_01572_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09374_ (.A1(_01437_),
    .A2(_01468_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09375_ (.A1(_01539_),
    .A2(_01573_),
    .B(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09376_ (.A1(_01311_),
    .A2(_01490_),
    .A3(_01521_),
    .A4(_01528_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _09377_ (.A1(_01551_),
    .A2(_01552_),
    .A3(_01572_),
    .B(_01576_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09378_ (.A1(_01532_),
    .A2(_01538_),
    .B(_01433_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09379_ (.A1(_01470_),
    .A2(_01529_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09380_ (.A1(_01577_),
    .A2(_01578_),
    .A3(_01579_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09381_ (.A1(_01531_),
    .A2(_01575_),
    .B(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09382_ (.A1(_01560_),
    .A2(_01563_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09383_ (.I(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09384_ (.A1(_01529_),
    .A2(_01552_),
    .B(_01551_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09385_ (.A1(_01583_),
    .A2(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09386_ (.A1(_01577_),
    .A2(_01578_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09387_ (.A1(_01471_),
    .A2(_01525_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09388_ (.A1(net22),
    .A2(_01516_),
    .A3(_01520_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09389_ (.A1(net22),
    .A2(_01587_),
    .B(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09390_ (.A1(_01489_),
    .A2(_01589_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09391_ (.A1(_01328_),
    .A2(_01397_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09392_ (.A1(_01425_),
    .A2(_01429_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09393_ (.A1(_01414_),
    .A2(_01483_),
    .A3(_01484_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09394_ (.I0(_01592_),
    .I1(_01593_),
    .S(net13),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09395_ (.A1(_01591_),
    .A2(_01536_),
    .B(_01534_),
    .C(_01594_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09396_ (.A1(_01311_),
    .A2(_01490_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09397_ (.A1(_01546_),
    .A2(_01550_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09398_ (.A1(_01437_),
    .A2(_01468_),
    .A3(_01469_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09399_ (.A1(_01564_),
    .A2(_01571_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _09400_ (.A1(_01596_),
    .A2(_01597_),
    .A3(_01598_),
    .A4(_01599_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09401_ (.A1(_01590_),
    .A2(_01595_),
    .B(_01600_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09402_ (.A1(_01491_),
    .A2(_01492_),
    .B(_01501_),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09403_ (.I0(_07301_),
    .I1(_01524_),
    .S(net22),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09404_ (.A1(_01384_),
    .A2(_01513_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09405_ (.A1(_01602_),
    .A2(_01603_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09406_ (.A1(_01515_),
    .A2(_01603_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09407_ (.A1(_01602_),
    .A2(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09408_ (.I0(_01604_),
    .I1(_01606_),
    .S(_01600_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09409_ (.I(_07359_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09410_ (.A1(_07342_),
    .A2(_07341_),
    .B(_07360_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09411_ (.A1(_01608_),
    .A2(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09412_ (.A1(_07357_),
    .A2(_01610_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09413_ (.A1(_01611_),
    .A2(_07356_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09414_ (.A1(_01612_),
    .A2(_07354_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09415_ (.A1(_01613_),
    .A2(_07353_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09416_ (.A1(_01614_),
    .A2(_07351_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09417_ (.A1(_01615_),
    .A2(_07350_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09418_ (.A1(_07348_),
    .A2(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09419_ (.A1(_01617_),
    .A2(_07347_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09420_ (.A1(_01618_),
    .A2(_07345_),
    .B(_07344_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09421_ (.A1(_01037_),
    .A2(_07220_),
    .ZN(_07233_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09422_ (.A1(_07235_),
    .A2(_00881_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09423_ (.I0(_07233_),
    .I1(_01620_),
    .S(_01233_),
    .Z(_07253_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09424_ (.A1(_07255_),
    .A2(_01022_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09425_ (.I0(_07253_),
    .I1(_01621_),
    .S(_01187_),
    .Z(_07270_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09426_ (.A1(_07272_),
    .A2(_01161_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09427_ (.I0(_07270_),
    .I1(_01622_),
    .S(_01381_),
    .Z(_07287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09428_ (.A1(_07289_),
    .A2(_01288_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09429_ (.I0(_07287_),
    .I1(_01623_),
    .S(_01491_),
    .Z(_07304_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09430_ (.A1(_07306_),
    .A2(_01408_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09431_ (.I0(_07304_),
    .I1(_01624_),
    .S(_01486_),
    .Z(_07321_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09432_ (.A1(_00574_),
    .A2(_07321_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _09433_ (.I(_00793_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09434_ (.A1(_01626_),
    .A2(_07321_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09435_ (.A1(_01619_),
    .A2(_01625_),
    .B(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09436_ (.A1(_07323_),
    .A2(_01512_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09437_ (.A1(_00573_),
    .A2(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09438_ (.A1(_00793_),
    .A2(_01629_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09439_ (.A1(_01619_),
    .A2(_01630_),
    .B(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09440_ (.A1(_01551_),
    .A2(_01529_),
    .A3(_01552_),
    .A4(_01572_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09441_ (.I0(_01628_),
    .I1(_01632_),
    .S(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09442_ (.A1(_01586_),
    .A2(_01601_),
    .A3(_01607_),
    .A4(_01634_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09443_ (.A1(_01581_),
    .A2(_01585_),
    .B(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09444_ (.A1(_01470_),
    .A2(_01577_),
    .B(_01579_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09445_ (.A1(_01636_),
    .A2(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09446_ (.A1(_01583_),
    .A2(_01584_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09447_ (.A1(_01467_),
    .A2(_01530_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09448_ (.A1(_01532_),
    .A2(_01538_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09449_ (.A1(_01597_),
    .A2(_01598_),
    .A3(_01599_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09450_ (.A1(_01641_),
    .A2(_01642_),
    .B(_01437_),
    .C(_01468_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09451_ (.A1(_01640_),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09452_ (.A1(_01577_),
    .A2(_01578_),
    .A3(_01579_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09453_ (.I(_01607_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09454_ (.I(_01634_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09455_ (.A1(_01645_),
    .A2(_01601_),
    .A3(_01646_),
    .A4(net30),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09456_ (.A1(_01644_),
    .A2(_01648_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09457_ (.A1(_01639_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09458_ (.A1(_01638_),
    .A2(_01650_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09459_ (.A1(_01384_),
    .A2(_01619_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09460_ (.I0(_07321_),
    .I1(_01629_),
    .S(_01633_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09461_ (.A1(_01601_),
    .A2(_01646_),
    .A3(_01652_),
    .A4(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09462_ (.A1(_00574_),
    .A2(_01619_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09463_ (.A1(_01653_),
    .A2(_01655_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09464_ (.A1(_01607_),
    .A2(_01647_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _09465_ (.A1(_01581_),
    .A2(_01585_),
    .A3(_01654_),
    .B1(_01656_),
    .B2(_01657_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09466_ (.A1(_01590_),
    .A2(_01595_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09467_ (.A1(_01531_),
    .A2(_01575_),
    .B1(_01600_),
    .B2(_01659_),
    .C(_01639_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09468_ (.A1(_01600_),
    .A2(_01590_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09469_ (.A1(_01646_),
    .A2(net30),
    .B(_01661_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09470_ (.A1(_01646_),
    .A2(net30),
    .A3(_01661_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09471_ (.A1(_01645_),
    .A2(_01660_),
    .B(_01662_),
    .C(_01663_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09472_ (.A1(_01658_),
    .A2(_01664_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09473_ (.A1(_01640_),
    .A2(_01643_),
    .B(_01585_),
    .C(_01601_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09474_ (.A1(_01646_),
    .A2(_01645_),
    .A3(_01647_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09475_ (.A1(_07345_),
    .A2(_01618_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09476_ (.I(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09477_ (.I(_01384_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09478_ (.I(_07373_),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09479_ (.I(_07362_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09480_ (.A1(_07365_),
    .A2(_07364_),
    .B(_07363_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09481_ (.A1(_01672_),
    .A2(_01673_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09482_ (.A1(_07380_),
    .A2(_01674_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09483_ (.A1(_01675_),
    .A2(_07379_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09484_ (.A1(_01676_),
    .A2(_07377_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09485_ (.A1(_01677_),
    .A2(_07376_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09486_ (.A1(_01678_),
    .A2(_07374_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09487_ (.A1(_01679_),
    .A2(_01671_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09488_ (.A1(_07368_),
    .A2(_01680_),
    .A3(_07371_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09489_ (.A1(_07368_),
    .A2(_07370_),
    .B(_07367_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09490_ (.A1(_01682_),
    .A2(_01681_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09491_ (.A1(_01683_),
    .A2(_01670_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09492_ (.A1(_01684_),
    .A2(_01586_),
    .A3(_01669_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09493_ (.A1(_01683_),
    .A2(_00574_),
    .B(_01281_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09494_ (.A1(_01668_),
    .A2(_01686_),
    .A3(_01586_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09495_ (.A1(_01666_),
    .A2(_01667_),
    .B1(_01687_),
    .B2(_01685_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09496_ (.A1(_01083_),
    .A2(_01040_),
    .B(_07237_),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09497_ (.A1(_07260_),
    .A2(_07258_),
    .A3(_07259_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09498_ (.A1(_01021_),
    .A2(_01689_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09499_ (.I0(_07256_),
    .I1(_01690_),
    .S(_01187_),
    .Z(_07261_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09500_ (.A1(_07263_),
    .A2(_01159_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09501_ (.I0(_07261_),
    .I1(_01691_),
    .S(_01381_),
    .Z(_07290_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09502_ (.A1(_07292_),
    .A2(_01286_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09503_ (.I0(_07290_),
    .I1(_01692_),
    .S(_01491_),
    .Z(_07307_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09504_ (.A1(_07311_),
    .A2(_01406_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09505_ (.A1(_07309_),
    .A2(_01693_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09506_ (.I0(_07307_),
    .I1(_01694_),
    .S(_01487_),
    .Z(_07324_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09507_ (.I(_07324_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09508_ (.A1(_07326_),
    .A2(_01510_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09509_ (.I0(_01695_),
    .I1(_01696_),
    .S(_01633_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09510_ (.A1(_01586_),
    .A2(_01697_),
    .A3(_01686_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09511_ (.I(_01697_),
    .ZN(_07343_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09512_ (.A1(_01586_),
    .A2(_07343_),
    .A3(_01684_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09513_ (.A1(_01645_),
    .A2(_01607_),
    .A3(_01634_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09514_ (.A1(_01698_),
    .A2(_01699_),
    .B(_01660_),
    .C(_01700_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09515_ (.A1(_01701_),
    .A2(_01688_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09516_ (.A1(_01640_),
    .A2(_01643_),
    .B(_01645_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09517_ (.A1(_01601_),
    .A2(_01646_),
    .A3(_01647_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09518_ (.A1(_01703_),
    .A2(_01639_),
    .B(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09519_ (.A1(_01311_),
    .A2(_01642_),
    .B(_01532_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09520_ (.A1(net13),
    .A2(_01592_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _09521_ (.A1(_01342_),
    .A2(net38),
    .B1(_01591_),
    .B2(_01420_),
    .C(_01593_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09522_ (.A1(_01516_),
    .A2(_01520_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09523_ (.A1(_01446_),
    .A2(_01477_),
    .A3(_01526_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09524_ (.A1(_01489_),
    .A2(net22),
    .A3(_01709_),
    .B(_01710_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09525_ (.A1(_01707_),
    .A2(_01708_),
    .A3(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09526_ (.A1(_01706_),
    .A2(_01712_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09527_ (.A1(_01600_),
    .A2(_01590_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09528_ (.A1(_01646_),
    .A2(_01647_),
    .A3(_01714_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09529_ (.A1(_01538_),
    .A2(_01706_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09530_ (.A1(_01713_),
    .A2(_01715_),
    .B(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _09531_ (.A1(_01646_),
    .A2(_01647_),
    .A3(_01714_),
    .B1(_01712_),
    .B2(_01706_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09532_ (.I(_01718_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09533_ (.A1(_01601_),
    .A2(_01713_),
    .A3(_01715_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09534_ (.A1(_01705_),
    .A2(_01717_),
    .A3(_01719_),
    .A4(_01720_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09535_ (.A1(_01665_),
    .A2(_01702_),
    .A3(_01721_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09536_ (.A1(_01668_),
    .A2(_01684_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09537_ (.A1(_01669_),
    .A2(_01686_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _09538_ (.A1(_01660_),
    .A2(_01700_),
    .B1(_01723_),
    .B2(_01724_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09539_ (.A1(_07343_),
    .A2(_01686_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09540_ (.A1(_01697_),
    .A2(_01684_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09541_ (.A1(_01726_),
    .A2(_01727_),
    .B(_01666_),
    .C(_01667_),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09542_ (.A1(_01725_),
    .A2(_01728_),
    .A3(_01658_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09543_ (.A1(_01651_),
    .A2(_01722_),
    .B(_01729_),
    .C(_01664_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09544_ (.A1(_01725_),
    .A2(_01728_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09545_ (.A1(_01660_),
    .A2(_01700_),
    .B(_01655_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09546_ (.A1(_01653_),
    .A2(_01732_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09547_ (.A1(_01646_),
    .A2(net30),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09548_ (.A1(_01580_),
    .A2(_01666_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09549_ (.A1(_01646_),
    .A2(net30),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09550_ (.A1(_01734_),
    .A2(_01735_),
    .B(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09551_ (.A1(_01731_),
    .A2(_01733_),
    .B(_01737_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09552_ (.A1(_01645_),
    .A2(_01660_),
    .B(_01715_),
    .C(_01713_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09553_ (.A1(_01718_),
    .A2(_01739_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09554_ (.A1(_01718_),
    .A2(_01739_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _09555_ (.A1(_01731_),
    .A2(_01665_),
    .A3(_01741_),
    .B1(_01717_),
    .B2(_01705_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09556_ (.A1(_01664_),
    .A2(_01729_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09557_ (.A1(_01740_),
    .A2(_01742_),
    .A3(_01743_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09558_ (.A1(_01730_),
    .A2(_01738_),
    .A3(_01744_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09559_ (.A1(_01638_),
    .A2(_01650_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09560_ (.A1(_01702_),
    .A2(_01665_),
    .A3(_01721_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09561_ (.I(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09562_ (.I(_07385_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09563_ (.A1(_07388_),
    .A2(_07387_),
    .B(_07386_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09564_ (.A1(_01750_),
    .A2(_01749_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09565_ (.A1(_07383_),
    .A2(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09566_ (.A1(_01752_),
    .A2(_07382_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09567_ (.A1(_07400_),
    .A2(_01753_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09568_ (.A1(_01754_),
    .A2(_07399_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09569_ (.A1(_07397_),
    .A2(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09570_ (.A1(_01756_),
    .A2(_07396_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09571_ (.A1(_07394_),
    .A2(_01757_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09572_ (.A1(_01758_),
    .A2(_07393_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09573_ (.A1(_01759_),
    .A2(_07391_),
    .B(_07390_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09574_ (.A1(_01670_),
    .A2(_01760_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09575_ (.A1(_01667_),
    .A2(_01666_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09576_ (.A1(_07348_),
    .A2(_01616_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09577_ (.A1(_07260_),
    .A2(_01198_),
    .ZN(_07264_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09578_ (.A1(_07266_),
    .A2(_07274_),
    .A3(_07273_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09579_ (.A1(_01158_),
    .A2(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09580_ (.I0(_07264_),
    .I1(_01765_),
    .S(_01381_),
    .Z(_07293_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09581_ (.A1(_07295_),
    .A2(_01284_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09582_ (.I0(_07293_),
    .I1(_01766_),
    .S(_01491_),
    .Z(_07310_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09583_ (.A1(_07312_),
    .A2(_01405_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09584_ (.I0(_07310_),
    .I1(_01767_),
    .S(_01487_),
    .Z(_07327_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09585_ (.A1(_07329_),
    .A2(_01508_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09586_ (.I0(_07327_),
    .I1(_01768_),
    .S(_01633_),
    .Z(_07346_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09587_ (.A1(_01666_),
    .A2(_01667_),
    .A3(_07346_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09588_ (.A1(_01762_),
    .A2(_01763_),
    .B(_01769_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09589_ (.A1(_01660_),
    .A2(_01700_),
    .B(_01668_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09590_ (.A1(_01660_),
    .A2(_01700_),
    .A3(_07343_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09591_ (.A1(_01771_),
    .A2(_01772_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09592_ (.A1(_01761_),
    .A2(_01770_),
    .B(_01773_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09593_ (.I(_01770_),
    .ZN(_07366_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09594_ (.A1(_01760_),
    .A2(_00574_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09595_ (.A1(_01775_),
    .A2(_01281_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09596_ (.A1(_07366_),
    .A2(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _09597_ (.A1(_01746_),
    .A2(_01748_),
    .A3(_01774_),
    .A4(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09598_ (.A1(_00574_),
    .A2(_01683_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09599_ (.I(_01779_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09600_ (.A1(_01771_),
    .A2(_01772_),
    .B(_01780_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09601_ (.A1(_01771_),
    .A2(_01772_),
    .A3(_01780_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09602_ (.A1(_07377_),
    .A2(_07379_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09603_ (.A1(_07376_),
    .A2(_01783_),
    .B(_07374_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09604_ (.A1(_01671_),
    .A2(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09605_ (.A1(_07371_),
    .A2(_07374_),
    .A3(_07377_),
    .A4(_07380_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _09606_ (.A1(_07371_),
    .A2(_01785_),
    .B1(_01786_),
    .B2(_01674_),
    .C(_07370_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09607_ (.A1(_07368_),
    .A2(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09608_ (.I0(_01761_),
    .I1(_01776_),
    .S(_01788_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09609_ (.A1(_01789_),
    .A2(_01782_),
    .A3(_01781_),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09610_ (.A1(_01731_),
    .A2(_01733_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09611_ (.A1(_01791_),
    .A2(_01790_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09612_ (.A1(_01792_),
    .A2(_01778_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09613_ (.A1(_01745_),
    .A2(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09614_ (.A1(_01665_),
    .A2(_01721_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09615_ (.A1(_01771_),
    .A2(_01772_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09616_ (.A1(_01670_),
    .A2(_01668_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09617_ (.A1(_00574_),
    .A2(_01669_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _09618_ (.A1(_01660_),
    .A2(_01700_),
    .B1(_01797_),
    .B2(_01798_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09619_ (.A1(_00574_),
    .A2(_07343_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09620_ (.A1(_01670_),
    .A2(_01697_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09621_ (.A1(_01800_),
    .A2(_01801_),
    .B(_01666_),
    .C(_01667_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09622_ (.A1(_01799_),
    .A2(_01802_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09623_ (.A1(_07368_),
    .A2(_07371_),
    .A3(_01680_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09624_ (.A1(_01804_),
    .A2(_01653_),
    .A3(_01655_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09625_ (.A1(_01666_),
    .A2(_01667_),
    .B(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09626_ (.A1(_01660_),
    .A2(_01700_),
    .A3(_01681_),
    .A4(_01653_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09627_ (.A1(_01681_),
    .A2(_01653_),
    .A3(_01655_),
    .B(_01682_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09628_ (.A1(_01806_),
    .A2(_01807_),
    .A3(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _09629_ (.A1(_01281_),
    .A2(_01796_),
    .B1(_01803_),
    .B2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09630_ (.A1(_01636_),
    .A2(_01637_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09631_ (.I(_01584_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09632_ (.A1(_01581_),
    .A2(_01704_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09633_ (.A1(_01437_),
    .A2(_01599_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09634_ (.A1(_01576_),
    .A2(_01598_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _09635_ (.A1(_01581_),
    .A2(_01583_),
    .A3(_01704_),
    .B1(_01814_),
    .B2(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09636_ (.A1(_01812_),
    .A2(_01813_),
    .B1(_01816_),
    .B2(_01597_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09637_ (.A1(_01531_),
    .A2(_01575_),
    .B(_01585_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09638_ (.I0(_01644_),
    .I1(_01818_),
    .S(_01648_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09639_ (.A1(_01586_),
    .A2(_01704_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09640_ (.A1(_01636_),
    .A2(_01819_),
    .A3(_01820_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09641_ (.A1(_01811_),
    .A2(_01817_),
    .A3(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09642_ (.A1(_01581_),
    .A2(_01704_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09643_ (.A1(_01551_),
    .A2(_01815_),
    .A3(_01814_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09644_ (.A1(_01582_),
    .A2(_01584_),
    .B(_01824_),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09645_ (.A1(_01823_),
    .A2(_01825_),
    .B(_01639_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09646_ (.A1(_07365_),
    .A2(_07368_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09647_ (.A1(_07363_),
    .A2(_01392_),
    .A3(_01786_),
    .A4(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09648_ (.A1(_01658_),
    .A2(_01799_),
    .A3(_01802_),
    .A4(_01828_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09649_ (.A1(_01826_),
    .A2(_01829_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09650_ (.A1(_01795_),
    .A2(_01810_),
    .A3(_01822_),
    .A4(_01830_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09651_ (.A1(_01815_),
    .A2(_01813_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09652_ (.A1(_01551_),
    .A2(_01832_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09653_ (.A1(_01582_),
    .A2(_01833_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09654_ (.A1(_07388_),
    .A2(_07394_),
    .A3(_07397_),
    .A4(_07400_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09655_ (.A1(_07386_),
    .A2(_07391_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09656_ (.A1(_07383_),
    .A2(_01392_),
    .A3(_01835_),
    .A4(_01836_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09657_ (.I(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09658_ (.A1(_01670_),
    .A2(_01770_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09659_ (.A1(_01838_),
    .A2(_01839_),
    .B(_01746_),
    .C(_01748_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09660_ (.A1(_01670_),
    .A2(_01788_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09661_ (.A1(_01837_),
    .A2(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09662_ (.A1(_01651_),
    .A2(_01722_),
    .B(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09663_ (.A1(_01831_),
    .A2(_01834_),
    .B1(_01840_),
    .B2(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09664_ (.A1(_01636_),
    .A2(_01820_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09665_ (.A1(_01795_),
    .A2(_01810_),
    .B(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09666_ (.A1(_01651_),
    .A2(_01748_),
    .B(_01638_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09667_ (.I0(_01832_),
    .I1(_01816_),
    .S(_01597_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09668_ (.A1(_01645_),
    .A2(_01704_),
    .A3(_01818_),
    .B(_01649_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09669_ (.A1(_01722_),
    .A2(_01848_),
    .B(_01849_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09670_ (.A1(_01702_),
    .A2(_01826_),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _09671_ (.A1(_01748_),
    .A2(_01848_),
    .B1(_01851_),
    .B2(_01795_),
    .C(_01819_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _09672_ (.A1(_01846_),
    .A2(_01847_),
    .A3(_01850_),
    .A4(_01852_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09673_ (.A1(_01844_),
    .A2(_01853_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09674_ (.A1(_07391_),
    .A2(_01759_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09675_ (.A1(_07403_),
    .A2(_07414_),
    .A3(_07417_),
    .A4(_07420_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09676_ (.A1(_07411_),
    .A2(_07406_),
    .A3(_07409_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09677_ (.A1(_01392_),
    .A2(_01856_),
    .A3(_01857_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09678_ (.A1(_01670_),
    .A2(_01858_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09679_ (.A1(_01846_),
    .A2(_01847_),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09680_ (.A1(_01855_),
    .A2(_01859_),
    .B(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09681_ (.A1(_01730_),
    .A2(_01738_),
    .A3(_01744_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09682_ (.A1(_01778_),
    .A2(_01792_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09683_ (.A1(_01855_),
    .A2(_01859_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09684_ (.A1(_01811_),
    .A2(_01650_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09685_ (.I0(_01811_),
    .I1(_01865_),
    .S(net27),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09686_ (.A1(_01864_),
    .A2(_01866_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09687_ (.A1(_01862_),
    .A2(_01863_),
    .B(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09688_ (.A1(_01794_),
    .A2(_01854_),
    .A3(_01861_),
    .B(_01868_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09689_ (.A1(_07391_),
    .A2(_01759_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09690_ (.A1(_00574_),
    .A2(_01858_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09691_ (.A1(_01870_),
    .A2(_01871_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09692_ (.A1(_01279_),
    .A2(_01277_),
    .B(_07274_),
    .ZN(_07296_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09693_ (.A1(_07300_),
    .A2(_07298_),
    .A3(_07299_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09694_ (.A1(_01283_),
    .A2(_01873_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09695_ (.I0(_07296_),
    .I1(_01874_),
    .S(_01491_),
    .Z(_07313_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09696_ (.A1(_07315_),
    .A2(_01403_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09697_ (.I0(_07313_),
    .I1(_01875_),
    .S(_01487_),
    .Z(_07330_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09698_ (.A1(_07332_),
    .A2(_01506_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09699_ (.I0(_07330_),
    .I1(_01876_),
    .S(_01633_),
    .Z(_07349_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09700_ (.A1(_07351_),
    .A2(_01614_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09701_ (.I0(_07349_),
    .I1(_01877_),
    .S(_01762_),
    .Z(_07369_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09702_ (.A1(_07371_),
    .A2(_01680_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09703_ (.A1(_01746_),
    .A2(_01747_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09704_ (.I0(_07369_),
    .I1(_01878_),
    .S(_01879_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09705_ (.I(_01880_),
    .Z(_07389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09706_ (.I0(_01859_),
    .I1(_01871_),
    .S(_07389_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _09707_ (.A1(_01745_),
    .A2(_01793_),
    .A3(_01844_),
    .A4(_01853_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09708_ (.I0(_01872_),
    .I1(_01881_),
    .S(_01882_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09709_ (.I0(_01817_),
    .I1(_01830_),
    .S(_01819_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09710_ (.A1(_01819_),
    .A2(_01817_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09711_ (.A1(_01665_),
    .A2(_01702_),
    .A3(_01721_),
    .A4(_01638_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09712_ (.I0(_01884_),
    .I1(_01885_),
    .S(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09713_ (.A1(_01746_),
    .A2(_01748_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09714_ (.A1(_01888_),
    .A2(_01790_),
    .B(_01778_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09715_ (.A1(_01651_),
    .A2(_01722_),
    .B(_01791_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09716_ (.A1(_01730_),
    .A2(_01738_),
    .A3(_01744_),
    .A4(_01890_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09717_ (.A1(_01889_),
    .A2(_01860_),
    .A3(_01891_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09718_ (.A1(_01844_),
    .A2(_01887_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09719_ (.A1(_01811_),
    .A2(_01821_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09720_ (.A1(_01795_),
    .A2(_01810_),
    .A3(_01894_),
    .B(_01848_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09721_ (.A1(_01831_),
    .A2(_01895_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09722_ (.A1(_01826_),
    .A2(_01829_),
    .B(_01819_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09723_ (.I0(_01897_),
    .I1(_01819_),
    .S(_01886_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09724_ (.A1(_01778_),
    .A2(_01792_),
    .B(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09725_ (.A1(_01745_),
    .A2(_01860_),
    .A3(_01896_),
    .A4(_01899_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09726_ (.A1(_01887_),
    .A2(_01892_),
    .B(_01893_),
    .C(_01900_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09727_ (.A1(_01831_),
    .A2(_01834_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09728_ (.A1(_01889_),
    .A2(_01860_),
    .A3(_01887_),
    .A4(_01891_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09729_ (.A1(_01638_),
    .A2(_01846_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _09730_ (.A1(_01902_),
    .A2(_01903_),
    .B1(_01904_),
    .B2(_01847_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09731_ (.A1(_01869_),
    .A2(_01883_),
    .A3(_01901_),
    .A4(_01905_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09732_ (.A1(_01745_),
    .A2(_01793_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09733_ (.A1(_01746_),
    .A2(net27),
    .B(_01788_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09734_ (.A1(_01746_),
    .A2(net27),
    .A3(_01770_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09735_ (.A1(_01908_),
    .A2(_01909_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09736_ (.A1(_01907_),
    .A2(_01854_),
    .A3(_01910_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09737_ (.A1(_01796_),
    .A2(_01909_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09738_ (.A1(_01888_),
    .A2(_01781_),
    .A3(_01782_),
    .A4(_01788_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09739_ (.I(_01670_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09740_ (.A1(_01912_),
    .A2(_01913_),
    .B(_01914_),
    .C(_01760_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09741_ (.A1(_00977_),
    .A2(_01760_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09742_ (.A1(_01670_),
    .A2(_01760_),
    .Z(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09743_ (.I0(_01916_),
    .I1(_01917_),
    .S(_01770_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09744_ (.I0(_01917_),
    .I1(_01916_),
    .S(_01788_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09745_ (.I0(_01918_),
    .I1(_01919_),
    .S(_01879_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09746_ (.A1(_01281_),
    .A2(_01775_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09747_ (.A1(_01670_),
    .A2(_01760_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09748_ (.A1(_01921_),
    .A2(_01908_),
    .A3(_01909_),
    .A4(_01922_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09749_ (.A1(_01746_),
    .A2(net27),
    .B(_01780_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09750_ (.A1(_01773_),
    .A2(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09751_ (.I0(_01920_),
    .I1(_01923_),
    .S(_01925_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09752_ (.A1(_01915_),
    .A2(_01926_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _09753_ (.A1(_01793_),
    .A2(_01745_),
    .A3(_01844_),
    .A4(_01853_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09754_ (.A1(_01725_),
    .A2(_01728_),
    .A3(_01658_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09755_ (.A1(_01781_),
    .A2(_01782_),
    .A3(_01789_),
    .B(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09756_ (.I0(_01790_),
    .I1(_01930_),
    .S(_01738_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09757_ (.A1(_01791_),
    .A2(_01931_),
    .B(_01879_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09758_ (.A1(_01778_),
    .A2(_01932_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09759_ (.A1(_01928_),
    .A2(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09760_ (.A1(_01844_),
    .A2(_01853_),
    .A3(_01891_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09761_ (.A1(_01730_),
    .A2(_01743_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09762_ (.A1(_01653_),
    .A2(_01732_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09763_ (.A1(_01799_),
    .A2(_01802_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09764_ (.A1(_01806_),
    .A2(_01807_),
    .A3(_01808_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09765_ (.A1(_01626_),
    .A2(_01773_),
    .B1(_01938_),
    .B2(_01939_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09766_ (.A1(_01734_),
    .A2(_01735_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09767_ (.A1(_01937_),
    .A2(_01940_),
    .B1(_01941_),
    .B2(_01736_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09768_ (.A1(_01778_),
    .A2(_01792_),
    .B(_01942_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09769_ (.A1(_01936_),
    .A2(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09770_ (.A1(_01741_),
    .A2(_01730_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09771_ (.A1(_01935_),
    .A2(_01944_),
    .B(_01945_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09772_ (.A1(_01911_),
    .A2(_01927_),
    .B(_01934_),
    .C(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09773_ (.A1(_01651_),
    .A2(net27),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09774_ (.A1(_01846_),
    .A2(_01948_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09775_ (.A1(_01844_),
    .A2(_01853_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09776_ (.A1(_01740_),
    .A2(_01730_),
    .A3(_01743_),
    .A4(_01738_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09777_ (.A1(_01665_),
    .A2(_01702_),
    .A3(_01651_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09778_ (.A1(_01795_),
    .A2(_01810_),
    .A3(_01952_),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09779_ (.A1(_01951_),
    .A2(_01793_),
    .B1(_01953_),
    .B2(_01742_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09780_ (.A1(_01907_),
    .A2(_01950_),
    .B(_01954_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09781_ (.A1(_01949_),
    .A2(_01955_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09782_ (.I(_07408_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09783_ (.A1(_07411_),
    .A2(_07410_),
    .B(_07409_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09784_ (.A1(_01957_),
    .A2(_01958_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09785_ (.A1(_01959_),
    .A2(_07406_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09786_ (.A1(_01960_),
    .A2(_07405_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09787_ (.A1(_07403_),
    .A2(_01961_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09788_ (.A1(_01962_),
    .A2(_07402_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09789_ (.A1(_07420_),
    .A2(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09790_ (.A1(_07419_),
    .A2(_01964_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09791_ (.A1(_07417_),
    .A2(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09792_ (.A1(_01966_),
    .A2(_07416_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09793_ (.A1(_07414_),
    .A2(_01967_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09794_ (.A1(_07413_),
    .A2(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09795_ (.A1(_01914_),
    .A2(_07389_),
    .A3(_01969_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09796_ (.A1(_01914_),
    .A2(_01870_),
    .A3(_01969_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09797_ (.I0(_01970_),
    .I1(_01971_),
    .S(_01928_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09798_ (.A1(_07413_),
    .A2(_01968_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09799_ (.A1(_01914_),
    .A2(_01973_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09800_ (.A1(_01974_),
    .A2(_07389_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09801_ (.A1(_01870_),
    .A2(_01974_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09802_ (.I0(_01975_),
    .I1(_01976_),
    .S(_01928_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09803_ (.A1(_01626_),
    .A2(_01870_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09804_ (.A1(_01626_),
    .A2(_07389_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09805_ (.I0(_01978_),
    .I1(_01979_),
    .S(_01882_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09806_ (.A1(_01972_),
    .A2(_01980_),
    .A3(_01977_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09807_ (.A1(_01981_),
    .A2(_01947_),
    .A3(_01956_),
    .A4(_01906_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _09808_ (.I(_01982_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09809_ (.A1(_07411_),
    .A2(_01983_),
    .ZN(_07430_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09810_ (.A1(_07434_),
    .A2(_07433_),
    .B(_07432_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09811_ (.A1(_07434_),
    .A2(_07432_),
    .A3(_07433_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09812_ (.A1(_01984_),
    .A2(_01985_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09813_ (.A1(_01906_),
    .A2(_01947_),
    .A3(_01956_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09814_ (.A1(_01936_),
    .A2(_01943_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09815_ (.I(_01928_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09816_ (.A1(_01933_),
    .A2(_01988_),
    .B(net17),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09817_ (.A1(_01911_),
    .A2(_01927_),
    .B(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09818_ (.I(_01945_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09819_ (.A1(_01936_),
    .A2(_01943_),
    .B(_01992_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09820_ (.A1(_01936_),
    .A2(_01935_),
    .A3(_01943_),
    .A4(_01992_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09821_ (.A1(_01742_),
    .A2(_01953_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09822_ (.A1(_01951_),
    .A2(_01793_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09823_ (.A1(_01846_),
    .A2(_01948_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09824_ (.A1(_01745_),
    .A2(_01793_),
    .B(_01997_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _09825_ (.A1(_01995_),
    .A2(_01996_),
    .B1(_01998_),
    .B2(_01854_),
    .C(_01866_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09826_ (.A1(_01993_),
    .A2(_01994_),
    .A3(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09827_ (.A1(net20),
    .A2(_01991_),
    .A3(_02000_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09828_ (.A1(_01831_),
    .A2(_01895_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09829_ (.A1(_01844_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09830_ (.A1(_01889_),
    .A2(_01860_),
    .A3(_01891_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09831_ (.A1(_01898_),
    .A2(_02004_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09832_ (.I0(_02002_),
    .I1(_02003_),
    .S(_02005_),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09833_ (.A1(_01987_),
    .A2(_02001_),
    .B(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09834_ (.A1(_01987_),
    .A2(_02006_),
    .A3(_02001_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09835_ (.A1(_01908_),
    .A2(_01909_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09836_ (.A1(_01794_),
    .A2(_01950_),
    .A3(_02009_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09837_ (.A1(_01915_),
    .A2(_01926_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09838_ (.A1(_02010_),
    .A2(_02011_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09839_ (.A1(_01972_),
    .A2(_01977_),
    .A3(_01980_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09840_ (.A1(_01890_),
    .A2(_02012_),
    .A3(_02013_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09841_ (.A1(_01738_),
    .A2(_01935_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09842_ (.A1(_01879_),
    .A2(_01729_),
    .B(_01942_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09843_ (.I0(_02015_),
    .I1(_02016_),
    .S(_01863_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09844_ (.A1(_01889_),
    .A2(_01890_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09845_ (.A1(_01793_),
    .A2(_01935_),
    .B(_02018_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09846_ (.A1(_02017_),
    .A2(_02019_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09847_ (.A1(_01987_),
    .A2(_02014_),
    .B(_02020_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09848_ (.A1(_01993_),
    .A2(_01994_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09849_ (.A1(_01911_),
    .A2(_01927_),
    .B(_01934_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09850_ (.A1(_02023_),
    .A2(net20),
    .B(_01944_),
    .C(_01935_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09851_ (.A1(_01955_),
    .A2(_02022_),
    .A3(_02024_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09852_ (.A1(_02007_),
    .A2(_02008_),
    .B(_02021_),
    .C(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09853_ (.A1(_01902_),
    .A2(_01903_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09854_ (.A1(_01898_),
    .A2(_02004_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09855_ (.A1(_01950_),
    .A2(_02005_),
    .B(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09856_ (.A1(_01901_),
    .A2(_01981_),
    .A3(_01991_),
    .A4(_02000_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09857_ (.A1(_02027_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_01987_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09858_ (.A1(_02009_),
    .A2(_01922_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09859_ (.A1(_01870_),
    .A2(_01882_),
    .A3(_02032_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _09860_ (.A1(net17),
    .A2(_07389_),
    .A3(_02009_),
    .B(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09861_ (.A1(_01914_),
    .A2(_01969_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09862_ (.A1(_00758_),
    .A2(_01973_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09863_ (.A1(_01980_),
    .A2(_02035_),
    .B(_02036_),
    .C(_01972_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09864_ (.A1(_02013_),
    .A2(_02034_),
    .Z(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09865_ (.A1(_01869_),
    .A2(_01883_),
    .A3(_01901_),
    .A4(_01905_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09866_ (.A1(_01844_),
    .A2(_01853_),
    .A3(_01891_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09867_ (.A1(_01936_),
    .A2(_01943_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09868_ (.A1(_02040_),
    .A2(_02041_),
    .B(_01992_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _09869_ (.A1(_02010_),
    .A2(_02011_),
    .B1(_01933_),
    .B2(net17),
    .C(_02042_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _09870_ (.A1(_01949_),
    .A2(_02039_),
    .A3(_02043_),
    .A4(_01955_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09871_ (.I(_07389_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09872_ (.I0(_01855_),
    .I1(_02045_),
    .S(_01882_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09873_ (.A1(_00575_),
    .A2(_01969_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09874_ (.I(_01922_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09875_ (.A1(_01928_),
    .A2(_02048_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09876_ (.A1(_01281_),
    .A2(_01910_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09877_ (.A1(_02049_),
    .A2(_02050_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09878_ (.A1(_01914_),
    .A2(_01969_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09879_ (.A1(_07389_),
    .A2(_01910_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09880_ (.A1(_01855_),
    .A2(_02048_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09881_ (.A1(_01855_),
    .A2(_01922_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09882_ (.I0(_02054_),
    .I1(_02055_),
    .S(_02009_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09883_ (.I0(_02053_),
    .I1(_02056_),
    .S(net17),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09884_ (.A1(_07389_),
    .A2(_01910_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09885_ (.A1(_01870_),
    .A2(_02048_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09886_ (.A1(_01870_),
    .A2(_01922_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09887_ (.I0(_02059_),
    .I1(_02060_),
    .S(_01910_),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09888_ (.I0(_02058_),
    .I1(_02061_),
    .S(net17),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09889_ (.A1(_02052_),
    .A2(_02057_),
    .B1(_02062_),
    .B2(_01974_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09890_ (.A1(_02046_),
    .A2(_02047_),
    .A3(_02051_),
    .B(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _09891_ (.A1(_02034_),
    .A2(_02037_),
    .B1(_02038_),
    .B2(_02044_),
    .C(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09892_ (.A1(_01981_),
    .A2(_01991_),
    .A3(_02000_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09893_ (.A1(_01907_),
    .A2(_01949_),
    .A3(_01950_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09894_ (.A1(_01866_),
    .A2(_02067_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09895_ (.A1(_02039_),
    .A2(_01991_),
    .A3(_02000_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09896_ (.A1(_01949_),
    .A2(_02043_),
    .A3(_01955_),
    .A4(_02013_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09897_ (.A1(_02066_),
    .A2(_02068_),
    .B1(_02069_),
    .B2(_02070_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09898_ (.A1(_02039_),
    .A2(_01947_),
    .A3(_01956_),
    .A4(net20),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09899_ (.A1(_01907_),
    .A2(_01949_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09900_ (.A1(_01950_),
    .A2(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09901_ (.A1(_07413_),
    .A2(_01911_),
    .A3(_01927_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09902_ (.A1(_01972_),
    .A2(_01977_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09903_ (.I0(_02075_),
    .I1(_01997_),
    .S(_02076_),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09904_ (.A1(_02043_),
    .A2(_01955_),
    .A3(_01980_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09905_ (.A1(_02072_),
    .A2(_02074_),
    .B1(_02077_),
    .B2(_02078_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09906_ (.A1(_02031_),
    .A2(_02065_),
    .A3(_02071_),
    .A4(_02079_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09907_ (.A1(_02012_),
    .A2(_02013_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09908_ (.A1(_02009_),
    .A2(_02049_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09909_ (.I0(_01761_),
    .I1(_01776_),
    .S(_02009_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09910_ (.A1(_01796_),
    .A2(_01924_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09911_ (.A1(_01889_),
    .A2(_01935_),
    .B1(_02083_),
    .B2(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09912_ (.A1(_02082_),
    .A2(_02013_),
    .B(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09913_ (.A1(_01987_),
    .A2(_02081_),
    .B(_02086_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _09914_ (.A1(_07414_),
    .A2(_01967_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09915_ (.A1(_01342_),
    .A2(_01344_),
    .B(_07300_),
    .ZN(_07316_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09916_ (.A1(_07320_),
    .A2(_07318_),
    .A3(_07319_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09917_ (.A1(_01402_),
    .A2(_02089_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09918_ (.I0(_07316_),
    .I1(_02090_),
    .S(_01487_),
    .Z(_07333_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09919_ (.A1(_07335_),
    .A2(_01504_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09920_ (.I0(_07333_),
    .I1(_02091_),
    .S(_01633_),
    .Z(_07352_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09921_ (.A1(_07354_),
    .A2(_01612_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09922_ (.I0(_07352_),
    .I1(_02092_),
    .S(_01762_),
    .Z(_07372_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09923_ (.A1(_07374_),
    .A2(_01678_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09924_ (.I0(_07372_),
    .I1(_02093_),
    .S(_01879_),
    .Z(_07392_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09925_ (.I(_07392_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09926_ (.A1(_07394_),
    .A2(_01757_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09927_ (.I0(_02094_),
    .I1(_02095_),
    .S(_01989_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09928_ (.A1(_02039_),
    .A2(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09929_ (.A1(_01947_),
    .A2(_01956_),
    .A3(_01981_),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09930_ (.A1(_01983_),
    .A2(_02088_),
    .B1(_02097_),
    .B2(_02098_),
    .C(_01626_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09931_ (.A1(_07414_),
    .A2(_01967_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09932_ (.I(_07439_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09933_ (.I(_07431_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09934_ (.A1(_01984_),
    .A2(_02102_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09935_ (.A1(_07429_),
    .A2(_02103_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09936_ (.A1(_02104_),
    .A2(_07428_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09937_ (.A1(_02105_),
    .A2(_07426_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09938_ (.A1(_02106_),
    .A2(_07425_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09939_ (.A1(_02107_),
    .A2(_07423_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09940_ (.A1(_02108_),
    .A2(_07422_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09941_ (.A1(_02109_),
    .A2(_07440_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09942_ (.A1(_02101_),
    .A2(_02110_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09943_ (.A1(_02111_),
    .A2(_07437_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09944_ (.A1(_02112_),
    .A2(_07436_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09945_ (.A1(_00574_),
    .A2(_02113_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09946_ (.A1(_02114_),
    .A2(_02100_),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09947_ (.A1(_02114_),
    .A2(_02096_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09948_ (.I0(_02115_),
    .I1(_02116_),
    .S(_01982_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09949_ (.A1(_01914_),
    .A2(_02113_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09950_ (.A1(_01982_),
    .A2(_02088_),
    .B1(_02097_),
    .B2(_02098_),
    .C(_02118_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _09951_ (.A1(_02087_),
    .A2(_02099_),
    .A3(_02119_),
    .A4(_02117_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09952_ (.A1(_02120_),
    .A2(_02080_),
    .A3(_02026_),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 clone40 (.A1(_02120_),
    .A2(_02080_),
    .A3(_02026_),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09954_ (.I0(_07430_),
    .I1(_01986_),
    .S(_02121_),
    .Z(_07450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09955_ (.I(_07454_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09956_ (.A1(_07457_),
    .A2(_07456_),
    .B(_07455_),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09957_ (.A1(_02123_),
    .A2(_02124_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09958_ (.A1(_07452_),
    .A2(_02125_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09959_ (.I(_02026_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _09960_ (.I(_02080_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09961_ (.A1(_02087_),
    .A2(_02099_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _09962_ (.I(_01914_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09963_ (.I0(_02100_),
    .I1(_02096_),
    .S(net9),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09964_ (.A1(_02130_),
    .A2(_02131_),
    .A3(_02113_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09965_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02129_),
    .B(_02132_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09966_ (.A1(_01866_),
    .A2(_02067_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _09967_ (.A1(_02039_),
    .A2(_01991_),
    .A3(_02000_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _09968_ (.A1(_02001_),
    .A2(_02134_),
    .B1(_02135_),
    .B2(_02098_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09969_ (.I(_01955_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09970_ (.A1(_02076_),
    .A2(_02075_),
    .B(_01980_),
    .C(_02043_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09971_ (.A1(_01949_),
    .A2(_02013_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _09972_ (.A1(_02039_),
    .A2(_01947_),
    .A3(_01956_),
    .A4(net20),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09973_ (.A1(_01950_),
    .A2(_02073_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _09974_ (.A1(_02137_),
    .A2(_02138_),
    .A3(_02139_),
    .B1(_02140_),
    .B2(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09975_ (.A1(_02136_),
    .A2(_02142_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _09976_ (.I(_02006_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09977_ (.A1(_02044_),
    .A2(_02066_),
    .B(_02144_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09978_ (.A1(_02044_),
    .A2(_02144_),
    .A3(_02066_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09979_ (.A1(_01890_),
    .A2(_02012_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _09980_ (.A1(_01906_),
    .A2(_01947_),
    .A3(_01956_),
    .B(_02013_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09981_ (.A1(_01955_),
    .A2(_02022_),
    .A3(_02017_),
    .A4(_02019_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09982_ (.A1(_02147_),
    .A2(_02148_),
    .B(_02024_),
    .C(_02149_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09983_ (.I(_02029_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _09984_ (.A1(_02145_),
    .A2(_02146_),
    .B(_02150_),
    .C(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09985_ (.A1(_02013_),
    .A2(_02034_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09986_ (.A1(_02046_),
    .A2(_02047_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09987_ (.A1(_02049_),
    .A2(_02050_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _09988_ (.A1(_02154_),
    .A2(_02155_),
    .B1(_02057_),
    .B2(_02052_),
    .C1(_01974_),
    .C2(_02062_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09989_ (.A1(_02034_),
    .A2(_02037_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09990_ (.A1(_01987_),
    .A2(_02153_),
    .B(_02156_),
    .C(_02157_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09991_ (.A1(_02158_),
    .A2(_02087_),
    .A3(_02099_),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09992_ (.A1(_01902_),
    .A2(_01903_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09993_ (.I(_02096_),
    .ZN(_07412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _09994_ (.I0(_02088_),
    .I1(_07412_),
    .S(_01983_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09995_ (.A1(_01981_),
    .A2(_01947_),
    .A3(_01956_),
    .A4(_01906_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09996_ (.A1(_02162_),
    .A2(_02030_),
    .A3(_02100_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09997_ (.A1(_02160_),
    .A2(_02161_),
    .B(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _09998_ (.A1(_02143_),
    .A2(_02152_),
    .A3(_02159_),
    .A4(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09999_ (.A1(_02161_),
    .A2(_02113_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10000_ (.A1(_02100_),
    .A2(_02114_),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10001_ (.A1(_02096_),
    .A2(_02114_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10002_ (.I0(_02167_),
    .I1(_02168_),
    .S(_01983_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10003_ (.A1(_02130_),
    .A2(_02166_),
    .B(_02169_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10004_ (.A1(_02133_),
    .A2(_02165_),
    .A3(_02170_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10005_ (.I(_07451_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10006_ (.A1(_07455_),
    .A2(_07456_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10007_ (.A1(_07454_),
    .A2(_02173_),
    .B(_07452_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10008_ (.A1(_02172_),
    .A2(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10009_ (.A1(_07449_),
    .A2(_07452_),
    .A3(_07455_),
    .A4(_07457_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10010_ (.A1(_07449_),
    .A2(_02175_),
    .B(_07448_),
    .C(_02176_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10011_ (.I(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10012_ (.A1(_02178_),
    .A2(_07446_),
    .B(_07445_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10013_ (.I(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10014_ (.A1(_07443_),
    .A2(_02180_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10015_ (.A1(_02181_),
    .A2(_07442_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10016_ (.A1(_02182_),
    .A2(_07460_),
    .B(_07459_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _10017_ (.I(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10018_ (.A1(_02184_),
    .A2(_00575_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10019_ (.A1(_02184_),
    .A2(_01914_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10020_ (.A1(_01446_),
    .A2(_07320_),
    .ZN(_07336_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10021_ (.A1(_07338_),
    .A2(_07340_),
    .A3(_07339_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10022_ (.A1(_01503_),
    .A2(_02187_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10023_ (.I0(_07336_),
    .I1(_02188_),
    .S(_01633_),
    .Z(_07355_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10024_ (.A1(_07357_),
    .A2(_01610_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10025_ (.I0(_07355_),
    .I1(_02189_),
    .S(_01762_),
    .Z(_07375_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10026_ (.A1(_07377_),
    .A2(_01676_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10027_ (.I0(_07375_),
    .I1(_02190_),
    .S(_01879_),
    .Z(_07395_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10028_ (.A1(_07397_),
    .A2(_01755_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10029_ (.I0(_07395_),
    .I1(_02191_),
    .S(_01989_),
    .Z(_07415_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10030_ (.A1(_07417_),
    .A2(_01965_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10031_ (.I0(_07415_),
    .I1(_02192_),
    .S(_02162_),
    .Z(_07435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10032_ (.I0(_02185_),
    .I1(_02186_),
    .S(_07435_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10033_ (.A1(_01626_),
    .A2(_07435_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10034_ (.A1(_02193_),
    .A2(_02194_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10035_ (.I(_01281_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10036_ (.A1(_07437_),
    .A2(_02111_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10037_ (.I0(_02186_),
    .I1(_02185_),
    .S(_02197_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10038_ (.A1(_02196_),
    .A2(_02197_),
    .B(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _10039_ (.I0(_02195_),
    .I1(_02199_),
    .S(_02121_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10040_ (.A1(_02200_),
    .A2(_02171_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10041_ (.I(_02201_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10042_ (.A1(_01626_),
    .A2(_02118_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10043_ (.A1(_02088_),
    .A2(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10044_ (.A1(_07412_),
    .A2(_02203_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10045_ (.I0(_02204_),
    .I1(_02205_),
    .S(_01982_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10046_ (.A1(_02158_),
    .A2(_02087_),
    .A3(_02117_),
    .A4(_02206_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10047_ (.A1(_02127_),
    .A2(_02080_),
    .B(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10048_ (.I(_02019_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10049_ (.A1(_01987_),
    .A2(_02081_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10050_ (.A1(_01987_),
    .A2(_02014_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10051_ (.A1(_02209_),
    .A2(_02210_),
    .B(_02211_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _10052_ (.A1(_02208_),
    .A2(_02212_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10053_ (.I(_01974_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10054_ (.A1(_02214_),
    .A2(_02047_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10055_ (.A1(net9),
    .A2(_02215_),
    .B(_02046_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10056_ (.A1(_02046_),
    .A2(net9),
    .A3(_02215_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _10057_ (.A1(_02161_),
    .A2(_02203_),
    .B1(_02216_),
    .B2(_02217_),
    .C(_02169_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10058_ (.A1(_02127_),
    .A2(_02128_),
    .B(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10059_ (.I(_02215_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10060_ (.A1(_02162_),
    .A2(_02220_),
    .B(_02046_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10061_ (.A1(_02046_),
    .A2(_02162_),
    .A3(_02220_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10062_ (.A1(_02087_),
    .A2(_02221_),
    .A3(_02222_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10063_ (.A1(_02216_),
    .A2(_02217_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10064_ (.A1(_02117_),
    .A2(_02206_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10065_ (.I0(_02223_),
    .I1(_02224_),
    .S(_02225_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10066_ (.A1(_02082_),
    .A2(_02148_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10067_ (.A1(_02218_),
    .A2(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10068_ (.A1(_02012_),
    .A2(_02013_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10069_ (.A1(_02085_),
    .A2(_02013_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _10070_ (.A1(_02085_),
    .A2(_02082_),
    .B1(_02044_),
    .B2(_02229_),
    .C(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10071_ (.A1(_02158_),
    .A2(_02117_),
    .A3(_02206_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10072_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02231_),
    .B(_02232_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10073_ (.A1(_02219_),
    .A2(_02226_),
    .A3(_02228_),
    .A4(_02233_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10074_ (.A1(_02031_),
    .A2(_02065_),
    .A3(_02071_),
    .A4(_02079_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10075_ (.A1(_02145_),
    .A2(_02146_),
    .B(_02150_),
    .C(_02231_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10076_ (.A1(_02235_),
    .A2(_02236_),
    .B(_02225_),
    .C(_02065_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _10077_ (.A1(_02231_),
    .A2(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _10078_ (.A1(_02213_),
    .A2(_02234_),
    .A3(_02238_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10079_ (.A1(_02145_),
    .A2(_02146_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10080_ (.A1(_02021_),
    .A2(_02025_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10081_ (.A1(_02240_),
    .A2(_02128_),
    .B(_02207_),
    .C(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10082_ (.A1(_01987_),
    .A2(_02001_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10083_ (.I(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10084_ (.A1(_02244_),
    .A2(_02029_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10085_ (.A1(_02144_),
    .A2(_02143_),
    .A3(_02242_),
    .A4(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10086_ (.A1(_02130_),
    .A2(_07435_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10087_ (.A1(_07443_),
    .A2(_07446_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10088_ (.A1(_07460_),
    .A2(_01392_),
    .A3(_02176_),
    .A4(_02248_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10089_ (.A1(_02247_),
    .A2(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10090_ (.A1(_00575_),
    .A2(_02249_),
    .A3(_02197_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10091_ (.A1(_02143_),
    .A2(_02152_),
    .A3(_02207_),
    .A4(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10092_ (.A1(_01901_),
    .A2(_01991_),
    .A3(_02000_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10093_ (.A1(_02148_),
    .A2(_02253_),
    .B(_02160_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10094_ (.A1(_02254_),
    .A2(_02251_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10095_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02120_),
    .B(_02255_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10096_ (.A1(_07437_),
    .A2(_02111_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10097_ (.A1(_02130_),
    .A2(_02249_),
    .A3(_02257_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10098_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02120_),
    .B(_02258_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _10099_ (.A1(net40),
    .A2(_02250_),
    .B1(_02252_),
    .B2(_02256_),
    .C(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10100_ (.A1(_01987_),
    .A2(_02138_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10101_ (.A1(_02022_),
    .A2(_02138_),
    .B(_01983_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10102_ (.A1(net20),
    .A2(_01991_),
    .A3(_02261_),
    .B(_02262_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10103_ (.A1(_01955_),
    .A2(_02263_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10104_ (.A1(_02242_),
    .A2(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _10105_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02120_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10106_ (.A1(_01991_),
    .A2(_02148_),
    .B(_02024_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10107_ (.A1(_02021_),
    .A2(_02207_),
    .B(_02267_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10108_ (.A1(_02017_),
    .A2(_02209_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10109_ (.A1(_02161_),
    .A2(_02118_),
    .B(_02269_),
    .C(_02169_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10110_ (.A1(_02159_),
    .A2(_02270_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10111_ (.A1(_02211_),
    .A2(_02017_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _10112_ (.A1(_02266_),
    .A2(_02268_),
    .B1(_02271_),
    .B2(_02272_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10113_ (.A1(_02246_),
    .A2(_02260_),
    .A3(_02265_),
    .A4(_02273_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _10114_ (.A1(_02274_),
    .A2(_02239_),
    .A3(_02202_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10115_ (.I(_02275_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10116_ (.I0(_07450_),
    .I1(_02126_),
    .S(_02276_),
    .Z(_07470_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10117_ (.I(_07477_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10118_ (.A1(_07480_),
    .A2(_07479_),
    .B(_07478_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10119_ (.A1(_02277_),
    .A2(_02278_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10120_ (.A1(_07475_),
    .A2(_02279_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10121_ (.A1(_07474_),
    .A2(_02280_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10122_ (.A1(_07472_),
    .A2(_02281_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10123_ (.A1(_02133_),
    .A2(_02165_),
    .A3(_02170_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10124_ (.A1(_02193_),
    .A2(_02194_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10125_ (.A1(_02130_),
    .A2(_02184_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10126_ (.A1(_02196_),
    .A2(_02257_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10127_ (.A1(_02285_),
    .A2(_02227_),
    .B(_02286_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10128_ (.A1(_02197_),
    .A2(_02185_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10129_ (.A1(_02088_),
    .A2(_02113_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10130_ (.A1(_07412_),
    .A2(_02113_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10131_ (.I0(_02289_),
    .I1(_02290_),
    .S(net9),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _10132_ (.A1(_02216_),
    .A2(_02217_),
    .B(_02291_),
    .C(_02286_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10133_ (.A1(_02196_),
    .A2(_02257_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10134_ (.A1(_02216_),
    .A2(_02217_),
    .A3(_02291_),
    .A4(_02293_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10135_ (.A1(_02287_),
    .A2(_02288_),
    .A3(_02292_),
    .A4(_02294_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10136_ (.I0(_02284_),
    .I1(_02295_),
    .S(net40),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10137_ (.A1(_02283_),
    .A2(_02234_),
    .A3(_02238_),
    .A4(_02296_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10138_ (.A1(_02087_),
    .A2(_02232_),
    .B(_02208_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10139_ (.A1(_02283_),
    .A2(_02234_),
    .A3(_02296_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10140_ (.A1(_02298_),
    .A2(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10141_ (.A1(_02171_),
    .A2(_02200_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10142_ (.A1(_02213_),
    .A2(_02234_),
    .A3(_02238_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10143_ (.A1(_02246_),
    .A2(_02260_),
    .A3(_02265_),
    .A4(_02273_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _10144_ (.A1(_02301_),
    .A2(_02302_),
    .A3(_02303_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10145_ (.A1(_02158_),
    .A2(_02087_),
    .A3(_02117_),
    .A4(_02206_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10146_ (.I(_02267_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10147_ (.A1(_02211_),
    .A2(_02020_),
    .A3(_02305_),
    .B(_02306_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10148_ (.A1(_02159_),
    .A2(_02270_),
    .B(_02272_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10149_ (.A1(net40),
    .A2(_02307_),
    .B(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _10150_ (.A1(_02213_),
    .A2(_02297_),
    .B1(_02300_),
    .B2(_02304_),
    .C(_02309_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _10151_ (.I(_02239_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10152_ (.I0(_07435_),
    .I1(_02257_),
    .S(net40),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10153_ (.A1(_01576_),
    .A2(_01642_),
    .B(_07340_),
    .ZN(_07358_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10154_ (.A1(_07360_),
    .A2(_07342_),
    .A3(_07341_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10155_ (.A1(_01609_),
    .A2(_02313_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10156_ (.I0(_07358_),
    .I1(_02314_),
    .S(_01762_),
    .Z(_07378_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10157_ (.A1(_07380_),
    .A2(_01674_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10158_ (.I0(_07378_),
    .I1(_02315_),
    .S(_01879_),
    .Z(_07398_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10159_ (.A1(_07400_),
    .A2(_01753_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10160_ (.I0(_07398_),
    .I1(_02316_),
    .S(_01989_),
    .Z(_07418_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10161_ (.I(_07418_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10162_ (.A1(_07420_),
    .A2(_01963_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10163_ (.I0(_02317_),
    .I1(_02318_),
    .S(_02162_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10164_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02120_),
    .A4(_02319_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10165_ (.A1(_07440_),
    .A2(_02109_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10166_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02120_),
    .B(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10167_ (.A1(_07472_),
    .A2(_02281_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10168_ (.A1(_02323_),
    .A2(_07471_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10169_ (.A1(_07469_),
    .A2(_02324_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10170_ (.A1(_02325_),
    .A2(_07468_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10171_ (.A1(_07466_),
    .A2(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10172_ (.A1(_02327_),
    .A2(_07465_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10173_ (.A1(_02328_),
    .A2(_07463_),
    .B(_07462_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _10174_ (.I(_02329_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10175_ (.A1(_02330_),
    .A2(_02130_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10176_ (.A1(_02320_),
    .A2(_02322_),
    .B1(_02196_),
    .B2(_02331_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10177_ (.A1(_00575_),
    .A2(_02330_),
    .A3(_02322_),
    .A4(_02320_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _10178_ (.A1(_02332_),
    .A2(_02312_),
    .A3(_02333_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10179_ (.A1(_02334_),
    .A2(_02311_),
    .A3(_02274_),
    .A4(_02202_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10180_ (.A1(_07460_),
    .A2(_02182_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10181_ (.A1(_07460_),
    .A2(_02182_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10182_ (.A1(_00575_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _10183_ (.A1(_02196_),
    .A2(_02336_),
    .B1(_02338_),
    .B2(_02329_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10184_ (.A1(_00575_),
    .A2(_02183_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10185_ (.A1(_02312_),
    .A2(_02340_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10186_ (.A1(_02299_),
    .A2(_02339_),
    .A3(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10187_ (.A1(_02246_),
    .A2(_02260_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10188_ (.A1(_02242_),
    .A2(_02264_),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10189_ (.A1(_02344_),
    .A2(_02309_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10190_ (.A1(_02343_),
    .A2(_02239_),
    .A3(_02345_),
    .B(_02301_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10191_ (.A1(_02171_),
    .A2(_02200_),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10192_ (.A1(_02234_),
    .A2(_02347_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10193_ (.A1(_02342_),
    .A2(_02335_),
    .B(_02346_),
    .C(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10194_ (.A1(_02349_),
    .A2(_02310_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10195_ (.A1(_02201_),
    .A2(_02239_),
    .A3(_02345_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10196_ (.A1(_02145_),
    .A2(_02146_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10197_ (.A1(_02352_),
    .A2(_02235_),
    .B(_02305_),
    .C(_02150_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10198_ (.A1(_02142_),
    .A2(_02353_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10199_ (.A1(_02241_),
    .A2(_02207_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10200_ (.A1(_02142_),
    .A2(_02355_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10201_ (.A1(_02071_),
    .A2(_02354_),
    .A3(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10202_ (.A1(_02136_),
    .A2(_02142_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10203_ (.A1(_02358_),
    .A2(_02242_),
    .B(_02244_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _10204_ (.A1(_02143_),
    .A2(_02355_),
    .B(_02243_),
    .C(_02029_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10205_ (.A1(_02029_),
    .A2(_02359_),
    .B(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10206_ (.A1(_02357_),
    .A2(_02361_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10207_ (.A1(_02029_),
    .A2(_02353_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10208_ (.A1(_02243_),
    .A2(_02029_),
    .B(_02144_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10209_ (.A1(_02363_),
    .A2(_02364_),
    .B(_02358_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10210_ (.A1(_02144_),
    .A2(_02143_),
    .A3(_02242_),
    .A4(_02245_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10211_ (.A1(_02366_),
    .A2(_02260_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10212_ (.A1(_02201_),
    .A2(_02239_),
    .A3(_02345_),
    .A4(_02367_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10213_ (.A1(_02029_),
    .A2(_02359_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10214_ (.A1(_02144_),
    .A2(_02369_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _10215_ (.A1(_02351_),
    .A2(_02362_),
    .A3(_02365_),
    .B1(_02368_),
    .B2(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10216_ (.A1(_02357_),
    .A2(_02361_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10217_ (.A1(_02354_),
    .A2(_02356_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10218_ (.A1(_02071_),
    .A2(_02354_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10219_ (.A1(_02373_),
    .A2(_02374_),
    .A3(_02361_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10220_ (.A1(_02246_),
    .A2(_02260_),
    .B(_02344_),
    .C(_02309_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _10221_ (.A1(_02201_),
    .A2(_02239_),
    .A3(_02376_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10222_ (.I0(_02372_),
    .I1(_02375_),
    .S(_02377_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10223_ (.A1(_02246_),
    .A2(_02260_),
    .A3(_02265_),
    .B(_02309_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10224_ (.A1(_02117_),
    .A2(_02119_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10225_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02380_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10226_ (.A1(_01914_),
    .A2(_02161_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10227_ (.A1(_07436_),
    .A2(_07439_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10228_ (.A1(_02110_),
    .A2(_02221_),
    .A3(_02222_),
    .B(_02383_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10229_ (.A1(_07437_),
    .A2(_07436_),
    .B(_02382_),
    .C(_02384_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10230_ (.A1(_02021_),
    .A2(_02159_),
    .A3(_02306_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10231_ (.A1(_02381_),
    .A2(_02385_),
    .A3(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10232_ (.A1(_02263_),
    .A2(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10233_ (.A1(_02201_),
    .A2(_02239_),
    .A3(_02379_),
    .B(_02388_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10234_ (.A1(_02246_),
    .A2(_02260_),
    .A3(_02265_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _10235_ (.A1(_02213_),
    .A2(_02234_),
    .A3(_02238_),
    .A4(_02309_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _10236_ (.A1(_02201_),
    .A2(_02388_),
    .A3(_02390_),
    .A4(_02391_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10237_ (.A1(_02143_),
    .A2(_02152_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10238_ (.A1(_02393_),
    .A2(_02207_),
    .B(_02254_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10239_ (.A1(_02201_),
    .A2(_02239_),
    .A3(_02345_),
    .A4(_02367_),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10240_ (.A1(net9),
    .A2(_02138_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10241_ (.A1(_02137_),
    .A2(_02396_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10242_ (.A1(_02381_),
    .A2(_02385_),
    .A3(_02263_),
    .A4(_02386_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10243_ (.A1(_02397_),
    .A2(_02398_),
    .B(_02242_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _10244_ (.A1(_02389_),
    .A2(_02392_),
    .B1(_02394_),
    .B2(_02395_),
    .C(_02399_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10245_ (.A1(_02371_),
    .A2(_02378_),
    .A3(_02400_),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _10246_ (.I(_02401_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10247_ (.A1(_02402_),
    .A2(_02350_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10248_ (.I(_02403_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10249_ (.I0(_07470_),
    .I1(_02282_),
    .S(_02404_),
    .Z(_07487_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10250_ (.I(_07494_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10251_ (.A1(_07498_),
    .A2(_07499_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10252_ (.A1(_07497_),
    .A2(_02406_),
    .B(_07495_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10253_ (.A1(_02405_),
    .A2(_02407_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10254_ (.A1(_07492_),
    .A2(_07495_),
    .A3(_07498_),
    .A4(_07500_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10255_ (.A1(_07492_),
    .A2(_02408_),
    .B(_07491_),
    .C(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10256_ (.A1(_07489_),
    .A2(_02410_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10257_ (.A1(_02346_),
    .A2(_02347_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10258_ (.A1(_02202_),
    .A2(_02311_),
    .A3(_02274_),
    .A4(_02334_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10259_ (.A1(_02304_),
    .A2(_02339_),
    .A3(_02341_),
    .B(_02413_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10260_ (.A1(_02412_),
    .A2(_02414_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10261_ (.A1(_07463_),
    .A2(_02328_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _10262_ (.I(_02416_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10263_ (.A1(_01626_),
    .A2(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10264_ (.A1(_02320_),
    .A2(_02322_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10265_ (.I0(_02419_),
    .I1(_02336_),
    .S(_02275_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10266_ (.A1(_02130_),
    .A2(_02329_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10267_ (.A1(_02420_),
    .A2(_02421_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10268_ (.A1(_02415_),
    .A2(_02418_),
    .A3(_02422_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10269_ (.A1(_01666_),
    .A2(_01667_),
    .B(_07342_),
    .ZN(_07361_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10270_ (.A1(_07363_),
    .A2(_07365_),
    .A3(_07364_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10271_ (.A1(_01673_),
    .A2(_02424_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10272_ (.I0(_07361_),
    .I1(_02425_),
    .S(_01879_),
    .Z(_07381_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10273_ (.A1(_07383_),
    .A2(_01751_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10274_ (.I0(_07381_),
    .I1(_02426_),
    .S(_01989_),
    .Z(_07401_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10275_ (.A1(_07403_),
    .A2(_01961_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10276_ (.I0(_07401_),
    .I1(_02427_),
    .S(_02162_),
    .Z(_07421_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10277_ (.A1(_07423_),
    .A2(_02107_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10278_ (.I0(_07421_),
    .I1(_02428_),
    .S(_02121_),
    .Z(_07441_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10279_ (.I(_07441_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10280_ (.A1(_07443_),
    .A2(_02179_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10281_ (.I0(_02429_),
    .I1(_02430_),
    .S(_02275_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10282_ (.I(_02431_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10283_ (.I(_02419_),
    .ZN(_07458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10284_ (.I0(_07458_),
    .I1(_02337_),
    .S(net44),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10285_ (.A1(_01626_),
    .A2(_02432_),
    .B(_02433_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10286_ (.A1(_02350_),
    .A2(_02402_),
    .A3(_02434_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10287_ (.A1(_02332_),
    .A2(_02333_),
    .B(_02312_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10288_ (.A1(_02339_),
    .A2(_02341_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10289_ (.I0(_02436_),
    .I1(_02437_),
    .S(net44),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10290_ (.A1(_02310_),
    .A2(_02349_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10291_ (.I(_02439_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _10292_ (.A1(_02371_),
    .A2(_02378_),
    .A3(_02400_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10293_ (.A1(_02440_),
    .A2(_02441_),
    .B(_02414_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10294_ (.A1(_02423_),
    .A2(_02435_),
    .B(_02438_),
    .C(_02442_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10295_ (.I(_02410_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10296_ (.A1(_02444_),
    .A2(_07489_),
    .B(_07488_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10297_ (.I(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10298_ (.A1(_07486_),
    .A2(_02446_),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10299_ (.A1(_02447_),
    .A2(_07485_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10300_ (.A1(_07483_),
    .A2(_02448_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10301_ (.A1(_02449_),
    .A2(_07482_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10302_ (.A1(_00575_),
    .A2(_02450_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10303_ (.A1(_02416_),
    .A2(_02451_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10304_ (.A1(_02130_),
    .A2(_02450_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10305_ (.A1(_02416_),
    .A2(_02453_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _10306_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02454_),
    .B2(_02452_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10307_ (.A1(_02432_),
    .A2(_02451_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10308_ (.A1(_02432_),
    .A2(_02453_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10309_ (.A1(_02456_),
    .A2(_02457_),
    .B(_02350_),
    .C(_02402_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10310_ (.A1(_02458_),
    .A2(_02455_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10311_ (.A1(_02350_),
    .A2(_02402_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _10312_ (.A1(_02202_),
    .A2(_02311_),
    .A3(_02303_),
    .B1(_02297_),
    .B2(_02213_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10313_ (.A1(_02235_),
    .A2(_02236_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10314_ (.A1(_02021_),
    .A2(_02207_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10315_ (.A1(_02462_),
    .A2(_02463_),
    .B(_02308_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10316_ (.A1(net43),
    .A2(_02311_),
    .A3(_02303_),
    .B(_02464_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10317_ (.A1(net43),
    .A2(_02311_),
    .A3(_02303_),
    .A4(_02464_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10318_ (.A1(_02465_),
    .A2(_02466_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10319_ (.A1(net44),
    .A2(_02299_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10320_ (.A1(_02298_),
    .A2(_02349_),
    .A3(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10321_ (.A1(_02349_),
    .A2(_02468_),
    .B(_02298_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10322_ (.A1(_02461_),
    .A2(_02467_),
    .A3(_02469_),
    .A4(_02470_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10323_ (.A1(_02218_),
    .A2(_02227_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10324_ (.A1(_02219_),
    .A2(_02226_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10325_ (.I(_02473_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _10326_ (.A1(_02472_),
    .A2(_02237_),
    .B1(_02346_),
    .B2(_02474_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10327_ (.A1(_02473_),
    .A2(_02346_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10328_ (.A1(_02468_),
    .A2(_02475_),
    .A3(_02476_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10329_ (.A1(_02460_),
    .A2(_02471_),
    .B(_02477_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10330_ (.A1(_02389_),
    .A2(_02392_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10331_ (.A1(_02310_),
    .A2(_02349_),
    .B(_02479_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10332_ (.A1(_02263_),
    .A2(_02387_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10333_ (.A1(_02298_),
    .A2(_02273_),
    .A3(_02399_),
    .A4(_02481_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10334_ (.A1(_02242_),
    .A2(_02397_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10335_ (.A1(_02263_),
    .A2(_02483_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10336_ (.I(_02397_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10337_ (.A1(_02387_),
    .A2(_02485_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _10338_ (.A1(net43),
    .A2(_02311_),
    .A3(_02379_),
    .B1(_02486_),
    .B2(_02353_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10339_ (.A1(net43),
    .A2(_02311_),
    .A3(_02265_),
    .A4(_02379_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10340_ (.A1(_02484_),
    .A2(_02487_),
    .A3(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10341_ (.A1(_02349_),
    .A2(_02461_),
    .A3(_02482_),
    .B(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _10342_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02480_),
    .B2(_02490_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10343_ (.A1(_02306_),
    .A2(_02463_),
    .B(_02387_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10344_ (.A1(_02301_),
    .A2(_02302_),
    .A3(_02274_),
    .A4(_02464_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10345_ (.A1(_02492_),
    .A2(_02493_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10346_ (.A1(_02346_),
    .A2(_02348_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10347_ (.A1(_02298_),
    .A2(_02461_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10348_ (.A1(_02465_),
    .A2(_02466_),
    .B1(_02389_),
    .B2(_02392_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _10349_ (.A1(_02495_),
    .A2(_02414_),
    .A3(_02496_),
    .A4(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10350_ (.A1(_02373_),
    .A2(_02377_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10351_ (.A1(_02494_),
    .A2(_02498_),
    .B(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10352_ (.A1(_02491_),
    .A2(_02500_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10353_ (.A1(_02459_),
    .A2(_02443_),
    .A3(_02478_),
    .A4(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10354_ (.A1(_07463_),
    .A2(_02328_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10355_ (.A1(_07483_),
    .A2(_07486_),
    .A3(_01392_),
    .A4(_02409_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10356_ (.A1(_07489_),
    .A2(_07177_),
    .A3(_02504_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10357_ (.A1(_02503_),
    .A2(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _10358_ (.I(_02130_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10359_ (.A1(_07489_),
    .A2(_02507_),
    .A3(_02504_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10360_ (.A1(_02417_),
    .A2(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _10361_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02506_),
    .B2(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _10362_ (.I(_02432_),
    .Z(_07461_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10363_ (.A1(_07461_),
    .A2(_02508_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10364_ (.A1(_02431_),
    .A2(_02505_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10365_ (.A1(_02511_),
    .A2(_02512_),
    .B(_02350_),
    .C(_02402_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10366_ (.A1(_02510_),
    .A2(_02513_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10367_ (.I(_02399_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10368_ (.A1(_02371_),
    .A2(_02378_),
    .A3(_02515_),
    .A4(_02479_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10369_ (.A1(_02343_),
    .A2(_02311_),
    .A3(_02345_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10370_ (.A1(_02299_),
    .A2(_02339_),
    .A3(_02341_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10371_ (.A1(_02234_),
    .A2(_02347_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _10372_ (.A1(_02301_),
    .A2(_02517_),
    .B1(_02413_),
    .B2(_02518_),
    .C(_02519_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10373_ (.A1(_02461_),
    .A2(_02482_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10374_ (.A1(_02520_),
    .A2(_02378_),
    .A3(_02521_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _10375_ (.A1(_02440_),
    .A2(_02516_),
    .A3(_02402_),
    .B1(_02522_),
    .B2(_02371_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10376_ (.A1(_02373_),
    .A2(_02377_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10377_ (.A1(_07177_),
    .A2(_02276_),
    .A3(_07458_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10378_ (.A1(_07463_),
    .A2(_07480_),
    .A3(_07466_),
    .A4(_07469_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10379_ (.A1(_07472_),
    .A2(_07475_),
    .A3(_07478_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10380_ (.A1(_01392_),
    .A2(_02374_),
    .A3(_02526_),
    .A4(_02527_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10381_ (.A1(_00575_),
    .A2(_07458_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10382_ (.A1(_02301_),
    .A2(_02302_),
    .A3(_02303_),
    .A4(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10383_ (.A1(net44),
    .A2(_02338_),
    .B(_02528_),
    .C(_02530_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10384_ (.A1(_02524_),
    .A2(_02525_),
    .A3(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10385_ (.A1(_02520_),
    .A2(_02521_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10386_ (.A1(_02071_),
    .A2(_02354_),
    .A3(_02356_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10387_ (.A1(_02402_),
    .A2(_02532_),
    .B(_02533_),
    .C(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10388_ (.A1(_02136_),
    .A2(_02461_),
    .A3(_02356_),
    .A4(_02482_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10389_ (.A1(net43),
    .A2(_02311_),
    .A3(_02376_),
    .B(_02242_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10390_ (.A1(_02071_),
    .A2(_02142_),
    .A3(_02537_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10391_ (.A1(_02142_),
    .A2(_02537_),
    .B(_02071_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10392_ (.A1(_02520_),
    .A2(_02536_),
    .B(_02538_),
    .C(_02539_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10393_ (.A1(_02395_),
    .A2(_02394_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10394_ (.A1(_02202_),
    .A2(_02311_),
    .A3(_02534_),
    .A4(_02376_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10395_ (.A1(_02361_),
    .A2(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10396_ (.A1(_02541_),
    .A2(_02543_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10397_ (.A1(_02540_),
    .A2(_02544_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _10398_ (.A1(_02523_),
    .A2(_02535_),
    .A3(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10399_ (.A1(_02514_),
    .A2(_02546_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10400_ (.A1(_02547_),
    .A2(_02502_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10401_ (.I(_02548_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _10402_ (.I(_02549_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10403_ (.I0(_07487_),
    .I1(_02411_),
    .S(_02550_),
    .Z(_07506_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10404_ (.I(_07519_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10405_ (.A1(_07502_),
    .A2(_07501_),
    .B(_07520_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10406_ (.A1(_02551_),
    .A2(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10407_ (.A1(_07517_),
    .A2(_02553_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10408_ (.A1(_02554_),
    .A2(_07516_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10409_ (.A1(_02555_),
    .A2(_07514_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10410_ (.A1(_02556_),
    .A2(_07513_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10411_ (.A1(_02557_),
    .A2(_07511_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10412_ (.A1(_02558_),
    .A2(_07510_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10413_ (.A1(_07508_),
    .A2(_02559_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _10414_ (.A1(_02443_),
    .A2(_02459_),
    .A3(_02478_),
    .A4(_02501_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10415_ (.A1(_02514_),
    .A2(_02546_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10416_ (.A1(_02443_),
    .A2(_02459_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10417_ (.A1(_02561_),
    .A2(_02562_),
    .B(_02477_),
    .C(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10418_ (.A1(_02130_),
    .A2(_02450_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10419_ (.A1(_02196_),
    .A2(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10420_ (.A1(_02417_),
    .A2(_02566_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _10421_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02452_),
    .B2(_02567_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10422_ (.A1(_07461_),
    .A2(_02566_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10423_ (.A1(_02456_),
    .A2(_02569_),
    .B(net4),
    .C(_02402_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10424_ (.A1(_02568_),
    .A2(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10425_ (.A1(_02438_),
    .A2(_02442_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10426_ (.A1(_02421_),
    .A2(_02415_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10427_ (.A1(net24),
    .A2(_02573_),
    .B(_02433_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10428_ (.A1(_07177_),
    .A2(_02329_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10429_ (.A1(net25),
    .A2(_02433_),
    .A3(_02575_),
    .A4(_02415_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10430_ (.A1(_02574_),
    .A2(_02576_),
    .B(_02476_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10431_ (.A1(_02468_),
    .A2(_02475_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10432_ (.A1(_02473_),
    .A2(_02412_),
    .A3(_02414_),
    .A4(_02403_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10433_ (.A1(_02578_),
    .A2(_02579_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10434_ (.A1(_02571_),
    .A2(_02572_),
    .A3(_02577_),
    .B(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10435_ (.A1(_02418_),
    .A2(_02422_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10436_ (.A1(net25),
    .A2(_02582_),
    .B(_02435_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10437_ (.A1(_02438_),
    .A2(_02442_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10438_ (.A1(_02583_),
    .A2(net15),
    .B(_02584_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10439_ (.A1(_02584_),
    .A2(_02583_),
    .A3(net15),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10440_ (.A1(_02561_),
    .A2(_02562_),
    .B(_02585_),
    .C(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10441_ (.I0(_02414_),
    .I1(_02442_),
    .S(_02412_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10442_ (.A1(_02476_),
    .A2(_02588_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10443_ (.A1(_02564_),
    .A2(_02581_),
    .A3(_02587_),
    .A4(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10444_ (.A1(_01888_),
    .A2(_07365_),
    .ZN(_07384_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10445_ (.A1(_07388_),
    .A2(_07386_),
    .A3(_07387_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10446_ (.A1(_01750_),
    .A2(_02591_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10447_ (.I0(_07384_),
    .I1(_02592_),
    .S(_01989_),
    .Z(_07404_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10448_ (.A1(_07406_),
    .A2(_01959_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10449_ (.I0(_07404_),
    .I1(_02593_),
    .S(_02162_),
    .Z(_07424_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10450_ (.A1(_07426_),
    .A2(_02105_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10451_ (.I0(_07424_),
    .I1(_02594_),
    .S(_02121_),
    .Z(_07444_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10452_ (.A1(_07446_),
    .A2(_02177_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10453_ (.I0(_07444_),
    .I1(_02595_),
    .S(_02276_),
    .Z(_07464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10454_ (.I(_07464_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10455_ (.A1(_07466_),
    .A2(_02326_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _10456_ (.I0(_02596_),
    .I1(_02597_),
    .S(_02403_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10457_ (.A1(_02507_),
    .A2(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10458_ (.A1(_07508_),
    .A2(_02559_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10459_ (.A1(_02600_),
    .A2(_07507_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10460_ (.A1(_02601_),
    .A2(_07505_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10461_ (.A1(_07504_),
    .A2(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _10462_ (.A1(_02196_),
    .A2(_02598_),
    .B1(_02599_),
    .B2(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10463_ (.I(_02452_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10464_ (.A1(_02417_),
    .A2(_02453_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10465_ (.A1(net4),
    .A2(_02402_),
    .B1(_02605_),
    .B2(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10466_ (.A1(_07461_),
    .A2(_02451_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10467_ (.A1(_07461_),
    .A2(_02453_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _10468_ (.A1(_02608_),
    .A2(_02609_),
    .B(_02440_),
    .C(_02441_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10469_ (.A1(_07482_),
    .A2(_02449_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10470_ (.A1(_00758_),
    .A2(_02611_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10471_ (.A1(_02417_),
    .A2(_02612_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _10472_ (.A1(_02607_),
    .A2(_02610_),
    .A3(_02613_),
    .B1(_02421_),
    .B2(_02433_),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10473_ (.A1(_07461_),
    .A2(_02612_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10474_ (.A1(_02460_),
    .A2(_02455_),
    .A3(_02458_),
    .A4(_02615_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10475_ (.A1(net25),
    .A2(_02575_),
    .B(_02420_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10476_ (.A1(net24),
    .A2(_02614_),
    .B(_02616_),
    .C(_02617_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10477_ (.I(_02460_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10478_ (.A1(_02619_),
    .A2(_02431_),
    .A3(_02420_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10479_ (.A1(net24),
    .A2(_02503_),
    .A3(_02422_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10480_ (.A1(_00575_),
    .A2(_02611_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10481_ (.A1(_02565_),
    .A2(_02622_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10482_ (.A1(_07461_),
    .A2(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10483_ (.A1(_02403_),
    .A2(_02420_),
    .A3(_02624_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10484_ (.A1(_02417_),
    .A2(_02623_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10485_ (.A1(_02460_),
    .A2(_02422_),
    .A3(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10486_ (.A1(_02625_),
    .A2(_02627_),
    .B(_02571_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10487_ (.A1(_02618_),
    .A2(_02620_),
    .A3(_02621_),
    .A4(_02628_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10488_ (.A1(_02602_),
    .A2(_07504_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _10489_ (.A1(_07483_),
    .A2(_02448_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10490_ (.A1(_07177_),
    .A2(_02631_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10491_ (.A1(_02196_),
    .A2(_02631_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10492_ (.A1(_02632_),
    .A2(_02630_),
    .B(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _10493_ (.A1(_02561_),
    .A2(_02562_),
    .B1(_02618_),
    .B2(_02628_),
    .C(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10494_ (.A1(_02548_),
    .A2(_02604_),
    .A3(_02629_),
    .B(_02635_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10495_ (.I(_02636_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10496_ (.A1(_02637_),
    .A2(_02590_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10497_ (.A1(_02440_),
    .A2(_02516_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10498_ (.A1(_02541_),
    .A2(_02639_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10499_ (.A1(_02371_),
    .A2(_02522_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10500_ (.A1(_02404_),
    .A2(_02639_),
    .B(_02641_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10501_ (.A1(_02535_),
    .A2(_02540_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10502_ (.A1(_02642_),
    .A2(_02543_),
    .A3(_02643_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10503_ (.A1(_02478_),
    .A2(_02501_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10504_ (.A1(_02563_),
    .A2(_02644_),
    .A3(_02645_),
    .A4(_02562_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10505_ (.A1(_02461_),
    .A2(_02469_),
    .A3(_02470_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10506_ (.A1(_02477_),
    .A2(_02415_),
    .A3(_02418_),
    .A4(_02422_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10507_ (.A1(_02647_),
    .A2(_02648_),
    .B(_02435_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _10508_ (.A1(_02495_),
    .A2(_02414_),
    .A3(_02496_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _10509_ (.A1(net4),
    .A2(_02402_),
    .B(_02650_),
    .C(_02467_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10510_ (.A1(_02650_),
    .A2(_02467_),
    .B(_02651_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10511_ (.A1(_02572_),
    .A2(_02459_),
    .A3(_02649_),
    .B(_02652_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10512_ (.A1(_02572_),
    .A2(_02459_),
    .A3(_02652_),
    .A4(_02649_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10513_ (.A1(_02561_),
    .A2(_02562_),
    .B(_02653_),
    .C(_02654_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10514_ (.A1(_02640_),
    .A2(_02646_),
    .B(_02655_),
    .C(_02642_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10515_ (.A1(_02650_),
    .A2(_02619_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10516_ (.A1(_02473_),
    .A2(_02238_),
    .A3(_02412_),
    .A4(_02414_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10517_ (.I(_02461_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10518_ (.A1(_02578_),
    .A2(_02658_),
    .B(_02659_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10519_ (.A1(_02657_),
    .A2(_02660_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10520_ (.I0(_02582_),
    .I1(_02434_),
    .S(_02460_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10521_ (.A1(_02455_),
    .A2(_02458_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10522_ (.A1(_02304_),
    .A2(_02300_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10523_ (.A1(_02664_),
    .A2(_02477_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10524_ (.A1(_02662_),
    .A2(_02588_),
    .A3(_02663_),
    .A4(_02665_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10525_ (.A1(_02561_),
    .A2(_02562_),
    .B(_02666_),
    .C(_02584_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10526_ (.I(_02477_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10527_ (.A1(_02524_),
    .A2(_02521_),
    .A3(_02525_),
    .A4(_02531_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10528_ (.A1(_02310_),
    .A2(_02441_),
    .A3(_02669_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10529_ (.A1(_02238_),
    .A2(_02520_),
    .A3(_02670_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10530_ (.A1(_02664_),
    .A2(_02520_),
    .B(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10531_ (.A1(_02668_),
    .A2(_02443_),
    .A3(net15),
    .B(_02672_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _10532_ (.A1(_02661_),
    .A2(_02667_),
    .A3(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10533_ (.A1(_02441_),
    .A2(_02669_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10534_ (.A1(_02520_),
    .A2(_02675_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10535_ (.A1(_02650_),
    .A2(_02467_),
    .B(_02494_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10536_ (.A1(_02310_),
    .A2(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10537_ (.A1(_02494_),
    .A2(_02676_),
    .B(_02678_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10538_ (.A1(net44),
    .A2(_02340_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10539_ (.A1(_02312_),
    .A2(_02680_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10540_ (.A1(_02495_),
    .A2(_02669_),
    .A3(_02681_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10541_ (.A1(_02441_),
    .A2(_02682_),
    .B(net4),
    .C(_02388_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10542_ (.A1(net4),
    .A2(_02479_),
    .B(_02683_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10543_ (.A1(_02484_),
    .A2(_02487_),
    .A3(_02488_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10544_ (.A1(_02440_),
    .A2(_02481_),
    .B(_02685_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10545_ (.A1(_02533_),
    .A2(_02686_),
    .B(_02619_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10546_ (.A1(_02499_),
    .A2(_02679_),
    .A3(_02684_),
    .A4(_02687_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10547_ (.A1(_02491_),
    .A2(_02500_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10548_ (.A1(_02443_),
    .A2(_02459_),
    .A3(_02478_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10549_ (.A1(_02689_),
    .A2(_02546_),
    .B(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _10550_ (.I0(_02501_),
    .I1(_02688_),
    .S(_02691_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10551_ (.A1(_02510_),
    .A2(_02513_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10552_ (.A1(_02523_),
    .A2(_02535_),
    .A3(_02545_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10553_ (.A1(_02693_),
    .A2(_02694_),
    .B(_02643_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _10554_ (.I0(_02643_),
    .I1(_02695_),
    .S(_02502_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10555_ (.A1(_02535_),
    .A2(_02543_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10556_ (.A1(_02696_),
    .A2(_02697_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _10557_ (.A1(_02656_),
    .A2(_02674_),
    .A3(_02692_),
    .A4(_02698_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10558_ (.A1(_02699_),
    .A2(_02638_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10559_ (.I(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10560_ (.I0(_07506_),
    .I1(_02560_),
    .S(_02701_),
    .Z(_07529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10561_ (.I(_07522_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10562_ (.A1(_07525_),
    .A2(_07524_),
    .B(_07523_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10563_ (.A1(_02702_),
    .A2(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10564_ (.A1(_07543_),
    .A2(_02704_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10565_ (.A1(_02705_),
    .A2(_07542_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10566_ (.A1(_02706_),
    .A2(_07540_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10567_ (.A1(_02707_),
    .A2(_07539_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10568_ (.A1(_02708_),
    .A2(_07537_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10569_ (.A1(_02709_),
    .A2(_07536_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10570_ (.A1(_02710_),
    .A2(_07534_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10571_ (.A1(_02711_),
    .A2(_07533_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10572_ (.A1(_07531_),
    .A2(_02712_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10573_ (.A1(_02696_),
    .A2(_02697_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _10574_ (.I(_02584_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10575_ (.A1(_02650_),
    .A2(_02479_),
    .B(_02619_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _10576_ (.A1(_02467_),
    .A2(_02494_),
    .A3(_02660_),
    .A4(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10577_ (.A1(_02666_),
    .A2(_02717_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10578_ (.A1(_02715_),
    .A2(_02549_),
    .A3(_02718_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10579_ (.I(_02684_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10580_ (.A1(_02679_),
    .A2(_02691_),
    .B(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10581_ (.A1(_02719_),
    .A2(_02721_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10582_ (.A1(_02679_),
    .A2(_02691_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _10583_ (.I(_02723_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10584_ (.A1(_02652_),
    .A2(_02661_),
    .A3(_02667_),
    .A4(_02673_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10585_ (.A1(_02590_),
    .A2(_02636_),
    .A3(_02725_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10586_ (.A1(_02724_),
    .A2(_02726_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10587_ (.A1(_02687_),
    .A2(_02722_),
    .A3(_02727_),
    .B(net29),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10588_ (.A1(_02656_),
    .A2(_02674_),
    .A3(_02692_),
    .A4(_02698_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10589_ (.A1(_02590_),
    .A2(_02729_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _10590_ (.A1(_02590_),
    .A2(_02637_),
    .A3(_02725_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10591_ (.A1(_02723_),
    .A2(_02722_),
    .A3(_02731_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10592_ (.A1(_02520_),
    .A2(_02521_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10593_ (.A1(net24),
    .A2(_02733_),
    .B1(_02686_),
    .B2(_02719_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10594_ (.A1(_02499_),
    .A2(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10595_ (.A1(_02687_),
    .A2(_02730_),
    .A3(_02732_),
    .B(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10596_ (.I(_02655_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10597_ (.A1(_02523_),
    .A2(_02737_),
    .A3(_02692_),
    .A4(_02698_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10598_ (.A1(_02640_),
    .A2(_02646_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10599_ (.I(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10600_ (.A1(_02638_),
    .A2(_02674_),
    .A3(_02738_),
    .B(_02740_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10601_ (.A1(_02692_),
    .A2(_02698_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10602_ (.I(_02687_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10603_ (.A1(_02524_),
    .A2(_02743_),
    .A3(_02543_),
    .A4(_02643_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10604_ (.A1(_02715_),
    .A2(_02549_),
    .A3(_02744_),
    .A4(_02718_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10605_ (.A1(_02642_),
    .A2(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10606_ (.A1(_02742_),
    .A2(_02731_),
    .B(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10607_ (.A1(_02657_),
    .A2(_02660_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10608_ (.A1(_02656_),
    .A2(_02748_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10609_ (.A1(_02742_),
    .A2(_02746_),
    .A3(_02731_),
    .A4(_02749_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10610_ (.A1(_02741_),
    .A2(_02747_),
    .A3(_02750_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10611_ (.A1(_02714_),
    .A2(_02728_),
    .A3(_02736_),
    .A4(_02751_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10612_ (.A1(_02588_),
    .A2(_02587_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10613_ (.A1(_02753_),
    .A2(_02637_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10614_ (.A1(_02715_),
    .A2(net14),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10615_ (.A1(_02563_),
    .A2(net14),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10616_ (.A1(_02412_),
    .A2(_02414_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10617_ (.A1(_02619_),
    .A2(_02757_),
    .B(_02346_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10618_ (.A1(_02474_),
    .A2(_02758_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _10619_ (.A1(_02571_),
    .A2(_02577_),
    .A3(_02755_),
    .B1(_02756_),
    .B2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10620_ (.A1(_02564_),
    .A2(_02581_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10621_ (.A1(_02754_),
    .A2(_02760_),
    .B(_02761_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10622_ (.A1(_02662_),
    .A2(_02663_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10623_ (.A1(net45),
    .A2(_02763_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10624_ (.A1(_02568_),
    .A2(_02570_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10625_ (.A1(_02420_),
    .A2(_02575_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10626_ (.A1(net24),
    .A2(_02766_),
    .B(_02617_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10627_ (.A1(_02765_),
    .A2(net45),
    .B(_02767_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10628_ (.A1(_02764_),
    .A2(_02768_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10629_ (.A1(_02502_),
    .A2(_02547_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _10630_ (.I0(_07461_),
    .I1(_02417_),
    .S(net25),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10631_ (.A1(_07177_),
    .A2(_02771_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10632_ (.A1(_02440_),
    .A2(_02441_),
    .A3(_07461_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10633_ (.A1(_02619_),
    .A2(_02417_),
    .B(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10634_ (.A1(_02774_),
    .A2(_02453_),
    .A3(_02630_),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10635_ (.A1(_02774_),
    .A2(_02450_),
    .A3(_02603_),
    .B(_02622_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10636_ (.A1(_02620_),
    .A2(_02621_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10637_ (.A1(_02772_),
    .A2(_02775_),
    .A3(_02776_),
    .B(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10638_ (.A1(_02770_),
    .A2(_02598_),
    .A3(_02778_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10639_ (.I(_02598_),
    .ZN(_07481_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10640_ (.A1(_00977_),
    .A2(_02771_),
    .A3(_02603_),
    .A4(_07481_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10641_ (.A1(_02507_),
    .A2(_02630_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10642_ (.A1(_02611_),
    .A2(_02781_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10643_ (.I0(_02622_),
    .I1(_02782_),
    .S(_02417_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10644_ (.I0(_02622_),
    .I1(_02782_),
    .S(_07461_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10645_ (.I0(_02783_),
    .I1(_02784_),
    .S(_02619_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10646_ (.A1(_02774_),
    .A2(_02451_),
    .B(_02631_),
    .C(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10647_ (.A1(_01626_),
    .A2(_02507_),
    .A3(_02630_),
    .A4(_02631_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10648_ (.A1(_02619_),
    .A2(_02417_),
    .B(_02773_),
    .C(_02623_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10649_ (.A1(_02771_),
    .A2(_02450_),
    .A3(_02787_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _10650_ (.A1(_02775_),
    .A2(_02786_),
    .B1(_02787_),
    .B2(_02788_),
    .C(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10651_ (.I0(_02780_),
    .I1(_02790_),
    .S(_02549_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10652_ (.A1(_02565_),
    .A2(_02622_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10653_ (.A1(_02771_),
    .A2(_02792_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10654_ (.A1(_02561_),
    .A2(_02562_),
    .B(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10655_ (.A1(_02774_),
    .A2(_02514_),
    .A3(_02546_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10656_ (.A1(_02774_),
    .A2(_02623_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10657_ (.A1(_02502_),
    .A2(_02795_),
    .B(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10658_ (.A1(_00758_),
    .A2(_02603_),
    .B(_02781_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10659_ (.A1(_02794_),
    .A2(_02797_),
    .B(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10660_ (.A1(_07531_),
    .A2(_02712_),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10661_ (.A1(_02800_),
    .A2(_07530_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10662_ (.A1(_02801_),
    .A2(_07528_),
    .B(_07527_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _10663_ (.A1(_02779_),
    .A2(_02791_),
    .A3(_02799_),
    .B(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10664_ (.A1(_02792_),
    .A2(_02634_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10665_ (.I0(_02604_),
    .I1(_02804_),
    .S(_02548_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10666_ (.A1(_02771_),
    .A2(_02805_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10667_ (.A1(_07177_),
    .A2(_02603_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10668_ (.A1(_02802_),
    .A2(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10669_ (.A1(_02631_),
    .A2(_02808_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10670_ (.A1(_02507_),
    .A2(_02603_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10671_ (.A1(_02810_),
    .A2(_02802_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10672_ (.A1(_02631_),
    .A2(_02811_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _10673_ (.A1(net3),
    .A2(_02547_),
    .B(_02809_),
    .C(_02812_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10674_ (.I(_02811_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10675_ (.I0(_02808_),
    .I1(_02814_),
    .S(_02598_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _10676_ (.A1(_02502_),
    .A2(_02547_),
    .A3(_02815_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10677_ (.A1(_02813_),
    .A2(_02816_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _10678_ (.A1(_02638_),
    .A2(_02699_),
    .A3(_02803_),
    .B1(_02817_),
    .B2(_02806_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10679_ (.A1(_02564_),
    .A2(_02581_),
    .A3(_02587_),
    .A4(_02589_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10680_ (.A1(_02715_),
    .A2(_02634_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10681_ (.A1(_02715_),
    .A2(_02763_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10682_ (.A1(_02618_),
    .A2(_02628_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10683_ (.I0(_02820_),
    .I1(_02821_),
    .S(_02822_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10684_ (.A1(_02715_),
    .A2(_02763_),
    .A3(_02634_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10685_ (.A1(_02715_),
    .A2(_02549_),
    .A3(_02763_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10686_ (.A1(net14),
    .A2(_02604_),
    .A3(_02629_),
    .B(_02588_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10687_ (.A1(_02823_),
    .A2(_02824_),
    .A3(_02825_),
    .A4(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10688_ (.A1(_02819_),
    .A2(_02699_),
    .B(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10689_ (.A1(_02762_),
    .A2(_02769_),
    .A3(_02828_),
    .A4(_02818_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10690_ (.A1(_02667_),
    .A2(_02673_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10691_ (.A1(_02590_),
    .A2(_02637_),
    .A3(_02830_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10692_ (.A1(_02656_),
    .A2(_02748_),
    .A3(_02692_),
    .A4(_02698_),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10693_ (.A1(_02590_),
    .A2(_02637_),
    .A3(_02661_),
    .A4(_02830_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10694_ (.A1(_02656_),
    .A2(_02692_),
    .A3(_02698_),
    .B(_02725_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10695_ (.A1(_02572_),
    .A2(net15),
    .A3(_02649_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _10696_ (.A1(net14),
    .A2(_02835_),
    .B1(_02748_),
    .B2(_02667_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10697_ (.A1(_02655_),
    .A2(_02836_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _10698_ (.A1(_02833_),
    .A2(_02834_),
    .B1(_02837_),
    .B2(_02731_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10699_ (.A1(_02590_),
    .A2(net11),
    .B(_02830_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10700_ (.A1(_02831_),
    .A2(_02832_),
    .B(_02838_),
    .C(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10701_ (.A1(_02829_),
    .A2(_02840_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10702_ (.I(_02841_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10703_ (.A1(_02842_),
    .A2(_02752_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10704_ (.I(_02843_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10705_ (.I0(_07529_),
    .I1(_02713_),
    .S(_02844_),
    .Z(_07552_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10706_ (.A1(_07457_),
    .A2(_02304_),
    .ZN(_07476_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10707_ (.A1(_07480_),
    .A2(_07478_),
    .A3(_07479_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10708_ (.A1(_02278_),
    .A2(_02845_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10709_ (.I0(_07476_),
    .I1(_02846_),
    .S(_02404_),
    .Z(_07493_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10710_ (.I(_07497_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10711_ (.A1(_07500_),
    .A2(_07499_),
    .B(_07498_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10712_ (.A1(_02847_),
    .A2(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10713_ (.A1(_07495_),
    .A2(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10714_ (.I0(_07493_),
    .I1(_02850_),
    .S(_02550_),
    .Z(_07512_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10715_ (.A1(_07514_),
    .A2(_02555_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10716_ (.I0(_07512_),
    .I1(_02851_),
    .S(_02701_),
    .Z(_07535_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10717_ (.A1(_07537_),
    .A2(_02708_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10718_ (.I0(_07535_),
    .I1(_02852_),
    .S(_02844_),
    .Z(_07558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10719_ (.I(_07550_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10720_ (.A1(_07545_),
    .A2(_07544_),
    .B(_07551_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10721_ (.A1(_02853_),
    .A2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10722_ (.A1(_07548_),
    .A2(_02855_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10723_ (.A1(_07547_),
    .A2(_02856_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10724_ (.A1(_07566_),
    .A2(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10725_ (.A1(_02858_),
    .A2(_07565_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10726_ (.A1(_07563_),
    .A2(_02859_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10727_ (.A1(_02860_),
    .A2(_07562_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10728_ (.A1(_07560_),
    .A2(_02861_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10729_ (.A1(_02829_),
    .A2(_02840_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10730_ (.A1(_02561_),
    .A2(_02695_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10731_ (.A1(_02864_),
    .A2(_02697_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10732_ (.I(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10733_ (.A1(_02866_),
    .A2(_02741_),
    .A3(_02747_),
    .A4(_02750_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _10734_ (.A1(_02696_),
    .A2(_02728_),
    .A3(_02736_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10735_ (.A1(_02692_),
    .A2(_02731_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10736_ (.A1(_02656_),
    .A2(_02742_),
    .B(_02869_),
    .C(_02696_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10737_ (.A1(_02742_),
    .A2(_02731_),
    .A3(_02749_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10738_ (.A1(_02865_),
    .A2(_02870_),
    .B(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10739_ (.A1(_02863_),
    .A2(_02867_),
    .A3(_02868_),
    .B(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10740_ (.A1(_02863_),
    .A2(_02872_),
    .A3(_02867_),
    .A4(_02868_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10741_ (.A1(_02698_),
    .A2(_02746_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10742_ (.A1(_02875_),
    .A2(_02728_),
    .A3(_02736_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10743_ (.A1(net41),
    .A2(_02876_),
    .B(_02741_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10744_ (.A1(_02873_),
    .A2(_02874_),
    .B(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10745_ (.A1(_02714_),
    .A2(_02728_),
    .A3(_02736_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10746_ (.A1(_02842_),
    .A2(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10747_ (.A1(_02747_),
    .A2(_02750_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10748_ (.A1(_02741_),
    .A2(_02881_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10749_ (.A1(_02714_),
    .A2(_02728_),
    .A3(_02736_),
    .A4(_02751_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10750_ (.A1(_07505_),
    .A2(_02601_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10751_ (.I0(_02598_),
    .I1(_02631_),
    .S(net14),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10752_ (.A1(_02810_),
    .A2(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10753_ (.A1(_02884_),
    .A2(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10754_ (.A1(_07388_),
    .A2(_01882_),
    .ZN(_07407_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10755_ (.A1(_07411_),
    .A2(_07409_),
    .A3(_07410_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10756_ (.A1(_01958_),
    .A2(_02888_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10757_ (.I0(_07407_),
    .I1(_02889_),
    .S(_02162_),
    .Z(_07427_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10758_ (.A1(_07429_),
    .A2(_02103_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10759_ (.I0(_07427_),
    .I1(_02890_),
    .S(_02121_),
    .Z(_07447_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10760_ (.A1(_07452_),
    .A2(_02125_),
    .B(_07451_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10761_ (.A1(_07449_),
    .A2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10762_ (.I0(_07447_),
    .I1(_02892_),
    .S(_02276_),
    .Z(_07467_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10763_ (.A1(_07469_),
    .A2(_02324_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10764_ (.I0(_07467_),
    .I1(_02893_),
    .S(_02404_),
    .Z(_07484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10765_ (.I(_07484_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10766_ (.A1(_07486_),
    .A2(_02445_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10767_ (.I0(_02894_),
    .I1(_02895_),
    .S(_02550_),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10768_ (.A1(_02885_),
    .A2(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10769_ (.I(_02699_),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10770_ (.A1(_02638_),
    .A2(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10771_ (.I0(_02887_),
    .I1(_02897_),
    .S(_02899_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10772_ (.A1(_07528_),
    .A2(_02801_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10773_ (.A1(_02638_),
    .A2(_02898_),
    .B(_02807_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _10774_ (.A1(_02802_),
    .A2(_02885_),
    .A3(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10775_ (.A1(_02901_),
    .A2(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10776_ (.A1(_02590_),
    .A2(_02729_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10777_ (.A1(_02572_),
    .A2(_02763_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10778_ (.A1(_02572_),
    .A2(_02763_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _10779_ (.A1(_02770_),
    .A2(_02906_),
    .A3(_02907_),
    .A4(_02635_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10780_ (.A1(_02656_),
    .A2(_02692_),
    .A3(_02698_),
    .B(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10781_ (.A1(_02587_),
    .A2(net11),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10782_ (.A1(_02905_),
    .A2(_02909_),
    .A3(_02910_),
    .Z(_02911_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _10783_ (.A1(_02883_),
    .A2(_02863_),
    .A3(_02900_),
    .B1(_02904_),
    .B2(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10784_ (.A1(_02476_),
    .A2(_02753_),
    .A3(net11),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10785_ (.A1(_02819_),
    .A2(_02898_),
    .B(_02913_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10786_ (.A1(_02831_),
    .A2(_02832_),
    .B(_02839_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10787_ (.A1(_02914_),
    .A2(_02762_),
    .A3(_02915_),
    .Z(_02916_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _10788_ (.A1(_02769_),
    .A2(_02818_),
    .A3(_02828_),
    .Z(_02917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10789_ (.A1(_02916_),
    .A2(_02917_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10790_ (.A1(_07545_),
    .A2(_07554_),
    .A3(_07557_),
    .A4(_07563_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10791_ (.A1(_07548_),
    .A2(_07551_),
    .A3(_07560_),
    .A4(_07566_),
    .Z(_02920_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10792_ (.A1(_01392_),
    .A2(_02919_),
    .A3(_02920_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10793_ (.A1(_02794_),
    .A2(_02797_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10794_ (.A1(net45),
    .A2(_02604_),
    .Z(_02923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10795_ (.A1(net45),
    .A2(net7),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10796_ (.A1(_02923_),
    .A2(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10797_ (.A1(net23),
    .A2(_02898_),
    .B(_02922_),
    .C(_02925_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10798_ (.A1(_02922_),
    .A2(_02925_),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10799_ (.A1(_02921_),
    .A2(_02926_),
    .A3(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10800_ (.A1(_02838_),
    .A2(_02928_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10801_ (.A1(_02813_),
    .A2(_02816_),
    .B(_02771_),
    .C(_02623_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10802_ (.A1(_02770_),
    .A2(_02604_),
    .A3(_02815_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10803_ (.A1(_02604_),
    .A2(_02815_),
    .B(_02771_),
    .C(_02770_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10804_ (.A1(_02930_),
    .A2(_02931_),
    .A3(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10805_ (.A1(net7),
    .A2(_02812_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _10806_ (.A1(net7),
    .A2(_02809_),
    .B(_02771_),
    .C(_02623_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10807_ (.A1(_02598_),
    .A2(_02811_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _10808_ (.A1(net3),
    .A2(_02547_),
    .A3(_02634_),
    .A4(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10809_ (.A1(_02770_),
    .A2(_02934_),
    .B(_02935_),
    .C(_02937_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10810_ (.A1(_02809_),
    .A2(_02788_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10811_ (.A1(net3),
    .A2(_02547_),
    .A3(_02936_),
    .A4(_02788_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10812_ (.A1(_02812_),
    .A2(_02788_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10813_ (.A1(net3),
    .A2(_02547_),
    .B(_02941_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10814_ (.A1(net7),
    .A2(_02939_),
    .A3(_02940_),
    .A4(_02942_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10815_ (.A1(_02938_),
    .A2(_02943_),
    .B(_02770_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10816_ (.A1(_02933_),
    .A2(_02944_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10817_ (.A1(net23),
    .A2(_02898_),
    .B(_02769_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _10818_ (.A1(_02764_),
    .A2(_02768_),
    .B1(_02933_),
    .B2(_02944_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _10819_ (.A1(net29),
    .A2(_02803_),
    .B1(_02945_),
    .B2(_02946_),
    .C(_02947_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _10820_ (.A1(_02883_),
    .A2(_02918_),
    .A3(_02929_),
    .B1(_02928_),
    .B2(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10821_ (.A1(_02747_),
    .A2(_02750_),
    .B1(_02842_),
    .B2(_02879_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _10822_ (.A1(_02880_),
    .A2(_02882_),
    .B1(_02912_),
    .B2(_02949_),
    .C(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10823_ (.A1(_02878_),
    .A2(_02951_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10824_ (.A1(_02696_),
    .A2(_02728_),
    .A3(_02867_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10825_ (.A1(_02842_),
    .A2(_02953_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10826_ (.A1(_02836_),
    .A2(_02914_),
    .A3(_02762_),
    .A4(_02915_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10827_ (.A1(_02833_),
    .A2(_02834_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10828_ (.A1(_02737_),
    .A2(_02726_),
    .B(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10829_ (.A1(_02917_),
    .A2(_02955_),
    .B(_02957_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _10830_ (.A1(_02868_),
    .A2(_02954_),
    .A3(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10831_ (.A1(_02883_),
    .A2(_02863_),
    .A3(_02900_),
    .B(_02904_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10832_ (.A1(_07560_),
    .A2(_02861_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10833_ (.A1(_07559_),
    .A2(_02961_),
    .Z(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10834_ (.A1(_07557_),
    .A2(_02962_),
    .Z(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10835_ (.A1(_02963_),
    .A2(_07556_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10836_ (.A1(_07554_),
    .A2(_02964_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10837_ (.A1(_02965_),
    .A2(_07553_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10838_ (.A1(_02960_),
    .A2(_02966_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10839_ (.A1(_02769_),
    .A2(_02818_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10840_ (.I(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10841_ (.A1(_02819_),
    .A2(_02898_),
    .B(_02909_),
    .C(_02910_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10842_ (.I(_02885_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10843_ (.A1(_02802_),
    .A2(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10844_ (.A1(_02802_),
    .A2(_02885_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10845_ (.I0(_02972_),
    .I1(_02973_),
    .S(_02902_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10846_ (.A1(_02819_),
    .A2(_02898_),
    .B(_02925_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10847_ (.A1(net45),
    .A2(_02777_),
    .B(_02822_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _10848_ (.A1(_02924_),
    .A2(_02793_),
    .A3(_02796_),
    .B1(_02923_),
    .B2(_02774_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10849_ (.A1(_02975_),
    .A2(_02976_),
    .B1(_02977_),
    .B2(_02769_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10850_ (.A1(_02974_),
    .A2(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10851_ (.A1(_02926_),
    .A2(_02927_),
    .Z(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10852_ (.A1(_02885_),
    .A2(_02902_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10853_ (.A1(_02948_),
    .A2(_02980_),
    .B(_02802_),
    .C(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10854_ (.A1(_02969_),
    .A2(_02970_),
    .A3(_02979_),
    .A4(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10855_ (.A1(_02412_),
    .A2(_02414_),
    .Z(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10856_ (.A1(_02619_),
    .A2(_02757_),
    .B(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10857_ (.A1(_02985_),
    .A2(_02764_),
    .A3(_02819_),
    .A4(_02699_),
    .Z(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10858_ (.A1(_02715_),
    .A2(_02985_),
    .A3(net11),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10859_ (.A1(_02764_),
    .A2(net11),
    .B(_02715_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10860_ (.A1(_02715_),
    .A2(_02985_),
    .A3(_02764_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10861_ (.A1(_02588_),
    .A2(_02988_),
    .B(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10862_ (.A1(_02986_),
    .A2(_02987_),
    .A3(_02990_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10863_ (.A1(_02769_),
    .A2(_02818_),
    .A3(_02970_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10864_ (.A1(_02991_),
    .A2(_02992_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _10865_ (.A1(_02752_),
    .A2(net41),
    .B1(_02993_),
    .B2(_02916_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10866_ (.A1(_02667_),
    .A2(_02673_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10867_ (.A1(_02995_),
    .A2(_02836_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10868_ (.A1(_02995_),
    .A2(_02836_),
    .Z(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10869_ (.A1(net23),
    .A2(_02997_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10870_ (.A1(net23),
    .A2(_02729_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10871_ (.A1(_02836_),
    .A2(_02999_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10872_ (.I0(_03000_),
    .I1(_02997_),
    .S(_02829_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10873_ (.A1(_02898_),
    .A2(_02996_),
    .A3(_02998_),
    .A4(_03001_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10874_ (.A1(_02843_),
    .A2(_02983_),
    .B(_02994_),
    .C(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _10875_ (.A1(_02959_),
    .A2(_02967_),
    .A3(_03003_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10876_ (.A1(_03004_),
    .A2(_02952_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _10877_ (.I(_03005_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10878_ (.I0(_07558_),
    .I1(_02862_),
    .S(_03006_),
    .Z(_07581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10879_ (.I(_07574_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10880_ (.A1(_07577_),
    .A2(_07576_),
    .B(_07575_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10881_ (.A1(_03007_),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10882_ (.A1(_03009_),
    .A2(_07572_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10883_ (.A1(_03010_),
    .A2(_07571_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10884_ (.A1(_07569_),
    .A2(_03011_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10885_ (.A1(_03012_),
    .A2(_07568_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10886_ (.A1(_07589_),
    .A2(_03013_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10887_ (.A1(_07588_),
    .A2(_03014_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10888_ (.A1(_07586_),
    .A2(_03015_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10889_ (.A1(_03016_),
    .A2(_07585_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10890_ (.A1(_07583_),
    .A2(_03017_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10891_ (.A1(_02959_),
    .A2(_02967_),
    .A3(_03003_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10892_ (.A1(_02728_),
    .A2(_02736_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10893_ (.A1(_02883_),
    .A2(net41),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10894_ (.A1(_03020_),
    .A2(_03021_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10895_ (.A1(_02696_),
    .A2(_02869_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10896_ (.A1(_02870_),
    .A2(_03023_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10897_ (.A1(_03022_),
    .A2(_03024_),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _10898_ (.A1(net41),
    .A2(_02953_),
    .B(_02958_),
    .C(_03020_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10899_ (.A1(_03026_),
    .A2(_02967_),
    .A3(_03003_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10900_ (.I0(_02881_),
    .I1(_02882_),
    .S(_02880_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10901_ (.A1(_03025_),
    .A2(_03027_),
    .B(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _10902_ (.A1(_02951_),
    .A2(_03019_),
    .B(_03029_),
    .C(_02878_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10903_ (.A1(_02878_),
    .A2(_02951_),
    .A3(_02959_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10904_ (.A1(_03002_),
    .A2(_02994_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10905_ (.A1(_02752_),
    .A2(_02842_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10906_ (.A1(_07528_),
    .A2(_02801_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10907_ (.A1(net29),
    .A2(_02884_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10908_ (.A1(_02899_),
    .A2(_02896_),
    .B(_03035_),
    .ZN(_07526_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _10909_ (.A1(_07529_),
    .A2(_02883_),
    .A3(_02863_),
    .A4(_07526_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10910_ (.A1(net384),
    .A2(_02713_),
    .A3(_03034_),
    .B(_03036_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10911_ (.A1(net23),
    .A2(_02898_),
    .A3(_02897_),
    .Z(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10912_ (.A1(_02899_),
    .A2(_02887_),
    .B(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _10913_ (.A1(_07553_),
    .A2(_02838_),
    .A3(_02965_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10914_ (.A1(_02916_),
    .A2(_02917_),
    .A3(_03039_),
    .A4(_03040_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10915_ (.A1(_02901_),
    .A2(_02903_),
    .A3(_02966_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10916_ (.A1(_02752_),
    .A2(_03041_),
    .B(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10917_ (.A1(_02843_),
    .A2(_02983_),
    .B(_03043_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10918_ (.A1(_03032_),
    .A2(_03037_),
    .A3(_03044_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10919_ (.A1(_07554_),
    .A2(_02964_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10920_ (.I(_03046_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10921_ (.I0(_03034_),
    .I1(_07526_),
    .S(_03033_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10922_ (.A1(_02966_),
    .A2(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _10923_ (.A1(_03031_),
    .A2(_03045_),
    .B1(_03047_),
    .B2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _10924_ (.A1(_02878_),
    .A2(_02951_),
    .A3(_02959_),
    .A4(_03003_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10925_ (.A1(_02968_),
    .A2(_02970_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10926_ (.A1(_07553_),
    .A2(_02904_),
    .A3(_02965_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10927_ (.A1(_02730_),
    .A2(_02754_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _10928_ (.A1(_02760_),
    .A2(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10929_ (.A1(_02991_),
    .A2(_03055_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10930_ (.A1(_03052_),
    .A2(_03053_),
    .B(_03056_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10931_ (.I(_02991_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10932_ (.A1(_03058_),
    .A2(_03052_),
    .A3(_03043_),
    .A4(_03055_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10933_ (.A1(_02843_),
    .A2(_02983_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10934_ (.A1(_03057_),
    .A2(_03059_),
    .B(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10935_ (.A1(net384),
    .A2(_03043_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10936_ (.A1(_03051_),
    .A2(_03061_),
    .A3(_03062_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10937_ (.A1(_07569_),
    .A2(_07577_),
    .A3(_07586_),
    .A4(_07589_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10938_ (.A1(_07580_),
    .A2(_07572_),
    .A3(_07575_),
    .A4(_07583_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10939_ (.A1(_01392_),
    .A2(_03064_),
    .A3(_03065_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _10940_ (.A1(_02878_),
    .A2(_02951_),
    .A3(_02959_),
    .A4(_03003_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10941_ (.A1(_02901_),
    .A2(_02966_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10942_ (.A1(_03033_),
    .A2(_02903_),
    .A3(_03068_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _10943_ (.A1(_03043_),
    .A2(_03067_),
    .B(_03069_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _10944_ (.A1(_03050_),
    .A2(_03063_),
    .A3(_03066_),
    .A4(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10945_ (.I(_02915_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10946_ (.A1(_02883_),
    .A2(_03072_),
    .A3(_02838_),
    .B(_02829_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10947_ (.A1(_02917_),
    .A2(_02843_),
    .A3(_03055_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10948_ (.I(_02761_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10949_ (.A1(_03075_),
    .A2(_02913_),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10950_ (.A1(_02999_),
    .A2(_03076_),
    .Z(_03077_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _10951_ (.A1(_03074_),
    .A2(_03077_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10952_ (.A1(_03073_),
    .A2(_03078_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10953_ (.A1(_02979_),
    .A2(_02982_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10954_ (.I(_07553_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10955_ (.A1(_03033_),
    .A2(_03080_),
    .B(_02912_),
    .C(_03081_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _10956_ (.A1(_02993_),
    .A2(_03055_),
    .B(net384),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10957_ (.A1(_02960_),
    .A2(_02980_),
    .A3(_02965_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10958_ (.A1(_03082_),
    .A2(_03083_),
    .A3(_03084_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10959_ (.A1(_02952_),
    .A2(_03004_),
    .B(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10960_ (.A1(_03079_),
    .A2(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10961_ (.A1(_03032_),
    .A2(_03044_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _10962_ (.A1(_07554_),
    .A2(_07557_),
    .A3(_02961_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10963_ (.A1(_07557_),
    .A2(_07559_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10964_ (.A1(_07556_),
    .A2(_03090_),
    .B(_07554_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10965_ (.A1(_03034_),
    .A2(_03089_),
    .B(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10966_ (.A1(_07526_),
    .A2(_03089_),
    .B(_03091_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10967_ (.I0(_03092_),
    .I1(_03093_),
    .S(_03033_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10968_ (.A1(_02994_),
    .A2(_03082_),
    .A3(_03094_),
    .B(_03002_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10969_ (.A1(_07583_),
    .A2(_03017_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10970_ (.A1(_03096_),
    .A2(_07582_),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10971_ (.A1(_07580_),
    .A2(_03097_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10972_ (.A1(_03098_),
    .A2(_07579_),
    .Z(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _10973_ (.I(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10974_ (.A1(_03026_),
    .A2(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10975_ (.A1(_03072_),
    .A2(_02829_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _10976_ (.A1(_02915_),
    .A2(_03073_),
    .B(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10977_ (.A1(_03103_),
    .A2(_03101_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _10978_ (.A1(_03031_),
    .A2(_03088_),
    .B(_03095_),
    .C(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _10979_ (.A1(_03063_),
    .A2(_03050_),
    .A3(_03070_),
    .A4(_03105_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _10980_ (.A1(_03106_),
    .A2(_03071_),
    .A3(_03087_),
    .A4(_03030_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _10981_ (.I(_03107_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10982_ (.I0(_07581_),
    .I1(_03018_),
    .S(_03108_),
    .Z(_07610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10983_ (.I(\butterfly_count[1] ),
    .ZN(_07636_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _10984_ (.I(\butterfly_count[0] ),
    .ZN(_07686_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10985_ (.A1(_07480_),
    .A2(_02619_),
    .ZN(_07496_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10986_ (.A1(_07500_),
    .A2(_07498_),
    .A3(_07499_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10987_ (.A1(_02848_),
    .A2(_03109_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10988_ (.I0(_07496_),
    .I1(_03110_),
    .S(_02550_),
    .Z(_07515_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10989_ (.A1(_07517_),
    .A2(_02553_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10990_ (.I0(_07515_),
    .I1(_03111_),
    .S(_02701_),
    .Z(_07538_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10991_ (.A1(_07540_),
    .A2(_02706_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10992_ (.I0(_07538_),
    .I1(_03112_),
    .S(_02844_),
    .Z(_07561_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10993_ (.A1(_07563_),
    .A2(_02859_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10994_ (.I0(_07561_),
    .I1(_03113_),
    .S(_03006_),
    .Z(_07584_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _10995_ (.A1(_07586_),
    .A2(_03015_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _10996_ (.I(_03108_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10997_ (.I0(_07584_),
    .I1(_03114_),
    .S(_03115_),
    .Z(_07604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10998_ (.I(_07596_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10999_ (.A1(_07591_),
    .A2(_07590_),
    .B(_07597_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11000_ (.A1(_03116_),
    .A2(_03117_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11001_ (.A1(_07594_),
    .A2(_03118_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11002_ (.A1(_03119_),
    .A2(_07593_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11003_ (.A1(_03120_),
    .A2(_07603_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11004_ (.A1(_07602_),
    .A2(_03121_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11005_ (.A1(_03122_),
    .A2(_07600_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11006_ (.A1(_03123_),
    .A2(_07599_),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11007_ (.A1(_03124_),
    .A2(_07609_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11008_ (.A1(_03125_),
    .A2(_07608_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11009_ (.A1(_07606_),
    .A2(net387),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11010_ (.A1(_02873_),
    .A2(_02874_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11011_ (.I(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11012_ (.A1(_03129_),
    .A2(_03004_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11013_ (.A1(_02880_),
    .A2(_02882_),
    .B(_02950_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11014_ (.A1(_02878_),
    .A2(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11015_ (.A1(net35),
    .A2(_02948_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11016_ (.A1(_02970_),
    .A2(_02921_),
    .A3(_02980_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11017_ (.A1(_02960_),
    .A2(_03133_),
    .A3(_03134_),
    .A4(_03032_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11018_ (.A1(_03132_),
    .A2(_03135_),
    .B(_03004_),
    .C(_03129_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11019_ (.I0(_03130_),
    .I1(_03136_),
    .S(_03131_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11020_ (.A1(_03129_),
    .A2(net380),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11021_ (.A1(_02877_),
    .A2(_03028_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11022_ (.A1(_02877_),
    .A2(_03138_),
    .B(_03139_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11023_ (.A1(_03137_),
    .A2(_03140_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11024_ (.I(_02722_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11025_ (.A1(_02724_),
    .A2(_03142_),
    .A3(_02726_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11026_ (.A1(_02905_),
    .A2(_03143_),
    .B(_02719_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11027_ (.A1(_02687_),
    .A2(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _11028_ (.A1(_02878_),
    .A2(_02951_),
    .A3(_02959_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11029_ (.A1(_03032_),
    .A2(_03044_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11030_ (.A1(_02722_),
    .A2(_02726_),
    .B(net29),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11031_ (.A1(_02723_),
    .A2(_03142_),
    .A3(_02726_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11032_ (.A1(_02724_),
    .A2(_03148_),
    .B(_03149_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11033_ (.A1(_02917_),
    .A2(_02955_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11034_ (.A1(_02957_),
    .A2(_03151_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11035_ (.A1(_03021_),
    .A2(_03152_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11036_ (.A1(_03150_),
    .A2(_03153_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11037_ (.A1(_03146_),
    .A2(_03147_),
    .A3(_03154_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11038_ (.A1(_03021_),
    .A2(_03150_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _11039_ (.A1(_03145_),
    .A2(_03155_),
    .A3(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11040_ (.A1(_03021_),
    .A2(_03152_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11041_ (.A1(_02728_),
    .A2(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11042_ (.A1(_02728_),
    .A2(net41),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11043_ (.A1(_02687_),
    .A2(_02735_),
    .A3(_02730_),
    .A4(_02732_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11044_ (.A1(_02736_),
    .A2(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11045_ (.A1(_03088_),
    .A2(_03159_),
    .B(_03160_),
    .C(_03162_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11046_ (.A1(_03026_),
    .A2(_02967_),
    .A3(_03003_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11047_ (.A1(_03132_),
    .A2(_03025_),
    .A3(_03135_),
    .B(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11048_ (.A1(_03022_),
    .A2(_03163_),
    .A3(_03165_),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11049_ (.A1(_02878_),
    .A2(_02951_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11050_ (.A1(_03025_),
    .A2(_03027_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11051_ (.A1(_03167_),
    .A2(net385),
    .B(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11052_ (.A1(_03128_),
    .A2(_03019_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11053_ (.A1(_03170_),
    .A2(_03154_),
    .A3(_03136_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _11054_ (.A1(_03157_),
    .A2(_03166_),
    .A3(_03169_),
    .A4(_03171_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11055_ (.A1(_03146_),
    .A2(_03147_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11056_ (.I(_03103_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11057_ (.A1(_03095_),
    .A2(_03174_),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11058_ (.A1(_03173_),
    .A2(_03175_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11059_ (.A1(_03051_),
    .A2(_03061_),
    .A3(_03062_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11060_ (.A1(_03079_),
    .A2(_03086_),
    .B(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11061_ (.A1(_03050_),
    .A2(_03070_),
    .A3(_03099_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11062_ (.A1(_03176_),
    .A2(_03178_),
    .A3(_03179_),
    .Z(_03180_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11063_ (.A1(_03030_),
    .A2(_03071_),
    .A3(_03106_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11064_ (.A1(_03137_),
    .A2(_03139_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _11065_ (.A1(_03172_),
    .A2(_03180_),
    .A3(_03181_),
    .A4(_03182_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _11066_ (.A1(_02878_),
    .A2(_02951_),
    .A3(_02959_),
    .A4(_03032_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11067_ (.A1(_02914_),
    .A2(_02762_),
    .A3(_02993_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11068_ (.A1(net384),
    .A2(_03185_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11069_ (.A1(_03044_),
    .A2(_03186_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11070_ (.I(_03145_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11071_ (.A1(_02898_),
    .A2(_02726_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11072_ (.I0(_02731_),
    .I1(_03189_),
    .S(_02724_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11073_ (.A1(_03021_),
    .A2(_03190_),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11074_ (.A1(_02724_),
    .A2(_02726_),
    .B(_03142_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11075_ (.A1(_03143_),
    .A2(_03192_),
    .B(net29),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11076_ (.A1(_03188_),
    .A2(_03191_),
    .A3(_03193_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11077_ (.A1(_03184_),
    .A2(_03187_),
    .B(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _11078_ (.A1(_03173_),
    .A2(_03175_),
    .A3(_03158_),
    .A4(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11079_ (.A1(_03178_),
    .A2(_03179_),
    .A3(_03196_),
    .B(_03166_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11080_ (.A1(_03178_),
    .A2(_03166_),
    .A3(_03179_),
    .A4(_03196_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11081_ (.A1(_03087_),
    .A2(net373),
    .B(_03169_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11082_ (.A1(_03087_),
    .A2(net373),
    .A3(_03169_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11083_ (.A1(_03197_),
    .A2(_03198_),
    .B1(_03199_),
    .B2(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _11084_ (.A1(_03106_),
    .A2(_03071_),
    .A3(_03087_),
    .A4(_03030_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11085_ (.A1(_03170_),
    .A2(_03136_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _11086_ (.A1(_03141_),
    .A2(_03183_),
    .B1(_03201_),
    .B2(_03202_),
    .C(_03203_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11087_ (.A1(_02967_),
    .A2(_03051_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11088_ (.A1(_03047_),
    .A2(_03100_),
    .B(_03049_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11089_ (.A1(_03005_),
    .A2(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11090_ (.A1(_03205_),
    .A2(_03069_),
    .A3(_03207_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11091_ (.I0(_07552_),
    .I1(_03046_),
    .S(_03005_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11092_ (.A1(_03099_),
    .A2(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11093_ (.A1(_03126_),
    .A2(_07606_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11094_ (.A1(_03211_),
    .A2(_07605_),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11095_ (.A1(_03212_),
    .A2(_07612_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11096_ (.A1(_03213_),
    .A2(_07611_),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11097_ (.A1(_07580_),
    .A2(_03097_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11098_ (.A1(_03214_),
    .A2(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11099_ (.A1(_03184_),
    .A2(_03187_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11100_ (.A1(_07434_),
    .A2(_02266_),
    .ZN(_07453_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11101_ (.A1(_07457_),
    .A2(_07455_),
    .A3(_07456_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11102_ (.A1(_02124_),
    .A2(_03218_),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11103_ (.I0(_07453_),
    .I1(_03219_),
    .S(_02276_),
    .Z(_07473_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11104_ (.A1(_07475_),
    .A2(_02279_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11105_ (.I0(_07473_),
    .I1(_03220_),
    .S(_02404_),
    .Z(_07490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11106_ (.A1(_07495_),
    .A2(_02849_),
    .B(_07494_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11107_ (.A1(_07492_),
    .A2(_03221_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11108_ (.I0(_07490_),
    .I1(_03222_),
    .S(_02550_),
    .Z(_07509_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11109_ (.A1(_07511_),
    .A2(_02557_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11110_ (.I0(_07509_),
    .I1(_03223_),
    .S(_02701_),
    .Z(_07532_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11111_ (.A1(_07534_),
    .A2(_02710_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11112_ (.I0(_07532_),
    .I1(_03224_),
    .S(_02843_),
    .Z(_07555_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11113_ (.A1(_07552_),
    .A2(_07555_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11114_ (.A1(_07557_),
    .A2(_02962_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11115_ (.A1(_03046_),
    .A2(_03226_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11116_ (.I0(_03225_),
    .I1(_03227_),
    .S(_03005_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11117_ (.A1(_03214_),
    .A2(_03217_),
    .A3(_03228_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _11118_ (.A1(_03210_),
    .A2(_03216_),
    .B1(_03107_),
    .B2(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11119_ (.A1(_03208_),
    .A2(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11120_ (.A1(_03178_),
    .A2(_03179_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11121_ (.A1(_03103_),
    .A2(_03232_),
    .A3(_03181_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11122_ (.A1(_03184_),
    .A2(_03187_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11123_ (.A1(_03103_),
    .A2(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11124_ (.A1(_03174_),
    .A2(_03217_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11125_ (.A1(_03232_),
    .A2(_03235_),
    .B(_03236_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11126_ (.A1(_03233_),
    .A2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11127_ (.A1(_03173_),
    .A2(_03095_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11128_ (.A1(_03050_),
    .A2(_03070_),
    .A3(_03099_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11129_ (.A1(_02926_),
    .A2(_02927_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11130_ (.A1(_02818_),
    .A2(net35),
    .B1(_02974_),
    .B2(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11131_ (.A1(_03205_),
    .A2(_03242_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11132_ (.A1(_03240_),
    .A2(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11133_ (.A1(_03239_),
    .A2(_03244_),
    .B(_03108_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11134_ (.A1(_02967_),
    .A2(_03051_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11135_ (.A1(_02979_),
    .A2(_02982_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11136_ (.A1(net35),
    .A2(_03247_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11137_ (.I(_03242_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11138_ (.I(_03133_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11139_ (.A1(_03246_),
    .A2(_03248_),
    .B1(_03249_),
    .B2(_03250_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _11140_ (.A1(_03133_),
    .A2(_03246_),
    .A3(_03240_),
    .B(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11141_ (.A1(_02952_),
    .A2(_03004_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11142_ (.A1(_02991_),
    .A2(_03052_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11143_ (.A1(_02917_),
    .A2(net35),
    .B(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11144_ (.A1(_02917_),
    .A2(_03055_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _11145_ (.A1(_03044_),
    .A2(_03074_),
    .A3(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11146_ (.A1(_03255_),
    .A2(_03257_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11147_ (.A1(_02969_),
    .A2(_02911_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11148_ (.A1(_03247_),
    .A2(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11149_ (.A1(_03052_),
    .A2(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11150_ (.A1(_03205_),
    .A2(_03259_),
    .B1(_03261_),
    .B2(net35),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11151_ (.A1(_03079_),
    .A2(_03086_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11152_ (.A1(_03253_),
    .A2(_03258_),
    .B(_03262_),
    .C(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11153_ (.A1(_03252_),
    .A2(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11154_ (.A1(_03245_),
    .A2(_03265_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11155_ (.A1(_03238_),
    .A2(_03231_),
    .A3(_03266_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11156_ (.A1(_03180_),
    .A2(_03181_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11157_ (.A1(_03173_),
    .A2(_03158_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11158_ (.A1(_03268_),
    .A2(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11159_ (.I(_03157_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11160_ (.A1(_03146_),
    .A2(_03147_),
    .B(_03158_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11161_ (.A1(_03190_),
    .A2(_03272_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11162_ (.A1(_03176_),
    .A2(_03273_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11163_ (.A1(_03173_),
    .A2(_03175_),
    .A3(_03158_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11164_ (.A1(_03153_),
    .A2(_03191_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11165_ (.A1(_03146_),
    .A2(_03147_),
    .A3(_03158_),
    .A4(_03190_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11166_ (.A1(_03173_),
    .A2(_03191_),
    .B(_03276_),
    .C(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11167_ (.A1(_03178_),
    .A2(_03179_),
    .A3(_03275_),
    .B(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _11168_ (.A1(_03232_),
    .A2(_03181_),
    .A3(_03274_),
    .B(_03279_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11169_ (.I(_03193_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _11170_ (.A1(_03232_),
    .A2(_03181_),
    .A3(_03281_),
    .A4(_03274_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11171_ (.A1(_03178_),
    .A2(_03179_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11172_ (.A1(_02958_),
    .A2(_03031_),
    .A3(_03088_),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11173_ (.A1(_03021_),
    .A2(_03284_),
    .B(_03190_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11174_ (.A1(_03193_),
    .A2(_03285_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11175_ (.A1(_03021_),
    .A2(_03284_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11176_ (.A1(_03287_),
    .A2(_03190_),
    .B1(_03273_),
    .B2(_03176_),
    .C(_03281_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11177_ (.A1(_03193_),
    .A2(_03285_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11178_ (.A1(_03283_),
    .A2(_03286_),
    .B(_03288_),
    .C(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11179_ (.A1(_03271_),
    .A2(_03280_),
    .A3(_03282_),
    .A4(_03290_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11180_ (.A1(_03270_),
    .A2(_03291_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11181_ (.A1(_03267_),
    .A2(_03204_),
    .A3(_03292_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _11182_ (.I(_03293_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 _11183_ (.I(_03294_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11184_ (.I0(_07604_),
    .I1(_03127_),
    .S(_03295_),
    .Z(_07630_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11185_ (.A1(_07502_),
    .A2(_02899_),
    .ZN(_07521_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11186_ (.A1(_07523_),
    .A2(_07525_),
    .A3(_07524_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11187_ (.A1(_02703_),
    .A2(_03296_),
    .Z(_03297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11188_ (.I0(_07521_),
    .I1(_03297_),
    .S(_02844_),
    .Z(_07546_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11189_ (.A1(_07548_),
    .A2(_02855_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11190_ (.I0(_07546_),
    .I1(_03298_),
    .S(_03006_),
    .Z(_07567_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11191_ (.A1(_07569_),
    .A2(_03011_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11192_ (.I0(_07567_),
    .I1(_03299_),
    .S(_03115_),
    .Z(_07598_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11193_ (.A1(_07600_),
    .A2(_03122_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11194_ (.I0(_07598_),
    .I1(_03300_),
    .S(_03295_),
    .Z(_07618_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11195_ (.I(_07614_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11196_ (.A1(_07617_),
    .A2(_07616_),
    .B(_07615_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11197_ (.A1(_03301_),
    .A2(_03302_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11198_ (.A1(_03303_),
    .A2(_07629_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11199_ (.A1(_03304_),
    .A2(_07628_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11200_ (.A1(_07626_),
    .A2(_03305_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11201_ (.A1(_03306_),
    .A2(_07625_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11202_ (.A1(_07623_),
    .A2(_03307_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11203_ (.A1(_07622_),
    .A2(_03308_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11204_ (.A1(_07620_),
    .A2(_03309_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11205_ (.I(_03267_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11206_ (.I(_03292_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11207_ (.I0(_07555_),
    .I1(_03226_),
    .S(net12),
    .Z(_07578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11208_ (.I0(_03215_),
    .I1(_07578_),
    .S(_03202_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11209_ (.A1(_07610_),
    .A2(_03313_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _11210_ (.A1(_03204_),
    .A2(_03311_),
    .A3(_03312_),
    .A4(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11211_ (.A1(_07612_),
    .A2(net386),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11212_ (.A1(_03214_),
    .A2(_03313_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11213_ (.A1(_03214_),
    .A2(_03313_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _11214_ (.A1(_03316_),
    .A2(_03317_),
    .A3(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11215_ (.I(_03319_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11216_ (.A1(_07615_),
    .A2(_07623_),
    .A3(_07626_),
    .A4(net391),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11217_ (.A1(_07620_),
    .A2(_07617_),
    .A3(_07632_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11218_ (.A1(_07635_),
    .A2(_07769_),
    .A3(_03321_),
    .A4(_03322_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11219_ (.A1(_03315_),
    .A2(_03320_),
    .B(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11220_ (.A1(_03141_),
    .A2(_03183_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11221_ (.A1(_03202_),
    .A2(_03201_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11222_ (.A1(_03166_),
    .A2(_03169_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11223_ (.A1(_03202_),
    .A2(_03232_),
    .A3(_03196_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11224_ (.A1(_03327_),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11225_ (.A1(_03203_),
    .A2(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11226_ (.A1(_03326_),
    .A2(_03311_),
    .A3(_03312_),
    .B(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11227_ (.A1(_03325_),
    .A2(_03331_),
    .Z(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11228_ (.A1(_03141_),
    .A2(_03183_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11229_ (.A1(_03202_),
    .A2(_03201_),
    .B(_03203_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11230_ (.A1(_03333_),
    .A2(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11231_ (.A1(_03166_),
    .A2(_03328_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11232_ (.A1(_03198_),
    .A2(_03336_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11233_ (.A1(_03335_),
    .A2(_03311_),
    .A3(_03312_),
    .B(_03337_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11234_ (.A1(_03335_),
    .A2(_03311_),
    .A3(_03312_),
    .A4(_03337_),
    .Z(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11235_ (.A1(_03087_),
    .A2(_03106_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11236_ (.I(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _11237_ (.A1(_03341_),
    .A2(_03169_),
    .B1(_03327_),
    .B2(_03328_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11238_ (.A1(_03338_),
    .A2(_03339_),
    .B(_03291_),
    .C(_03342_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _11239_ (.A1(_03324_),
    .A2(_03332_),
    .A3(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11240_ (.I(_03344_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11241_ (.A1(net383),
    .A2(_03238_),
    .A3(_03266_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11242_ (.I(_03270_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11243_ (.A1(_03233_),
    .A2(_03237_),
    .Z(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11244_ (.A1(_03248_),
    .A2(_03240_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11245_ (.A1(net378),
    .A2(_03349_),
    .B(_03264_),
    .C(_03252_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11246_ (.A1(_03208_),
    .A2(net377),
    .A3(_03243_),
    .A4(_03350_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11247_ (.A1(_03239_),
    .A2(_03233_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _11248_ (.A1(_03269_),
    .A2(_03348_),
    .A3(_03351_),
    .A4(_03352_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11249_ (.A1(_03346_),
    .A2(_03347_),
    .B(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11250_ (.A1(net376),
    .A2(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11251_ (.A1(_03334_),
    .A2(_03238_),
    .A3(_03266_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11252_ (.A1(_03348_),
    .A2(_03351_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11253_ (.A1(_03333_),
    .A2(_03312_),
    .A3(_03356_),
    .B(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11254_ (.A1(_03204_),
    .A2(_03270_),
    .A3(_03291_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11255_ (.A1(_03348_),
    .A2(_03351_),
    .B(_03352_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11256_ (.A1(_03346_),
    .A2(_03359_),
    .B(_03360_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11257_ (.A1(_03348_),
    .A2(_03351_),
    .B(_03358_),
    .C(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11258_ (.A1(_03355_),
    .A2(_03362_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11259_ (.I(_03363_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11260_ (.A1(_03204_),
    .A2(_03311_),
    .A3(_03292_),
    .A4(_03314_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11261_ (.A1(_07620_),
    .A2(_03309_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11262_ (.A1(_07619_),
    .A2(_03366_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11263_ (.A1(_07635_),
    .A2(_03367_),
    .Z(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11264_ (.A1(_07634_),
    .A2(_03368_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11265_ (.A1(_03369_),
    .A2(_07632_),
    .Z(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11266_ (.A1(_03370_),
    .A2(_07631_),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11267_ (.A1(_03365_),
    .A2(_03319_),
    .B(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11268_ (.A1(_03333_),
    .A2(_03312_),
    .A3(_03356_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11269_ (.A1(_03263_),
    .A2(_03234_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11270_ (.A1(_03177_),
    .A2(net39),
    .A3(_03240_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11271_ (.A1(_03374_),
    .A2(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11272_ (.I(_03376_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11273_ (.A1(_03060_),
    .A2(_03240_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11274_ (.A1(net39),
    .A2(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11275_ (.A1(_02991_),
    .A2(_03052_),
    .A3(_03055_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11276_ (.A1(_02992_),
    .A2(_03056_),
    .B(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11277_ (.I(_03255_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11278_ (.A1(net39),
    .A2(_03382_),
    .A3(_03257_),
    .A4(_03378_),
    .Z(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _11279_ (.A1(_03258_),
    .A2(_03379_),
    .B1(_03381_),
    .B2(_03044_),
    .C(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11280_ (.A1(_03108_),
    .A2(_03349_),
    .B(_03252_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11281_ (.A1(net12),
    .A2(_03044_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11282_ (.A1(_03386_),
    .A2(_03262_),
    .Z(_03387_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11283_ (.A1(_03385_),
    .A2(_03387_),
    .A3(_03379_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11284_ (.A1(_03208_),
    .A2(net377),
    .A3(_03243_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11285_ (.A1(net12),
    .A2(_03384_),
    .B(_03388_),
    .C(_03389_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11286_ (.A1(_03204_),
    .A2(_03311_),
    .A3(_03312_),
    .B(_03390_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11287_ (.A1(_03351_),
    .A2(_03373_),
    .B1(_03377_),
    .B2(_03391_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11288_ (.A1(_03044_),
    .A2(_03255_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11289_ (.A1(net12),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11290_ (.A1(_03379_),
    .A2(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11291_ (.A1(_03389_),
    .A2(_03388_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11292_ (.A1(_03204_),
    .A2(_03311_),
    .A3(_03292_),
    .B(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11293_ (.A1(_03395_),
    .A2(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11294_ (.I(_03385_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _11295_ (.A1(_03210_),
    .A2(_03216_),
    .B1(net381),
    .B2(net39),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11296_ (.A1(net47),
    .A2(_03210_),
    .A3(_03216_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11297_ (.A1(_03050_),
    .A2(_03099_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11298_ (.I(_03243_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11299_ (.A1(_03402_),
    .A2(_03403_),
    .B(net47),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11300_ (.A1(_03208_),
    .A2(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _11301_ (.A1(_03399_),
    .A2(_03400_),
    .A3(_03401_),
    .A4(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11302_ (.I(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11303_ (.A1(_03074_),
    .A2(_03256_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11304_ (.A1(_03060_),
    .A2(_03240_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11305_ (.A1(_03386_),
    .A2(_03409_),
    .B(_03382_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11306_ (.A1(_03408_),
    .A2(_03410_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11307_ (.A1(net47),
    .A2(_03411_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11308_ (.A1(net47),
    .A2(_03349_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11309_ (.A1(_03413_),
    .A2(_03387_),
    .B(_03379_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11310_ (.A1(_03294_),
    .A2(_03407_),
    .B(_03412_),
    .C(_03414_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _11311_ (.A1(_03415_),
    .A2(_03392_),
    .A3(_03398_),
    .A4(_03372_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11312_ (.A1(_03416_),
    .A2(_03364_),
    .A3(_03345_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11313_ (.I0(_07618_),
    .I1(_03310_),
    .S(net10),
    .Z(_07648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11314_ (.A1(_03294_),
    .A2(_03400_),
    .B(_03401_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _11315_ (.A1(_03392_),
    .A2(_03398_),
    .A3(_03415_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11316_ (.A1(_03345_),
    .A2(_03364_),
    .A3(_03419_),
    .B(_03372_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11317_ (.A1(_03418_),
    .A2(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11318_ (.A1(net39),
    .A2(_03402_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11319_ (.A1(net12),
    .A2(_03206_),
    .B(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11320_ (.A1(_03207_),
    .A2(_03400_),
    .B(_03422_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11321_ (.A1(_03070_),
    .A2(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11322_ (.A1(_03243_),
    .A2(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11323_ (.A1(net37),
    .A2(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11324_ (.A1(_03372_),
    .A2(_03418_),
    .A3(_03423_),
    .A4(_03427_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11325_ (.A1(_03344_),
    .A2(_03363_),
    .A3(_03416_),
    .B(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11326_ (.A1(_03311_),
    .A2(_03204_),
    .A3(_03312_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11327_ (.A1(_03430_),
    .A2(_03389_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _11328_ (.A1(_03385_),
    .A2(_03429_),
    .A3(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11329_ (.A1(_03421_),
    .A2(_03432_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11330_ (.A1(_03345_),
    .A2(_03364_),
    .A3(_03419_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11331_ (.I(_03423_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11332_ (.A1(_03372_),
    .A2(_03418_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11333_ (.A1(_03435_),
    .A2(_03436_),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11334_ (.A1(_03207_),
    .A2(net37),
    .A3(_03400_),
    .Z(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11335_ (.A1(_03422_),
    .A2(_03438_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11336_ (.A1(_03070_),
    .A2(_03439_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11337_ (.A1(net47),
    .A2(_03231_),
    .A3(_03244_),
    .Z(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11338_ (.A1(_03431_),
    .A2(_03441_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11339_ (.A1(_03434_),
    .A2(_03437_),
    .A3(_03440_),
    .B(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11340_ (.A1(_03434_),
    .A2(_03437_),
    .A3(_03442_),
    .A4(_03440_),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11341_ (.A1(net370),
    .A2(_03317_),
    .B(_03318_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11342_ (.A1(_03207_),
    .A2(net46),
    .Z(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11343_ (.I0(_03435_),
    .I1(_03446_),
    .S(_03400_),
    .Z(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11344_ (.A1(_03440_),
    .A2(_03445_),
    .A3(_03447_),
    .Z(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11345_ (.A1(_03443_),
    .A2(_03444_),
    .B(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11346_ (.A1(_07630_),
    .A2(net10),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11347_ (.I(_07610_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11348_ (.I0(_03451_),
    .I1(_03316_),
    .S(net37),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11349_ (.A1(_07631_),
    .A2(_03452_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11350_ (.A1(_07632_),
    .A2(_03369_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11351_ (.A1(_03370_),
    .A2(_03452_),
    .B1(_03453_),
    .B2(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11352_ (.A1(_07631_),
    .A2(_03370_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11353_ (.A1(_03315_),
    .A2(_03320_),
    .B(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11354_ (.A1(_07500_),
    .A2(_02770_),
    .ZN(_07518_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11355_ (.A1(_07502_),
    .A2(_07520_),
    .A3(_07501_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11356_ (.A1(_02552_),
    .A2(_03458_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11357_ (.I0(_07518_),
    .I1(_03459_),
    .S(_02701_),
    .Z(_07541_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11358_ (.A1(_07543_),
    .A2(_02704_),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11359_ (.I0(_07541_),
    .I1(_03460_),
    .S(_02844_),
    .Z(_07564_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11360_ (.A1(_07566_),
    .A2(_02857_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11361_ (.I0(_07564_),
    .I1(_03461_),
    .S(_03006_),
    .Z(_07587_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11362_ (.A1(_07589_),
    .A2(_03013_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11363_ (.I0(_07587_),
    .I1(_03462_),
    .S(_03115_),
    .Z(_07607_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11364_ (.A1(_07609_),
    .A2(net389),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11365_ (.I0(_07607_),
    .I1(_03463_),
    .S(net374),
    .Z(_07633_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11366_ (.A1(_03457_),
    .A2(_07633_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11367_ (.A1(_03344_),
    .A2(_03364_),
    .A3(_03419_),
    .A4(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11368_ (.A1(_07635_),
    .A2(_03367_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _11369_ (.A1(_03345_),
    .A2(_03364_),
    .A3(_03416_),
    .B1(_03466_),
    .B2(_03368_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11370_ (.I(_07653_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11371_ (.I(_07658_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11372_ (.I(_07646_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11373_ (.A1(_07639_),
    .A2(_07640_),
    .B(_07647_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11374_ (.A1(_03471_),
    .A2(_03470_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11375_ (.A1(_03472_),
    .A2(_07644_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11376_ (.A1(_03473_),
    .A2(_07643_),
    .B(_07659_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11377_ (.A1(_03474_),
    .A2(_03469_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11378_ (.A1(_03475_),
    .A2(_07656_),
    .B(_07655_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11379_ (.I(_07652_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11380_ (.A1(_03476_),
    .A2(_03468_),
    .B(_03477_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11381_ (.A1(_03478_),
    .A2(_07650_),
    .B(_07649_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11382_ (.A1(_07177_),
    .A2(_03479_),
    .B(_02196_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11383_ (.A1(_03480_),
    .A2(_03467_),
    .A3(_03465_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11384_ (.A1(_03465_),
    .A2(_03467_),
    .B(_03479_),
    .C(_02507_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11385_ (.A1(_03450_),
    .A2(_03455_),
    .B(_03482_),
    .C(_03481_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11386_ (.A1(_03483_),
    .A2(_03449_),
    .A3(_03433_),
    .Z(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11387_ (.A1(net46),
    .A2(_03407_),
    .B(_03457_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _11388_ (.A1(_03345_),
    .A2(_03364_),
    .A3(_03416_),
    .B(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11389_ (.A1(_03385_),
    .A2(_03431_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11390_ (.A1(_03486_),
    .A2(_03487_),
    .B(_03414_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11391_ (.A1(_03414_),
    .A2(_03486_),
    .A3(_03487_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11392_ (.A1(_03346_),
    .A2(_03359_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11393_ (.A1(_03360_),
    .A2(_03490_),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11394_ (.A1(_03348_),
    .A2(_03351_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11395_ (.A1(_03373_),
    .A2(_03357_),
    .B(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11396_ (.A1(_03372_),
    .A2(_03392_),
    .A3(_03398_),
    .A4(_03415_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11397_ (.A1(_03493_),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11398_ (.A1(_03324_),
    .A2(_03332_),
    .A3(_03343_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11399_ (.A1(net46),
    .A2(_03354_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11400_ (.A1(_03493_),
    .A2(_03372_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11401_ (.A1(_03496_),
    .A2(_03497_),
    .B(_03419_),
    .C(_03498_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11402_ (.A1(_03491_),
    .A2(_03495_),
    .A3(_03499_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11403_ (.A1(_03395_),
    .A2(_03397_),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11404_ (.I(_03412_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11405_ (.A1(net46),
    .A2(_03396_),
    .A3(_03395_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11406_ (.A1(_03502_),
    .A2(_03503_),
    .B(_03391_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11407_ (.A1(_03377_),
    .A2(_03504_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11408_ (.A1(_03203_),
    .A2(_03329_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11409_ (.A1(_03506_),
    .A2(_03137_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11410_ (.A1(_03138_),
    .A2(_03506_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11411_ (.A1(_03028_),
    .A2(_03508_),
    .B(_03507_),
    .C(_02877_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11412_ (.A1(_03334_),
    .A2(_03311_),
    .A3(_03312_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11413_ (.I0(_03507_),
    .I1(_03509_),
    .S(_03510_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11414_ (.I(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11415_ (.A1(_03501_),
    .A2(_03505_),
    .A3(_03512_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11416_ (.A1(_03488_),
    .A2(_03489_),
    .A3(_03500_),
    .A4(_03513_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11417_ (.A1(net372),
    .A2(_03353_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11418_ (.A1(_03280_),
    .A2(_03515_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11419_ (.A1(_03282_),
    .A2(_03290_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11420_ (.A1(_03280_),
    .A2(net371),
    .A3(_03353_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11421_ (.A1(_03517_),
    .A2(_03518_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11422_ (.A1(_03355_),
    .A2(_03362_),
    .A3(_03457_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11423_ (.A1(_07631_),
    .A2(_03430_),
    .A3(_03406_),
    .B(_03371_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _11424_ (.A1(_03365_),
    .A2(_03319_),
    .B1(_03373_),
    .B2(_03357_),
    .C(_03492_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11425_ (.A1(net37),
    .A2(_03354_),
    .B(_03280_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11426_ (.A1(_03361_),
    .A2(_03521_),
    .A3(_03522_),
    .A4(_03523_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11427_ (.A1(_03392_),
    .A2(_03398_),
    .A3(_03415_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11428_ (.A1(_03344_),
    .A2(_03520_),
    .B(_03524_),
    .C(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11429_ (.A1(_03519_),
    .A2(_03526_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11430_ (.A1(_03345_),
    .A2(_03497_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11431_ (.A1(_03362_),
    .A2(_03457_),
    .A3(_03419_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11432_ (.I0(_03528_),
    .I1(_03355_),
    .S(_03529_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11433_ (.A1(_03338_),
    .A2(_03339_),
    .Z(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11434_ (.A1(_03342_),
    .A2(_03531_),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11435_ (.A1(_03157_),
    .A2(_03282_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11436_ (.A1(_03328_),
    .A2(_03533_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11437_ (.A1(_03517_),
    .A2(_03518_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11438_ (.A1(_03534_),
    .A2(_03535_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11439_ (.A1(_03532_),
    .A2(_03536_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11440_ (.A1(_03516_),
    .A2(_03527_),
    .A3(_03530_),
    .A4(_03537_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11441_ (.A1(_03333_),
    .A2(_03510_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11442_ (.A1(_03331_),
    .A2(_03539_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _11443_ (.A1(_07635_),
    .A2(_07769_),
    .A3(_03321_),
    .A4(_03322_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11444_ (.A1(_03365_),
    .A2(_03319_),
    .B(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11445_ (.A1(_03325_),
    .A2(_03331_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11446_ (.A1(_03542_),
    .A2(_03543_),
    .B(_03343_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11447_ (.A1(_03497_),
    .A2(_03361_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _11448_ (.A1(_03419_),
    .A2(_03498_),
    .A3(_03544_),
    .A4(_03545_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11449_ (.A1(_03540_),
    .A2(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11450_ (.A1(_03519_),
    .A2(_03534_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11451_ (.I(_03507_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11452_ (.A1(_03532_),
    .A2(_03549_),
    .A3(_03540_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11453_ (.A1(_03028_),
    .A2(_03508_),
    .B(_02877_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11454_ (.A1(_03510_),
    .A2(_03507_),
    .B(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _11455_ (.A1(_03526_),
    .A2(_03548_),
    .A3(_03550_),
    .B(_03552_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11456_ (.A1(_03547_),
    .A2(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11457_ (.A1(_03514_),
    .A2(_03538_),
    .A3(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11458_ (.A1(_03555_),
    .A2(_03484_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11459_ (.I(_03556_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11460_ (.A1(_07650_),
    .A2(_03478_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11461_ (.A1(_03557_),
    .A2(_03558_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11462_ (.A1(_07648_),
    .A2(net16),
    .B(_03559_),
    .ZN(_07661_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11463_ (.A1(_07525_),
    .A2(_03033_),
    .ZN(_07549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11464_ (.A1(_07545_),
    .A2(_07551_),
    .A3(_07544_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11465_ (.A1(_02854_),
    .A2(_03560_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11466_ (.I0(_07549_),
    .I1(_03561_),
    .S(_03006_),
    .Z(_07570_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11467_ (.A1(_07572_),
    .A2(_03009_),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11468_ (.I0(_07570_),
    .I1(_03562_),
    .S(_03115_),
    .Z(_07601_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11469_ (.A1(_07603_),
    .A2(_03120_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11470_ (.I0(_07601_),
    .I1(_03563_),
    .S(net401),
    .Z(_07621_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11471_ (.A1(_07623_),
    .A2(_03307_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11472_ (.I0(_07621_),
    .I1(_03564_),
    .S(_03417_),
    .Z(_07651_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11473_ (.I(_07643_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11474_ (.I(_07647_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11475_ (.A1(_03566_),
    .A2(_07638_),
    .B(_03470_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11476_ (.A1(_07644_),
    .A2(_03567_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11477_ (.A1(_03565_),
    .A2(_03568_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11478_ (.A1(_07659_),
    .A2(_03569_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11479_ (.A1(_07658_),
    .A2(_03570_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11480_ (.A1(_07656_),
    .A2(_03571_),
    .B(_07655_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11481_ (.A1(_03468_),
    .A2(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11482_ (.A1(_03557_),
    .A2(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11483_ (.A1(_03557_),
    .A2(_07651_),
    .B(_03574_),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11484_ (.A1(_07545_),
    .A2(_03253_),
    .ZN(_07573_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11485_ (.A1(_07577_),
    .A2(_07575_),
    .A3(_07576_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11486_ (.A1(_03008_),
    .A2(_03575_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11487_ (.I0(_07573_),
    .I1(_03576_),
    .S(_03115_),
    .Z(_07592_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11488_ (.A1(_07594_),
    .A2(_03118_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11489_ (.I0(_07592_),
    .I1(_03577_),
    .S(net401),
    .Z(_07624_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11490_ (.A1(_07626_),
    .A2(net388),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11491_ (.I0(_07624_),
    .I1(_03578_),
    .S(_03417_),
    .Z(_07654_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11492_ (.A1(_07656_),
    .A2(_03475_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11493_ (.A1(_03579_),
    .A2(_03557_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11494_ (.A1(net16),
    .A2(_07654_),
    .B(_03580_),
    .ZN(_07669_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11495_ (.A1(_07577_),
    .A2(_03202_),
    .ZN(_07595_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11496_ (.A1(_07597_),
    .A2(_07591_),
    .A3(_07590_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11497_ (.A1(_03117_),
    .A2(_03581_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11498_ (.I0(_07595_),
    .I1(_03582_),
    .S(_03295_),
    .Z(_07627_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _11499_ (.A1(net382),
    .A2(_03303_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11500_ (.I0(net379),
    .I1(_03583_),
    .S(_03417_),
    .Z(_07657_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11501_ (.A1(_07659_),
    .A2(_03569_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11502_ (.A1(_03570_),
    .A2(_03584_),
    .B(_03557_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11503_ (.A1(net16),
    .A2(_07657_),
    .B(_03585_),
    .ZN(_07673_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11504_ (.A1(_07591_),
    .A2(_03430_),
    .ZN(_07613_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11505_ (.A1(_07615_),
    .A2(_07617_),
    .A3(_07616_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11506_ (.A1(_03302_),
    .A2(_03586_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11507_ (.I0(_07613_),
    .I1(_03587_),
    .S(_03417_),
    .Z(_07642_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11508_ (.A1(_07644_),
    .A2(_03472_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11509_ (.A1(_03473_),
    .A2(_03588_),
    .B(net16),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11510_ (.A1(net16),
    .A2(_07642_),
    .B(_03589_),
    .ZN(_07677_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11511_ (.I(_07617_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11512_ (.I0(\butterfly_count[2] ),
    .I1(_03590_),
    .S(_03417_),
    .Z(_07645_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _11513_ (.I(_05877_),
    .ZN(_05862_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11514_ (.I(\state[0] ),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11515_ (.A1(net80),
    .A2(_07803_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11516_ (.A1(\state[2] ),
    .A2(_03592_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11517_ (.A1(_03591_),
    .A2(_00565_),
    .B(_03593_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _11518_ (.I(\state[1] ),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11519_ (.I(_03594_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11520_ (.I(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11521_ (.A1(\state[2] ),
    .A2(net80),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11522_ (.A1(_03596_),
    .A2(_07789_),
    .B1(_03597_),
    .B2(_07803_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11523_ (.I(_03598_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11524_ (.I(\idx1[1] ),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11525_ (.I(_03599_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11526_ (.I(\idx1[2] ),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11527_ (.I(\idx1[0] ),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11528_ (.A1(_03601_),
    .A2(_03602_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11529_ (.I(_03602_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11530_ (.A1(\idx1[2] ),
    .A2(_03604_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11531_ (.A1(\samples_real[3][0] ),
    .A2(_03603_),
    .B1(_03605_),
    .B2(\samples_real[6][0] ),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11532_ (.A1(_03600_),
    .A2(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11533_ (.I0(\samples_real[4][0] ),
    .I1(\samples_real[5][0] ),
    .S(_03602_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11534_ (.I(_03602_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11535_ (.A1(_03609_),
    .A2(\samples_real[7][0] ),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11536_ (.I(\idx1[1] ),
    .Z(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11537_ (.I0(_03608_),
    .I1(_03610_),
    .S(_03611_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11538_ (.I(_03609_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11539_ (.I(\samples_real[1][0] ),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11540_ (.A1(_03604_),
    .A2(\samples_real[2][0] ),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11541_ (.A1(_03613_),
    .A2(_03614_),
    .B1(_03615_),
    .B2(_03611_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11542_ (.I(_03601_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11543_ (.I0(_03612_),
    .I1(_03616_),
    .S(_03617_),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11544_ (.A1(_03599_),
    .A2(_03604_),
    .Z(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11545_ (.A1(_03601_),
    .A2(_03619_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11546_ (.A1(_03607_),
    .A2(_03618_),
    .B1(_03620_),
    .B2(\samples_real[0][0] ),
    .ZN(_07704_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11547_ (.I0(\samples_real[4][1] ),
    .I1(\samples_real[5][1] ),
    .I2(\samples_real[6][1] ),
    .I3(\samples_real[7][1] ),
    .S0(_03609_),
    .S1(_03611_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11548_ (.I(_03611_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11549_ (.I0(\samples_real[2][1] ),
    .I1(\samples_real[3][1] ),
    .S(_03609_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11550_ (.I(_03623_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11551_ (.A1(_03599_),
    .A2(_03602_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11552_ (.I(_03625_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11553_ (.I(\samples_real[1][1] ),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11554_ (.A1(_03622_),
    .A2(_03624_),
    .B1(_03626_),
    .B2(_03627_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11555_ (.I0(_03621_),
    .I1(_03628_),
    .S(_03601_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11556_ (.A1(\samples_real[0][1] ),
    .A2(_03620_),
    .B(_03629_),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _11557_ (.I(\temp_real[0] ),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11558_ (.I(_05861_),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11559_ (.I(\stage[1] ),
    .ZN(_07774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11560_ (.I0(\butterfly_in_group[0] ),
    .I1(\butterfly_in_group[1] ),
    .S(\stage[0] ),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11561_ (.A1(_07787_),
    .A2(\stage[1] ),
    .A3(_03630_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _11562_ (.I(\stage[0] ),
    .ZN(_07773_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11563_ (.A1(_00567_),
    .A2(_07773_),
    .A3(\butterfly_in_group[2] ),
    .A4(_07774_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11564_ (.A1(_03631_),
    .A2(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11565_ (.A1(_00581_),
    .A2(_03594_),
    .Z(_03634_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11566_ (.A1(_07789_),
    .A2(net81),
    .A3(_03634_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11567_ (.I(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _11568_ (.I0(\twiddle_idx[0] ),
    .I1(_03633_),
    .S(_03636_),
    .Z(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11569_ (.I0(\butterfly_in_group[0] ),
    .I1(\butterfly_in_group[2] ),
    .S(\stage[1] ),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11570_ (.A1(\butterfly_in_group[1] ),
    .A2(\stage[1] ),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11571_ (.I0(_03637_),
    .I1(_03638_),
    .S(_07773_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11572_ (.A1(_07787_),
    .A2(_03639_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _11573_ (.I0(\twiddle_idx[1] ),
    .I1(_03640_),
    .S(_03636_),
    .Z(_00007_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11574_ (.A1(_00000_),
    .A2(_00007_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11575_ (.I(_00021_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11576_ (.A1(_00000_),
    .A2(_00007_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11577_ (.A1(_00018_),
    .A2(_00020_),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11578_ (.I(_00007_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11579_ (.I(_03620_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11580_ (.I(_03613_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11581_ (.I(_03642_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11582_ (.I(_03622_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11583_ (.I(_03644_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11584_ (.I0(\samples_imag[4][0] ),
    .I1(\samples_imag[5][0] ),
    .I2(\samples_imag[6][0] ),
    .I3(\samples_imag[7][0] ),
    .S0(_03643_),
    .S1(_03645_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11585_ (.I(\samples_imag[1][0] ),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11586_ (.I(_03626_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11587_ (.I(_03609_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11588_ (.I(_03649_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11589_ (.I0(\samples_imag[2][0] ),
    .I1(\samples_imag[3][0] ),
    .S(_03650_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11590_ (.I(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11591_ (.A1(_03647_),
    .A2(_03648_),
    .B1(_03652_),
    .B2(_03645_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11592_ (.I(_03617_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11593_ (.I(_03654_),
    .Z(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11594_ (.I0(_03646_),
    .I1(_03653_),
    .S(_03655_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11595_ (.A1(\samples_imag[0][0] ),
    .A2(_03641_),
    .B(_03656_),
    .ZN(_07818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11596_ (.A1(\samples_imag[3][1] ),
    .A2(_03603_),
    .B1(_03605_),
    .B2(\samples_imag[6][1] ),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11597_ (.A1(_03600_),
    .A2(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11598_ (.I0(\samples_imag[4][1] ),
    .I1(\samples_imag[5][1] ),
    .S(_03642_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11599_ (.A1(_03650_),
    .A2(\samples_imag[7][1] ),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11600_ (.I(_03622_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11601_ (.I0(_03659_),
    .I1(_03660_),
    .S(_03661_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11602_ (.I(\samples_imag[1][1] ),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11603_ (.I(_03604_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11604_ (.I(_03664_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11605_ (.A1(_03665_),
    .A2(\samples_imag[2][1] ),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11606_ (.A1(_03643_),
    .A2(_03663_),
    .B1(_03666_),
    .B2(_03645_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11607_ (.I0(_03662_),
    .I1(_03667_),
    .S(_03655_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _11608_ (.A1(\samples_imag[0][1] ),
    .A2(_03641_),
    .B1(_03658_),
    .B2(_03668_),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _11609_ (.I(\temp_imag[0] ),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11610_ (.I(_05876_),
    .ZN(_05873_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11611_ (.A1(_07787_),
    .A2(_07773_),
    .A3(_07774_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11612_ (.A1(\group[0] ),
    .A2(_02507_),
    .A3(_03669_),
    .Z(_07883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11613_ (.A1(\group[1] ),
    .A2(_02507_),
    .A3(_03669_),
    .Z(_07885_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11614_ (.I(_07790_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11615_ (.A1(\group[0] ),
    .A2(_07777_),
    .A3(_03670_),
    .A4(_03669_),
    .Z(_07888_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11616_ (.I(\idx2[1] ),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11617_ (.I(_03671_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11618_ (.I(_03672_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11619_ (.I(\idx2[0] ),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11620_ (.I(_03674_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11621_ (.I(_03675_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11622_ (.I(\idx2[2] ),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11623_ (.I(_03677_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11624_ (.I(_03678_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11625_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11626_ (.I0(\samples_real[2][12] ),
    .I1(\samples_real[3][12] ),
    .I2(\samples_real[6][12] ),
    .I3(\samples_real[7][12] ),
    .S0(_03676_),
    .S1(_03680_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11627_ (.A1(_03673_),
    .A2(_03681_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11628_ (.I(_03674_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11629_ (.I(_03683_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11630_ (.I(_03684_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11631_ (.I0(\samples_real[1][12] ),
    .I1(\samples_real[5][12] ),
    .S(_03680_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11632_ (.I(_03677_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11633_ (.I(_03687_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11634_ (.I(_03688_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11635_ (.A1(_03676_),
    .A2(_03689_),
    .A3(\samples_real[4][12] ),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11636_ (.I(\idx2[1] ),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11637_ (.I(_03691_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11638_ (.I(_03692_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11639_ (.A1(_03685_),
    .A2(_03686_),
    .B(_03690_),
    .C(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11640_ (.A1(_03683_),
    .A2(_03687_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11641_ (.I(_03695_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11642_ (.A1(_03692_),
    .A2(_03696_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _11643_ (.I(_03697_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11644_ (.I(\samples_real[0][12] ),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11645_ (.A1(_03682_),
    .A2(_03694_),
    .B1(_03698_),
    .B2(_03699_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11646_ (.A1(_00010_),
    .A2(_03700_),
    .ZN(_05917_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11647_ (.A1(_03688_),
    .A2(\samples_imag[4][12] ),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11648_ (.A1(_03689_),
    .A2(\samples_imag[1][12] ),
    .B1(_03701_),
    .B2(_03684_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11649_ (.A1(_03691_),
    .A2(_03678_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11650_ (.A1(_03671_),
    .A2(_03687_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11651_ (.A1(\samples_imag[5][12] ),
    .A2(_03703_),
    .B1(_03704_),
    .B2(\samples_imag[3][12] ),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11652_ (.A1(\idx2[1] ),
    .A2(_03677_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11653_ (.I(_03706_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11654_ (.I0(\samples_imag[6][12] ),
    .I1(\samples_imag[7][12] ),
    .S(_03675_),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11655_ (.A1(\samples_imag[2][12] ),
    .A2(_03696_),
    .B1(_03707_),
    .B2(_03708_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11656_ (.A1(_03672_),
    .A2(_03702_),
    .B1(_03705_),
    .B2(_03684_),
    .C(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11657_ (.A1(_03692_),
    .A2(_03695_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _11658_ (.I(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11659_ (.A1(\samples_imag[0][12] ),
    .A2(_03712_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11660_ (.A1(_03710_),
    .A2(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11661_ (.A1(_00008_),
    .A2(_03714_),
    .Z(_07908_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _11662_ (.I(_00010_),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11663_ (.A1(\samples_real[5][11] ),
    .A2(_03703_),
    .B1(_03704_),
    .B2(\samples_real[3][11] ),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11664_ (.I(_03687_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11665_ (.A1(_03687_),
    .A2(\samples_real[4][11] ),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11666_ (.A1(_03717_),
    .A2(\samples_real[1][11] ),
    .B1(_03718_),
    .B2(_03683_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11667_ (.I0(\samples_real[6][11] ),
    .I1(\samples_real[7][11] ),
    .S(_03674_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11668_ (.A1(\samples_real[2][11] ),
    .A2(_03696_),
    .B1(_03706_),
    .B2(_03720_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11669_ (.A1(_03684_),
    .A2(_03716_),
    .B1(_03719_),
    .B2(_03671_),
    .C(_03721_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11670_ (.A1(\samples_real[0][11] ),
    .A2(_03711_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11671_ (.A1(_03722_),
    .A2(_03723_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11672_ (.A1(_03715_),
    .A2(_03724_),
    .Z(_05922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11673_ (.I(_05922_),
    .ZN(_05881_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11674_ (.I(_00008_),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11675_ (.I(_03725_),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11676_ (.I(\samples_imag[0][11] ),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _11677_ (.I(_03698_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _11678_ (.I(_03676_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11679_ (.I(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11680_ (.I(_03680_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11681_ (.I0(\samples_imag[2][11] ),
    .I1(\samples_imag[3][11] ),
    .I2(\samples_imag[6][11] ),
    .I3(\samples_imag[7][11] ),
    .S0(_03730_),
    .S1(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11682_ (.A1(_03673_),
    .A2(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11683_ (.I0(\samples_imag[1][11] ),
    .I1(\samples_imag[5][11] ),
    .S(_03731_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11684_ (.I(_03689_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11685_ (.A1(_03730_),
    .A2(_03735_),
    .A3(\samples_imag[4][11] ),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11686_ (.I(_03693_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11687_ (.A1(_03685_),
    .A2(_03734_),
    .B(_03736_),
    .C(_03737_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11688_ (.A1(_03727_),
    .A2(_03728_),
    .B1(_03733_),
    .B2(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11689_ (.A1(_03726_),
    .A2(_03739_),
    .Z(_05882_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11690_ (.I(_03725_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11691_ (.I(\samples_imag[0][10] ),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11692_ (.I0(\samples_imag[3][10] ),
    .I1(\samples_imag[7][10] ),
    .S(_03731_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11693_ (.A1(_03673_),
    .A2(_03730_),
    .A3(_03742_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11694_ (.I0(\samples_imag[4][10] ),
    .I1(\samples_imag[5][10] ),
    .S(_03729_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11695_ (.A1(_03671_),
    .A2(_03683_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11696_ (.A1(_03737_),
    .A2(_03744_),
    .B1(_03745_),
    .B2(\samples_imag[6][10] ),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11697_ (.A1(_03685_),
    .A2(\samples_imag[2][10] ),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11698_ (.A1(_03685_),
    .A2(\samples_imag[1][10] ),
    .B1(_03747_),
    .B2(_03737_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11699_ (.I0(_03746_),
    .I1(_03748_),
    .S(_03735_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11700_ (.A1(_03741_),
    .A2(_03728_),
    .B1(_03743_),
    .B2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11701_ (.A1(_03740_),
    .A2(_03750_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11702_ (.I(_05891_),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11703_ (.I(\samples_imag[0][9] ),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11704_ (.A1(_03674_),
    .A2(_03706_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11705_ (.I(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11706_ (.A1(_03691_),
    .A2(_03674_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11707_ (.A1(_03687_),
    .A2(_03754_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11708_ (.A1(\samples_imag[7][9] ),
    .A2(_03753_),
    .B1(_03755_),
    .B2(\samples_imag[1][9] ),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11709_ (.A1(_03683_),
    .A2(_03677_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11710_ (.I(_03757_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11711_ (.A1(_03691_),
    .A2(_03758_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11712_ (.I(_03759_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11713_ (.A1(\idx2[1] ),
    .A2(_03695_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11714_ (.I(_03761_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11715_ (.A1(\samples_imag[4][9] ),
    .A2(_03760_),
    .B1(_03762_),
    .B2(\samples_imag[2][9] ),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11716_ (.A1(_03674_),
    .A2(_03687_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11717_ (.A1(\samples_imag[6][9] ),
    .A2(_03758_),
    .B1(_03764_),
    .B2(\samples_imag[3][9] ),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11718_ (.A1(_03674_),
    .A2(_03678_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11719_ (.I(_03766_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11720_ (.A1(\samples_imag[5][9] ),
    .A2(_03767_),
    .B(_03696_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11721_ (.I0(_03765_),
    .I1(_03768_),
    .S(_03693_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11722_ (.A1(_03756_),
    .A2(_03763_),
    .A3(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11723_ (.A1(_03751_),
    .A2(_03698_),
    .B(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11724_ (.A1(_03725_),
    .A2(_03771_),
    .ZN(_05892_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11725_ (.I(_05892_),
    .ZN(_05907_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11726_ (.I(\samples_real[0][10] ),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11727_ (.A1(\samples_real[7][10] ),
    .A2(_03753_),
    .B1(_03755_),
    .B2(\samples_real[1][10] ),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11728_ (.A1(\samples_real[4][10] ),
    .A2(_03760_),
    .B1(_03762_),
    .B2(\samples_real[2][10] ),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11729_ (.A1(\samples_real[6][10] ),
    .A2(_03758_),
    .B1(_03764_),
    .B2(\samples_real[3][10] ),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11730_ (.A1(\samples_real[5][10] ),
    .A2(_03767_),
    .B(_03696_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11731_ (.I0(_03775_),
    .I1(_03776_),
    .S(_03693_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11732_ (.A1(_03773_),
    .A2(_03774_),
    .A3(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11733_ (.A1(_03772_),
    .A2(_03698_),
    .B(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11734_ (.A1(_00010_),
    .A2(_03779_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11735_ (.I(_05964_),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11736_ (.I(\samples_imag[0][8] ),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11737_ (.I0(\samples_imag[4][8] ),
    .I1(\samples_imag[5][8] ),
    .S(_03674_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11738_ (.A1(_03675_),
    .A2(\samples_imag[7][8] ),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11739_ (.I0(_03781_),
    .I1(_03782_),
    .S(_03671_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11740_ (.A1(\samples_imag[6][8] ),
    .A2(_03758_),
    .B1(_03764_),
    .B2(\samples_imag[3][8] ),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11741_ (.A1(_03683_),
    .A2(\samples_imag[2][8] ),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11742_ (.A1(_03684_),
    .A2(\samples_imag[1][8] ),
    .B1(_03785_),
    .B2(_03692_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11743_ (.A1(_03692_),
    .A2(_03784_),
    .B1(_03786_),
    .B2(_03679_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11744_ (.A1(_03680_),
    .A2(_03783_),
    .B(_03787_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11745_ (.A1(_03780_),
    .A2(_03697_),
    .B(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11746_ (.A1(_03726_),
    .A2(_03789_),
    .Z(_05908_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11747_ (.I(\samples_imag[0][7] ),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11748_ (.I0(\samples_imag[2][7] ),
    .I1(\samples_imag[3][7] ),
    .I2(\samples_imag[6][7] ),
    .I3(\samples_imag[7][7] ),
    .S0(_03675_),
    .S1(_03680_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11749_ (.A1(_03672_),
    .A2(_03791_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11750_ (.I0(\samples_imag[1][7] ),
    .I1(\samples_imag[5][7] ),
    .S(_03679_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11751_ (.A1(_03676_),
    .A2(_03688_),
    .A3(\samples_imag[4][7] ),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11752_ (.A1(_03684_),
    .A2(_03793_),
    .B(_03794_),
    .C(_03693_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11753_ (.A1(_03790_),
    .A2(_03698_),
    .B1(_03792_),
    .B2(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11754_ (.A1(_00008_),
    .A2(_03796_),
    .Z(_05950_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11755_ (.I(\samples_imag[0][6] ),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11756_ (.A1(_03735_),
    .A2(\samples_imag[1][6] ),
    .B1(_03767_),
    .B2(\samples_imag[5][6] ),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11757_ (.A1(_03673_),
    .A2(_03798_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11758_ (.A1(_03691_),
    .A2(_03687_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11759_ (.A1(\samples_imag[6][6] ),
    .A2(_03707_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11760_ (.A1(_03800_),
    .A2(_03801_),
    .B(_03685_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11761_ (.A1(\samples_imag[4][6] ),
    .A2(_03760_),
    .B1(_03762_),
    .B2(\samples_imag[2][6] ),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11762_ (.A1(\idx2[1] ),
    .A2(_03674_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11763_ (.A1(_03677_),
    .A2(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11764_ (.I(_03805_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11765_ (.A1(\samples_imag[7][6] ),
    .A2(_03753_),
    .B1(_03806_),
    .B2(\samples_imag[3][6] ),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11766_ (.A1(_03799_),
    .A2(_03802_),
    .A3(_03803_),
    .A4(_03807_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11767_ (.A1(_03797_),
    .A2(_03728_),
    .B(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11768_ (.A1(_03740_),
    .A2(_03809_),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11769_ (.I(_06040_),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11770_ (.A1(_03688_),
    .A2(\samples_imag[2][4] ),
    .B1(_03707_),
    .B2(\samples_imag[6][4] ),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11771_ (.A1(\samples_imag[5][4] ),
    .A2(_03766_),
    .B(_03696_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11772_ (.A1(\samples_imag[4][4] ),
    .A2(_03759_),
    .B1(_03806_),
    .B2(\samples_imag[3][4] ),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11773_ (.A1(\samples_imag[7][4] ),
    .A2(_03752_),
    .B1(_03755_),
    .B2(\samples_imag[1][4] ),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11774_ (.A1(_03812_),
    .A2(_03813_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11775_ (.A1(_03676_),
    .A2(_03810_),
    .B1(_03811_),
    .B2(_03671_),
    .C(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11776_ (.A1(\samples_imag[0][4] ),
    .A2(_03711_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11777_ (.A1(_03815_),
    .A2(_03816_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11778_ (.A1(_03726_),
    .A2(_03817_),
    .Z(_06145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11779_ (.I(\samples_real[0][9] ),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11780_ (.A1(\samples_real[7][9] ),
    .A2(_03753_),
    .B1(_03806_),
    .B2(\samples_real[3][9] ),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11781_ (.A1(_03692_),
    .A2(_03767_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11782_ (.I(\samples_real[4][9] ),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11783_ (.I(\samples_real[6][9] ),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11784_ (.I(\samples_real[2][9] ),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11785_ (.I0(_03822_),
    .I1(_03823_),
    .S(_03717_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _11786_ (.A1(_03821_),
    .A2(_03703_),
    .B1(_03824_),
    .B2(_03671_),
    .C(_03676_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11787_ (.A1(\samples_real[1][9] ),
    .A2(_03755_),
    .B1(_03820_),
    .B2(\samples_real[5][9] ),
    .C(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11788_ (.A1(_03818_),
    .A2(_03698_),
    .B1(_03819_),
    .B2(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11789_ (.A1(_03715_),
    .A2(_03827_),
    .Z(_05927_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11790_ (.I(_05927_),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11791_ (.A1(_03688_),
    .A2(\samples_imag[1][5] ),
    .B1(_03767_),
    .B2(\samples_imag[5][5] ),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11792_ (.A1(\samples_imag[6][5] ),
    .A2(_03707_),
    .B(_03800_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11793_ (.A1(\samples_imag[4][5] ),
    .A2(_03759_),
    .B1(_03762_),
    .B2(\samples_imag[2][5] ),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11794_ (.A1(\samples_imag[7][5] ),
    .A2(_03752_),
    .B1(_03806_),
    .B2(\samples_imag[3][5] ),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11795_ (.A1(_03830_),
    .A2(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11796_ (.A1(_03672_),
    .A2(_03828_),
    .B1(_03829_),
    .B2(_03676_),
    .C(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11797_ (.A1(\samples_imag[0][5] ),
    .A2(_03712_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11798_ (.A1(_03833_),
    .A2(_03834_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11799_ (.A1(_03725_),
    .A2(_03835_),
    .Z(_06094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11800_ (.I(\samples_imag[0][3] ),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11801_ (.I0(\samples_imag[1][3] ),
    .I1(\samples_imag[5][3] ),
    .S(_03678_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11802_ (.A1(_03717_),
    .A2(\samples_imag[4][3] ),
    .B(_03691_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11803_ (.A1(_03717_),
    .A2(\samples_imag[2][3] ),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11804_ (.A1(_03838_),
    .A2(_03839_),
    .B(_03675_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11805_ (.I0(\samples_imag[3][3] ),
    .I1(\samples_imag[7][3] ),
    .S(_03677_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11806_ (.A1(\samples_imag[6][3] ),
    .A2(_03758_),
    .B1(_03841_),
    .B2(_03674_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11807_ (.A1(_03692_),
    .A2(_03842_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11808_ (.A1(_03754_),
    .A2(_03837_),
    .B(_03840_),
    .C(_03843_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11809_ (.A1(_03836_),
    .A2(_03697_),
    .B(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11810_ (.A1(_03740_),
    .A2(_03845_),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11811_ (.I(_06255_),
    .ZN(_06205_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11812_ (.I(\samples_imag[0][2] ),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11813_ (.A1(_03717_),
    .A2(\samples_imag[2][2] ),
    .B1(_03706_),
    .B2(\samples_imag[6][2] ),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11814_ (.A1(_03675_),
    .A2(_03847_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11815_ (.A1(\samples_imag[5][2] ),
    .A2(_03766_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11816_ (.A1(_03696_),
    .A2(_03849_),
    .B(_03692_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11817_ (.A1(\samples_imag[4][2] ),
    .A2(_03760_),
    .B1(_03806_),
    .B2(\samples_imag[3][2] ),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11818_ (.A1(\samples_imag[7][2] ),
    .A2(_03752_),
    .B1(_03755_),
    .B2(\samples_imag[1][2] ),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11819_ (.A1(_03848_),
    .A2(_03850_),
    .A3(_03851_),
    .A4(_03852_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11820_ (.A1(_03846_),
    .A2(_03697_),
    .B(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11821_ (.A1(_03725_),
    .A2(_03854_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11822_ (.I(_06256_),
    .ZN(_06471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11823_ (.I(\samples_real[0][8] ),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11824_ (.I0(\samples_real[4][8] ),
    .I1(\samples_real[5][8] ),
    .S(_03729_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11825_ (.A1(_03729_),
    .A2(\samples_real[7][8] ),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11826_ (.I0(_03856_),
    .I1(_03857_),
    .S(_03673_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11827_ (.A1(\samples_real[6][8] ),
    .A2(_03758_),
    .B1(_03764_),
    .B2(\samples_real[3][8] ),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11828_ (.I(\samples_real[1][8] ),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11829_ (.A1(_03729_),
    .A2(_03860_),
    .B(_03672_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11830_ (.A1(_03685_),
    .A2(\samples_real[2][8] ),
    .B(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11831_ (.A1(_03693_),
    .A2(_03859_),
    .B1(_03862_),
    .B2(_03680_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11832_ (.A1(_03731_),
    .A2(_03858_),
    .B(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11833_ (.A1(_03855_),
    .A2(_03728_),
    .B(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11834_ (.A1(_03715_),
    .A2(_03865_),
    .Z(_05928_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11835_ (.I(_05928_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11836_ (.I(\samples_imag[0][1] ),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11837_ (.I0(\samples_imag[3][1] ),
    .I1(\samples_imag[7][1] ),
    .S(_03677_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11838_ (.A1(_03678_),
    .A2(\samples_imag[5][1] ),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11839_ (.I0(_03867_),
    .I1(_03868_),
    .S(_03691_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11840_ (.I0(\samples_imag[2][1] ),
    .I1(\samples_imag[6][1] ),
    .S(_03678_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11841_ (.A1(_03717_),
    .A2(\samples_imag[4][1] ),
    .B(_03683_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11842_ (.A1(_03717_),
    .A2(\samples_imag[1][1] ),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11843_ (.A1(_03871_),
    .A2(_03872_),
    .B(_03671_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11844_ (.A1(_03675_),
    .A2(_03869_),
    .B1(_03870_),
    .B2(_03745_),
    .C(_03873_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11845_ (.A1(_03866_),
    .A2(_03697_),
    .B(_03874_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11846_ (.A1(_03740_),
    .A2(_03875_),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _11847_ (.I(_06303_),
    .ZN(_07898_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11848_ (.I(_00009_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11849_ (.I(_03876_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11850_ (.I(\samples_real[0][13] ),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11851_ (.I0(\samples_real[1][13] ),
    .I1(\samples_real[5][13] ),
    .S(_03678_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11852_ (.A1(_03717_),
    .A2(\samples_real[4][13] ),
    .B(_03691_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11853_ (.A1(_03717_),
    .A2(\samples_real[2][13] ),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11854_ (.A1(_03880_),
    .A2(_03881_),
    .B(_03675_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11855_ (.I0(\samples_real[3][13] ),
    .I1(\samples_real[7][13] ),
    .S(_03677_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11856_ (.A1(\samples_real[6][13] ),
    .A2(_03758_),
    .B1(_03883_),
    .B2(_03675_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11857_ (.A1(_03692_),
    .A2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11858_ (.A1(_03754_),
    .A2(_03879_),
    .B(_03882_),
    .C(_03885_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11859_ (.A1(_03878_),
    .A2(_03697_),
    .B(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11860_ (.A1(_03877_),
    .A2(_03887_),
    .Z(_05924_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11861_ (.I(\samples_real[0][7] ),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11862_ (.A1(_03688_),
    .A2(\samples_real[2][7] ),
    .B1(_03707_),
    .B2(\samples_real[6][7] ),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11863_ (.A1(_03676_),
    .A2(_03889_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11864_ (.A1(\samples_real[5][7] ),
    .A2(_03767_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11865_ (.A1(_03696_),
    .A2(_03891_),
    .B(_03693_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11866_ (.A1(\samples_real[4][7] ),
    .A2(_03760_),
    .B1(_03806_),
    .B2(\samples_real[3][7] ),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11867_ (.A1(\samples_real[7][7] ),
    .A2(_03753_),
    .B1(_03755_),
    .B2(\samples_real[1][7] ),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11868_ (.A1(_03890_),
    .A2(_03892_),
    .A3(_03893_),
    .A4(_03894_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11869_ (.A1(_03888_),
    .A2(_03698_),
    .B(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11870_ (.A1(_00010_),
    .A2(_03896_),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11871_ (.I(_05969_),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11872_ (.I(_00012_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11873_ (.I(_03897_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11874_ (.A1(_03898_),
    .A2(_03724_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11875_ (.A1(_03735_),
    .A2(\samples_real[1][6] ),
    .B1(_03767_),
    .B2(\samples_real[5][6] ),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11876_ (.A1(\samples_real[6][6] ),
    .A2(_03707_),
    .B(_03800_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11877_ (.A1(\samples_real[4][6] ),
    .A2(_03760_),
    .B1(_03762_),
    .B2(\samples_real[2][6] ),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11878_ (.A1(\samples_real[7][6] ),
    .A2(_03753_),
    .B1(_03806_),
    .B2(\samples_real[3][6] ),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11879_ (.A1(_03901_),
    .A2(_03902_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11880_ (.A1(_03673_),
    .A2(_03899_),
    .B1(_03900_),
    .B2(_03730_),
    .C(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11881_ (.I(_03712_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11882_ (.A1(\samples_real[0][6] ),
    .A2(_03905_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11883_ (.A1(_03904_),
    .A2(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11884_ (.A1(_03715_),
    .A2(_03907_),
    .Z(_05932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11885_ (.I(_05932_),
    .ZN(_06095_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11886_ (.I(\samples_real[0][5] ),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11887_ (.I0(\samples_real[6][5] ),
    .I1(\samples_real[7][5] ),
    .S(_03730_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11888_ (.A1(\samples_real[1][5] ),
    .A2(_03755_),
    .B1(_03909_),
    .B2(_03707_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11889_ (.A1(\samples_real[5][5] ),
    .A2(_03703_),
    .B1(_03704_),
    .B2(\samples_real[3][5] ),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11890_ (.A1(_03735_),
    .A2(\samples_real[4][5] ),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11891_ (.A1(_03735_),
    .A2(\samples_real[2][5] ),
    .B1(_03912_),
    .B2(_03737_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11892_ (.I0(_03911_),
    .I1(_03913_),
    .S(_03685_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11893_ (.A1(_03908_),
    .A2(_03728_),
    .B1(_03910_),
    .B2(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11894_ (.A1(_00011_),
    .A2(_03915_),
    .Z(_05933_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11895_ (.I(\samples_imag[0][0] ),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11896_ (.I0(\samples_imag[3][0] ),
    .I1(\samples_imag[7][0] ),
    .S(_03677_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11897_ (.A1(_03677_),
    .A2(\samples_imag[5][0] ),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11898_ (.I0(_03917_),
    .I1(_03918_),
    .S(_03691_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11899_ (.I0(\samples_imag[2][0] ),
    .I1(\samples_imag[6][0] ),
    .S(_03678_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11900_ (.A1(_03687_),
    .A2(\samples_imag[4][0] ),
    .B(_03683_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11901_ (.A1(_03687_),
    .A2(\samples_imag[1][0] ),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11902_ (.A1(_03921_),
    .A2(_03922_),
    .B(_03671_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11903_ (.A1(_03675_),
    .A2(_03919_),
    .B1(_03920_),
    .B2(_03745_),
    .C(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11904_ (.A1(_03916_),
    .A2(_03697_),
    .B(_03924_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11905_ (.A1(_00008_),
    .A2(_03925_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11906_ (.I(_06337_),
    .ZN(_06341_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11907_ (.A1(_03877_),
    .A2(_03724_),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11908_ (.A1(_03715_),
    .A2(_03915_),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _11909_ (.I(_06065_),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11910_ (.I(\samples_real[0][4] ),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11911_ (.I0(\samples_real[2][4] ),
    .I1(\samples_real[3][4] ),
    .I2(\samples_real[6][4] ),
    .I3(\samples_real[7][4] ),
    .S0(_03730_),
    .S1(_03731_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11912_ (.A1(_03673_),
    .A2(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11913_ (.I0(\samples_real[1][4] ),
    .I1(\samples_real[5][4] ),
    .S(_03731_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11914_ (.A1(_03730_),
    .A2(_03735_),
    .A3(\samples_real[4][4] ),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11915_ (.A1(_03685_),
    .A2(_03929_),
    .B(_03930_),
    .C(_03737_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11916_ (.A1(_03926_),
    .A2(_03728_),
    .B1(_03928_),
    .B2(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11917_ (.A1(_03715_),
    .A2(_03932_),
    .Z(_06011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11918_ (.I(_06011_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _11919_ (.I(_00011_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11920_ (.I(\samples_real[0][3] ),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11921_ (.A1(\samples_real[7][3] ),
    .A2(_03753_),
    .B1(_03755_),
    .B2(\samples_real[1][3] ),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11922_ (.A1(\samples_real[4][3] ),
    .A2(_03760_),
    .B1(_03762_),
    .B2(\samples_real[2][3] ),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11923_ (.A1(\samples_real[6][3] ),
    .A2(_03758_),
    .B1(_03764_),
    .B2(\samples_real[3][3] ),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11924_ (.A1(\samples_real[5][3] ),
    .A2(_03767_),
    .B(_03696_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11925_ (.I0(_03937_),
    .I1(_03938_),
    .S(_03737_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11926_ (.A1(_03935_),
    .A2(_03936_),
    .A3(_03939_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11927_ (.A1(_03934_),
    .A2(_03728_),
    .B(_03940_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11928_ (.A1(_03933_),
    .A2(_03941_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11929_ (.I(_05988_),
    .ZN(_06001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11930_ (.A1(_03688_),
    .A2(\samples_real[1][2] ),
    .B1(_03766_),
    .B2(\samples_real[5][2] ),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11931_ (.A1(\samples_real[6][2] ),
    .A2(_03706_),
    .B(_03800_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11932_ (.A1(\samples_real[4][2] ),
    .A2(_03759_),
    .B1(_03762_),
    .B2(\samples_real[2][2] ),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11933_ (.A1(\samples_real[7][2] ),
    .A2(_03752_),
    .B1(_03805_),
    .B2(\samples_real[3][2] ),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11934_ (.A1(_03944_),
    .A2(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11935_ (.A1(_03672_),
    .A2(_03942_),
    .B1(_03943_),
    .B2(_03676_),
    .C(_03946_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11936_ (.A1(\samples_real[0][2] ),
    .A2(_03711_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11937_ (.A1(_03947_),
    .A2(_03948_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11938_ (.A1(_03933_),
    .A2(_03949_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11939_ (.I(_05989_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _11940_ (.I(_00010_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11941_ (.A1(_03950_),
    .A2(_03941_),
    .ZN(_05997_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11942_ (.I(_05997_),
    .ZN(_06169_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11943_ (.A1(_03735_),
    .A2(\samples_real[4][1] ),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11944_ (.A1(_03735_),
    .A2(\samples_real[2][1] ),
    .B1(_03951_),
    .B2(_03737_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11945_ (.I0(\samples_real[3][1] ),
    .I1(\samples_real[7][1] ),
    .S(_03731_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11946_ (.A1(\samples_real[6][1] ),
    .A2(_03758_),
    .B1(_03953_),
    .B2(_03730_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11947_ (.I0(\samples_real[1][1] ),
    .I1(\samples_real[5][1] ),
    .S(_03731_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11948_ (.A1(_03754_),
    .A2(_03955_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11949_ (.A1(_03730_),
    .A2(_03952_),
    .B1(_03954_),
    .B2(_03737_),
    .C(_03956_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11950_ (.A1(\samples_real[0][1] ),
    .A2(_03905_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11951_ (.A1(_03957_),
    .A2(_03958_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11952_ (.A1(_03933_),
    .A2(_03959_),
    .ZN(_05998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11953_ (.I(_05998_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11954_ (.A1(_03950_),
    .A2(_03949_),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _11955_ (.I(_06016_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11956_ (.I(\samples_real[0][0] ),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11957_ (.I0(\samples_real[3][0] ),
    .I1(\samples_real[7][0] ),
    .S(_03678_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11958_ (.A1(_03679_),
    .A2(\samples_real[5][0] ),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11959_ (.I0(_03961_),
    .I1(_03962_),
    .S(_03692_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11960_ (.I0(\samples_real[2][0] ),
    .I1(\samples_real[6][0] ),
    .S(_03679_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11961_ (.A1(_03688_),
    .A2(\samples_real[4][0] ),
    .B(_03684_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11962_ (.A1(_03688_),
    .A2(\samples_real[1][0] ),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11963_ (.A1(_03965_),
    .A2(_03966_),
    .B(_03671_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11964_ (.A1(_03729_),
    .A2(_03963_),
    .B1(_03964_),
    .B2(_03745_),
    .C(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11965_ (.A1(_03960_),
    .A2(_03698_),
    .B(_03968_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11966_ (.A1(_03933_),
    .A2(_03969_),
    .ZN(_06017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11967_ (.I(_06017_),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11968_ (.A1(_03950_),
    .A2(_03959_),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11969_ (.I(_06404_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11970_ (.I(\samples_imag[0][13] ),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11971_ (.I0(\samples_imag[3][13] ),
    .I1(\samples_imag[7][13] ),
    .S(_03679_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11972_ (.A1(_03679_),
    .A2(\samples_imag[5][13] ),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11973_ (.I0(_03971_),
    .I1(_03972_),
    .S(_03693_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11974_ (.I0(\samples_imag[2][13] ),
    .I1(\samples_imag[6][13] ),
    .S(_03680_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11975_ (.A1(_03689_),
    .A2(\samples_imag[4][13] ),
    .B(_03684_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11976_ (.A1(_03689_),
    .A2(\samples_imag[1][13] ),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11977_ (.A1(_03975_),
    .A2(_03976_),
    .B(_03672_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11978_ (.A1(_03729_),
    .A2(_03973_),
    .B1(_03974_),
    .B2(_03745_),
    .C(_03977_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11979_ (.A1(_03970_),
    .A2(_03698_),
    .B(_03978_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11980_ (.A1(_03725_),
    .A2(_03979_),
    .Z(_07909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11981_ (.A1(_03950_),
    .A2(_03969_),
    .ZN(_06435_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _11982_ (.I(_06435_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11983_ (.A1(_03877_),
    .A2(_03779_),
    .Z(_06104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11984_ (.A1(_03898_),
    .A2(_03865_),
    .ZN(_06153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11985_ (.A1(_03877_),
    .A2(_03865_),
    .Z(_06214_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _11986_ (.I(_03876_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11987_ (.A1(_03980_),
    .A2(_03896_),
    .Z(_06264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11988_ (.A1(_03980_),
    .A2(_03907_),
    .Z(_06311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11989_ (.A1(_03898_),
    .A2(_03932_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11990_ (.A1(_03898_),
    .A2(_03949_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11991_ (.A1(_03980_),
    .A2(_03932_),
    .Z(_08021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11992_ (.A1(_03898_),
    .A2(_03959_),
    .ZN(_06436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11993_ (.A1(_03980_),
    .A2(_03959_),
    .Z(_08052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11994_ (.A1(_03898_),
    .A2(_03969_),
    .Z(_08053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11995_ (.A1(_08039_),
    .A2(_07926_),
    .Z(_06441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11996_ (.A1(_00009_),
    .A2(_03969_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11997_ (.I(_03981_),
    .ZN(_08090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11998_ (.I(_08078_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11999_ (.A1(_06301_),
    .A2(_08082_),
    .Z(_06488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12000_ (.A1(_03933_),
    .A2(_03925_),
    .ZN(_06856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12001_ (.I(_06856_),
    .ZN(_08101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12002_ (.A1(_03726_),
    .A2(_03887_),
    .Z(_08102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12003_ (.A1(_00011_),
    .A2(_03875_),
    .Z(_06501_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12004_ (.I(_06501_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12005_ (.A1(_00010_),
    .A2(_03854_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12006_ (.I(_06567_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12007_ (.A1(_03715_),
    .A2(_03875_),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12008_ (.I(_06496_),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12009_ (.A1(_03933_),
    .A2(_03854_),
    .ZN(_06632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12010_ (.I(_06632_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12011_ (.A1(_00011_),
    .A2(_03845_),
    .ZN(_06568_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12012_ (.I(_06568_),
    .ZN(_06498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12013_ (.A1(_03933_),
    .A2(_03817_),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12014_ (.A1(_00010_),
    .A2(_03835_),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12015_ (.I(_06534_),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12016_ (.A1(_00010_),
    .A2(_03817_),
    .Z(_06505_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12017_ (.I(_06505_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12018_ (.A1(_00011_),
    .A2(_03835_),
    .Z(_06506_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12019_ (.I(_06506_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12020_ (.A1(_03950_),
    .A2(_03809_),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12021_ (.I(_06578_),
    .ZN(_06507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12022_ (.A1(_03740_),
    .A2(_03700_),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12023_ (.I(_06613_),
    .ZN(_06616_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12024_ (.A1(_00011_),
    .A2(_03809_),
    .Z(_08107_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12025_ (.I(_08107_),
    .ZN(_06546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12026_ (.A1(_03950_),
    .A2(_03796_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12027_ (.I(_06547_),
    .ZN(_06691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12028_ (.A1(_03933_),
    .A2(_03796_),
    .ZN(_06520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12029_ (.A1(_03950_),
    .A2(_03789_),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12030_ (.I(_06521_),
    .ZN(_06692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12031_ (.A1(_03950_),
    .A2(_03771_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12032_ (.I(_06522_),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12033_ (.A1(_03950_),
    .A2(_03750_),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12034_ (.I(_06580_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12035_ (.A1(_03715_),
    .A2(_03739_),
    .Z(_06517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12036_ (.A1(_03715_),
    .A2(_03714_),
    .Z(_06525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12037_ (.A1(_03740_),
    .A2(_03724_),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12038_ (.I(_06600_),
    .ZN(_06663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12039_ (.A1(_03898_),
    .A2(_03979_),
    .Z(_08111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12040_ (.A1(_03689_),
    .A2(\samples_imag[1][14] ),
    .B1(_03767_),
    .B2(\samples_imag[5][14] ),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12041_ (.A1(\samples_imag[6][14] ),
    .A2(_03707_),
    .B(_03800_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12042_ (.A1(\samples_imag[4][14] ),
    .A2(_03760_),
    .B1(_03762_),
    .B2(\samples_imag[2][14] ),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12043_ (.A1(\samples_imag[7][14] ),
    .A2(_03753_),
    .B1(_03806_),
    .B2(\samples_imag[3][14] ),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12044_ (.A1(_03984_),
    .A2(_03985_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12045_ (.A1(_03672_),
    .A2(_03982_),
    .B1(_03983_),
    .B2(_03729_),
    .C(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12046_ (.A1(\samples_imag[0][14] ),
    .A2(_03712_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12047_ (.A1(_03987_),
    .A2(_03988_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12048_ (.A1(_03980_),
    .A2(_03989_),
    .Z(_08112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12049_ (.A1(_00008_),
    .A2(_03949_),
    .ZN(_06918_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12050_ (.I(_06918_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12051_ (.A1(_03726_),
    .A2(_03959_),
    .Z(_06748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12052_ (.A1(_03726_),
    .A2(_03932_),
    .Z(_08116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12053_ (.I(_08116_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12054_ (.A1(_03726_),
    .A2(_03779_),
    .Z(_06601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12055_ (.A1(_03725_),
    .A2(_03969_),
    .Z(_06803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12056_ (.A1(_03740_),
    .A2(_03941_),
    .ZN(_06873_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12057_ (.I(_06873_),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12058_ (.A1(_03740_),
    .A2(_03915_),
    .ZN(_06767_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12059_ (.I(_06767_),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12060_ (.A1(_03725_),
    .A2(_03896_),
    .Z(_08126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12061_ (.I(_08126_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12062_ (.A1(_03740_),
    .A2(_03865_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12063_ (.I(_06668_),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12064_ (.A1(_03726_),
    .A2(_03907_),
    .ZN(_06719_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12065_ (.I(_06719_),
    .ZN(_06913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12066_ (.A1(_03726_),
    .A2(_03827_),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12067_ (.I(_06605_),
    .ZN(_06602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12068_ (.A1(_08305_),
    .A2(_06803_),
    .Z(_08306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12069_ (.I(_07789_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12070_ (.A1(_03594_),
    .A2(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12071_ (.I(_03991_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12072_ (.A1(_03933_),
    .A2(_03907_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12073_ (.A1(_03933_),
    .A2(_03932_),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12074_ (.I(_07912_),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12075_ (.I(_08125_),
    .ZN(_06606_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12076_ (.I(_06676_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12077_ (.I(_08181_),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12078_ (.I(_08195_),
    .ZN(_06865_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12079_ (.I(_06868_),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12080_ (.I(_06842_),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12081_ (.I(_06849_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12082_ (.I(_06901_),
    .ZN(_06903_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12083_ (.I(_08212_),
    .ZN(_06908_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12084_ (.I(_08226_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12085_ (.I(_08244_),
    .ZN(_06997_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12086_ (.I(_06900_),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12087_ (.I(_08246_),
    .ZN(_07039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12088_ (.A1(_03898_),
    .A2(_03887_),
    .ZN(_05918_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12089_ (.I(_07918_),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12090_ (.I(_07950_),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12091_ (.I(_07961_),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12092_ (.I(_06466_),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12093_ (.I(_06476_),
    .ZN(_06472_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12094_ (.I(_08084_),
    .ZN(_06492_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12095_ (.I(_08122_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12096_ (.I(_08140_),
    .ZN(_06659_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12097_ (.I(_08153_),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12098_ (.I(_08165_),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12099_ (.I(_08178_),
    .ZN(_06816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12100_ (.I(_08183_),
    .ZN(_06847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12101_ (.I(_06874_),
    .ZN(_06914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12102_ (.I(_06934_),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12103_ (.I(_08276_),
    .ZN(_07040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12104_ (.I(_07065_),
    .ZN(_07062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12105_ (.I(_08287_),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12106_ (.I(_07075_),
    .ZN(_07070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12107_ (.I(_07701_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12108_ (.I(_07815_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12109_ (.I(\samples_real[0][14] ),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12110_ (.I0(\samples_real[3][14] ),
    .I1(\samples_real[7][14] ),
    .S(_03679_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12111_ (.A1(_03679_),
    .A2(\samples_real[5][14] ),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12112_ (.I0(_03993_),
    .I1(_03994_),
    .S(_03693_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12113_ (.I0(\samples_real[2][14] ),
    .I1(\samples_real[6][14] ),
    .S(_03680_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12114_ (.A1(_03689_),
    .A2(\samples_real[4][14] ),
    .B(_03684_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12115_ (.A1(_03689_),
    .A2(\samples_real[1][14] ),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12116_ (.A1(_03997_),
    .A2(_03998_),
    .B(_03672_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12117_ (.A1(_03729_),
    .A2(_03995_),
    .B1(_03996_),
    .B2(_03745_),
    .C(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12118_ (.A1(_03992_),
    .A2(_03698_),
    .B(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12119_ (.A1(_03877_),
    .A2(_04001_),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12120_ (.A1(_03877_),
    .A2(_03700_),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12121_ (.A1(_03877_),
    .A2(_03827_),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12122_ (.I(_07949_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12123_ (.I(_07960_),
    .ZN(_06273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12124_ (.A1(_03877_),
    .A2(_03915_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12125_ (.A1(_03877_),
    .A2(_03941_),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12126_ (.A1(_03877_),
    .A2(_03949_),
    .ZN(_06437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12127_ (.I(_06454_),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12128_ (.I(_06477_),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12129_ (.I(_08133_),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12130_ (.I(_08121_),
    .ZN(_06629_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12131_ (.I(_08139_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12132_ (.I(_08152_),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12133_ (.I(_08164_),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12134_ (.I(_08186_),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12135_ (.I(_08177_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12136_ (.I(_08182_),
    .ZN(_06848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12137_ (.I(_08201_),
    .ZN(_06867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12138_ (.I(_06869_),
    .ZN(_06894_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12139_ (.I(_08217_),
    .ZN(_06910_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12140_ (.I(_06919_),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12141_ (.A1(_03950_),
    .A2(_03845_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12142_ (.I(_08231_),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12143_ (.I(_08251_),
    .ZN(_06999_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12144_ (.I(_08257_),
    .ZN(_07019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12145_ (.I(_08286_),
    .ZN(_07068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12146_ (.I(_05926_),
    .ZN(_07906_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12147_ (.I(_05938_),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12148_ (.I(_05963_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12149_ (.I(_06019_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12150_ (.I(_06053_),
    .ZN(_07933_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12151_ (.I(_06057_),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12152_ (.I(_06106_),
    .ZN(_07942_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12153_ (.I(_06109_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12154_ (.I(_06160_),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12155_ (.I(_06164_),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12156_ (.I(_06167_),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12157_ (.I(_06216_),
    .ZN(_07965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12158_ (.I(_06220_),
    .ZN(_06260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12159_ (.I(_06250_),
    .ZN(_07974_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12160_ (.I(_06266_),
    .ZN(_07976_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12161_ (.I(_06270_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12162_ (.I(_06298_),
    .ZN(_07984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12163_ (.I(_06302_),
    .ZN(_07986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12164_ (.I(_06313_),
    .ZN(_07989_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12165_ (.I(_06317_),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12166_ (.I(_06340_),
    .ZN(_08018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12167_ (.I(_06378_),
    .ZN(_08007_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12168_ (.I(_06401_),
    .ZN(_08022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12169_ (.I(_06425_),
    .ZN(_08042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12170_ (.I(_06432_),
    .ZN(_08033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12171_ (.I(_06500_),
    .ZN(_08105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12172_ (.I(_06509_),
    .ZN(_06511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12173_ (.I(_06532_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12174_ (.I(_06545_),
    .ZN(_06551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12175_ (.I(_06566_),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12176_ (.I(_06586_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12177_ (.I(_06590_),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12178_ (.I(_06604_),
    .ZN(_06611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12179_ (.I(_06649_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12180_ (.I(_06682_),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12181_ (.I(_06702_),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12182_ (.I(_06739_),
    .ZN(_06785_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12183_ (.I(_06758_),
    .ZN(_06787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12184_ (.I(_06793_),
    .ZN(_06843_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12185_ (.I(_06805_),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12186_ (.I(_06830_),
    .ZN(_06841_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12187_ (.I(_06879_),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12188_ (.I(_06896_),
    .ZN(_06935_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12189_ (.I(_06925_),
    .ZN(_06937_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12190_ (.I(_06943_),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12191_ (.I(_06962_),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12192_ (.I(_06967_),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12193_ (.I(_07038_),
    .ZN(_07041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12194_ (.I(_05925_),
    .ZN(_07901_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12195_ (.I(_05999_),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12196_ (.I(_05981_),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12197_ (.I(_06018_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12198_ (.I(_06052_),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12199_ (.I(_06105_),
    .ZN(_07934_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12200_ (.I(_06215_),
    .ZN(_07954_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12201_ (.I(_06265_),
    .ZN(_07966_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12202_ (.I(_06297_),
    .ZN(_07975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12203_ (.I(_06312_),
    .ZN(_07977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12204_ (.I(_06339_),
    .ZN(_07987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12205_ (.I(_06377_),
    .ZN(_07992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12206_ (.I(_06400_),
    .ZN(_08008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12207_ (.I(_06424_),
    .ZN(_08019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12208_ (.I(_06431_),
    .ZN(_08023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12209_ (.I(_06503_),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12210_ (.I(_06540_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12211_ (.I(_06565_),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12212_ (.I(_06574_),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12213_ (.I(_06585_),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12214_ (.I(_06617_),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12215_ (.I(_06644_),
    .ZN(_06654_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12216_ (.I(_06648_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12217_ (.I(_06681_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12218_ (.I(_06697_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12219_ (.I(_06701_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12220_ (.I(_06738_),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12221_ (.I(_06750_),
    .ZN(_06708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12222_ (.I(_06757_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12223_ (.I(_06792_),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12224_ (.I(_06895_),
    .ZN(_06889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12225_ (.I(_06942_),
    .ZN(_06936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12226_ (.I(_06984_),
    .ZN(_06978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12227_ (.I(_06995_),
    .ZN(_06992_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _12228_ (.I(_07680_),
    .ZN(_07082_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12229_ (.I0(\samples_real[4][14] ),
    .I1(\samples_real[5][14] ),
    .I2(\samples_real[6][14] ),
    .I3(\samples_real[7][14] ),
    .S0(_03609_),
    .S1(_03611_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12230_ (.I(\samples_real[1][14] ),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12231_ (.I0(\samples_real[2][14] ),
    .I1(\samples_real[3][14] ),
    .S(_03609_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12232_ (.I(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12233_ (.A1(_04003_),
    .A2(_03626_),
    .B1(_04005_),
    .B2(_03622_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12234_ (.I0(_04002_),
    .I1(_04006_),
    .S(_03617_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12235_ (.A1(_03601_),
    .A2(_03619_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12236_ (.A1(_03992_),
    .A2(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12237_ (.A1(_04007_),
    .A2(_04009_),
    .Z(_07691_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12238_ (.I(_04008_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12239_ (.A1(\idx1[2] ),
    .A2(_03611_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12240_ (.A1(_03613_),
    .A2(_04011_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12241_ (.I(_04012_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12242_ (.A1(_03601_),
    .A2(\idx1[1] ),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12243_ (.I(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12244_ (.A1(_03613_),
    .A2(_04015_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12245_ (.I(_04016_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12246_ (.A1(\samples_real[7][13] ),
    .A2(_04013_),
    .B1(_04017_),
    .B2(\samples_real[3][13] ),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12247_ (.A1(\idx1[2] ),
    .A2(_03626_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12248_ (.I(_04019_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12249_ (.A1(_03601_),
    .A2(_03626_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12250_ (.I(_04021_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12251_ (.A1(\samples_real[5][13] ),
    .A2(_04020_),
    .B1(_04022_),
    .B2(\samples_real[1][13] ),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12252_ (.I0(\samples_real[4][13] ),
    .I1(\samples_real[6][13] ),
    .S(_03622_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12253_ (.A1(\idx1[2] ),
    .A2(_03599_),
    .A3(\samples_real[2][13] ),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12254_ (.A1(_03617_),
    .A2(_04024_),
    .B(_04025_),
    .C(_03664_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12255_ (.A1(_04018_),
    .A2(_04023_),
    .A3(_04026_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12256_ (.A1(_03878_),
    .A2(_04010_),
    .B(_04027_),
    .ZN(_07696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12257_ (.A1(\samples_real[3][15] ),
    .A2(_03603_),
    .B1(_03605_),
    .B2(\samples_real[6][15] ),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12258_ (.A1(_03599_),
    .A2(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12259_ (.I0(\samples_real[4][15] ),
    .I1(\samples_real[5][15] ),
    .S(_03602_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12260_ (.A1(_03602_),
    .A2(\samples_real[7][15] ),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12261_ (.I0(_04030_),
    .I1(_04031_),
    .S(\idx1[1] ),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12262_ (.I(\samples_real[1][15] ),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12263_ (.A1(_03604_),
    .A2(\samples_real[2][15] ),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12264_ (.A1(_03602_),
    .A2(_04033_),
    .B1(_04034_),
    .B2(\idx1[1] ),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12265_ (.I0(_04032_),
    .I1(_04035_),
    .S(_03601_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12266_ (.A1(\samples_real[0][15] ),
    .A2(_03620_),
    .B1(_04029_),
    .B2(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12267_ (.I(_04037_),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12268_ (.I(_04010_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12269_ (.A1(_03604_),
    .A2(_04011_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12270_ (.I(_04039_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12271_ (.I(_04040_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12272_ (.I0(\samples_real[4][12] ),
    .I1(\samples_real[5][12] ),
    .S(_03643_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12273_ (.A1(_03643_),
    .A2(\samples_real[7][12] ),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12274_ (.A1(_03665_),
    .A2(\samples_real[1][12] ),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12275_ (.I0(\samples_real[2][12] ),
    .I1(\samples_real[3][12] ),
    .S(_03650_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12276_ (.I0(_04042_),
    .I1(_04043_),
    .I2(_04044_),
    .I3(_04045_),
    .S0(_03645_),
    .S1(_03655_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12277_ (.A1(\samples_real[6][12] ),
    .A2(_04041_),
    .B(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12278_ (.A1(_03699_),
    .A2(_04038_),
    .B(_04047_),
    .ZN(_07710_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12279_ (.I0(\samples_real[4][11] ),
    .I1(\samples_real[5][11] ),
    .I2(\samples_real[6][11] ),
    .I3(\samples_real[7][11] ),
    .S0(_03609_),
    .S1(_03611_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12280_ (.I(\samples_real[1][11] ),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12281_ (.I0(\samples_real[2][11] ),
    .I1(\samples_real[3][11] ),
    .S(_03609_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12282_ (.I(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12283_ (.A1(_04049_),
    .A2(_03626_),
    .B1(_04051_),
    .B2(_03611_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12284_ (.I0(_04048_),
    .I1(_04052_),
    .S(_03617_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12285_ (.A1(\samples_real[0][11] ),
    .A2(_03620_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12286_ (.A1(_04053_),
    .A2(_04054_),
    .Z(_07715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12287_ (.I0(\samples_real[5][10] ),
    .I1(\samples_real[7][10] ),
    .S(_03611_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12288_ (.A1(_03622_),
    .A2(\samples_real[3][10] ),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12289_ (.I0(_04055_),
    .I1(_04056_),
    .S(_03617_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12290_ (.I(\idx1[2] ),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12291_ (.I0(\samples_real[2][10] ),
    .I1(\samples_real[6][10] ),
    .S(_04058_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12292_ (.A1(_03611_),
    .A2(_03604_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12293_ (.A1(_03664_),
    .A2(\samples_real[1][10] ),
    .B(_03617_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12294_ (.A1(_03664_),
    .A2(\samples_real[4][10] ),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12295_ (.A1(_04061_),
    .A2(_04062_),
    .B(_03644_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12296_ (.A1(_03643_),
    .A2(_04057_),
    .B1(_04059_),
    .B2(_04060_),
    .C(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12297_ (.A1(_03772_),
    .A2(_04010_),
    .B(_04064_),
    .ZN(_07720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12298_ (.A1(\samples_real[7][9] ),
    .A2(_04013_),
    .B1(_04022_),
    .B2(\samples_real[1][9] ),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12299_ (.I0(_03822_),
    .I1(_03821_),
    .S(_03599_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12300_ (.A1(_03823_),
    .A2(_04015_),
    .B1(_04066_),
    .B2(_04058_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _12301_ (.A1(\samples_real[3][9] ),
    .A2(_04017_),
    .B1(_04020_),
    .B2(\samples_real[5][9] ),
    .C1(_03664_),
    .C2(_04067_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12302_ (.A1(_03818_),
    .A2(_04010_),
    .B1(_04065_),
    .B2(_04068_),
    .ZN(_07725_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12303_ (.I0(\samples_real[4][8] ),
    .I1(\samples_real[5][8] ),
    .I2(\samples_real[6][8] ),
    .I3(\samples_real[7][8] ),
    .S0(_03649_),
    .S1(_03622_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12304_ (.I0(\samples_real[2][8] ),
    .I1(\samples_real[3][8] ),
    .S(_03613_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12305_ (.I(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12306_ (.A1(_03860_),
    .A2(_03626_),
    .B1(_04071_),
    .B2(_03644_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12307_ (.I0(_04069_),
    .I1(_04072_),
    .S(_03654_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12308_ (.A1(_03855_),
    .A2(_04010_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12309_ (.A1(_04073_),
    .A2(_04074_),
    .Z(_07730_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12310_ (.A1(_03604_),
    .A2(_04015_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12311_ (.I(_04075_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12312_ (.A1(\samples_real[7][7] ),
    .A2(_04013_),
    .B1(_04076_),
    .B2(\samples_real[2][7] ),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12313_ (.A1(\idx1[2] ),
    .A2(_03619_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12314_ (.I(_04078_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12315_ (.A1(\samples_real[1][7] ),
    .A2(_04021_),
    .B1(_04079_),
    .B2(\samples_real[4][7] ),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12316_ (.A1(_03622_),
    .A2(_03649_),
    .A3(\samples_real[3][7] ),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12317_ (.A1(\samples_real[5][7] ),
    .A2(_03626_),
    .B1(_04060_),
    .B2(\samples_real[6][7] ),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12318_ (.A1(_04058_),
    .A2(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12319_ (.A1(_04058_),
    .A2(_03619_),
    .A3(_04081_),
    .B(_04083_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12320_ (.A1(_04077_),
    .A2(_04080_),
    .A3(_04084_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12321_ (.A1(_03888_),
    .A2(_04010_),
    .B(_04085_),
    .ZN(_07735_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12322_ (.A1(\samples_real[0][6] ),
    .A2(_03641_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12323_ (.A1(_03664_),
    .A2(\samples_real[1][6] ),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12324_ (.A1(_03665_),
    .A2(\samples_real[4][6] ),
    .B1(_04087_),
    .B2(_03654_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12325_ (.I0(\samples_real[6][6] ),
    .I1(\samples_real[7][6] ),
    .S(_03649_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12326_ (.A1(\samples_real[5][6] ),
    .A2(_03648_),
    .B1(_04089_),
    .B2(_03661_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12327_ (.I0(\samples_real[2][6] ),
    .I1(\samples_real[3][6] ),
    .S(_03649_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12328_ (.A1(_04015_),
    .A2(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12329_ (.A1(_03661_),
    .A2(_04088_),
    .B1(_04090_),
    .B2(_03654_),
    .C(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12330_ (.A1(_04086_),
    .A2(_04093_),
    .Z(_07740_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12331_ (.I(_04021_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12332_ (.I0(\samples_real[6][5] ),
    .I1(\samples_real[7][5] ),
    .S(_03642_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12333_ (.A1(\samples_real[1][5] ),
    .A2(_04094_),
    .B1(_04095_),
    .B2(_04011_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12334_ (.A1(\idx1[2] ),
    .A2(_03599_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12335_ (.A1(\samples_real[3][5] ),
    .A2(_04015_),
    .B1(_04097_),
    .B2(\samples_real[5][5] ),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12336_ (.A1(_03599_),
    .A2(\samples_real[2][5] ),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12337_ (.A1(_03600_),
    .A2(\samples_real[4][5] ),
    .B1(_04099_),
    .B2(_03617_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12338_ (.I0(_04098_),
    .I1(_04100_),
    .S(_03664_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12339_ (.A1(_03908_),
    .A2(_04010_),
    .B1(_04096_),
    .B2(_04101_),
    .ZN(_07745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12340_ (.I0(\samples_real[4][4] ),
    .I1(\samples_real[5][4] ),
    .S(_03650_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12341_ (.A1(_03643_),
    .A2(\samples_real[7][4] ),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12342_ (.A1(_03665_),
    .A2(\samples_real[1][4] ),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12343_ (.I0(\samples_real[2][4] ),
    .I1(\samples_real[3][4] ),
    .S(_03650_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12344_ (.I0(_04102_),
    .I1(_04103_),
    .I2(_04104_),
    .I3(_04105_),
    .S0(_03645_),
    .S1(_03655_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12345_ (.A1(\samples_real[6][4] ),
    .A2(_04041_),
    .B(_04106_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12346_ (.A1(_03926_),
    .A2(_04038_),
    .B(_04107_),
    .ZN(_07750_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12347_ (.I0(\samples_real[4][3] ),
    .I1(\samples_real[5][3] ),
    .I2(\samples_real[6][3] ),
    .I3(\samples_real[7][3] ),
    .S0(_03642_),
    .S1(_03661_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12348_ (.I(\samples_real[1][3] ),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12349_ (.I0(\samples_real[2][3] ),
    .I1(\samples_real[3][3] ),
    .S(_03649_),
    .Z(_04110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12350_ (.I(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12351_ (.A1(_04109_),
    .A2(_03648_),
    .B1(_04111_),
    .B2(_03661_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12352_ (.I0(_04108_),
    .I1(_04112_),
    .S(_03655_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12353_ (.A1(_03934_),
    .A2(_04038_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12354_ (.A1(_04113_),
    .A2(_04114_),
    .Z(_07755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12355_ (.A1(\samples_real[3][2] ),
    .A2(_03603_),
    .B1(_03605_),
    .B2(\samples_real[6][2] ),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12356_ (.A1(_03600_),
    .A2(_04115_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12357_ (.I0(\samples_real[4][2] ),
    .I1(\samples_real[5][2] ),
    .S(_03609_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12358_ (.A1(_03613_),
    .A2(\samples_real[7][2] ),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12359_ (.I0(_04117_),
    .I1(_04118_),
    .S(_03622_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12360_ (.I(\samples_real[1][2] ),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12361_ (.A1(_03664_),
    .A2(\samples_real[2][2] ),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12362_ (.A1(_03642_),
    .A2(_04120_),
    .B1(_04121_),
    .B2(_03644_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12363_ (.I0(_04119_),
    .I1(_04122_),
    .S(_03617_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12364_ (.A1(\samples_real[0][2] ),
    .A2(_03641_),
    .B1(_04116_),
    .B2(_04123_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12365_ (.I(_04124_),
    .ZN(_07760_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12366_ (.I(_05853_),
    .ZN(_05857_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12367_ (.I(\sample_count[0] ),
    .ZN(_07797_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12368_ (.I0(\samples_imag[4][14] ),
    .I1(\samples_imag[5][14] ),
    .I2(\samples_imag[6][14] ),
    .I3(\samples_imag[7][14] ),
    .S0(_03650_),
    .S1(_03661_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12369_ (.I(\samples_imag[1][14] ),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12370_ (.I0(\samples_imag[2][14] ),
    .I1(\samples_imag[3][14] ),
    .S(_03649_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12371_ (.I(_04127_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12372_ (.A1(_04126_),
    .A2(_03648_),
    .B1(_04128_),
    .B2(_03645_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12373_ (.I0(_04125_),
    .I1(_04129_),
    .S(_03655_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12374_ (.A1(\samples_imag[0][14] ),
    .A2(_03641_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12375_ (.A1(_04130_),
    .A2(_04131_),
    .Z(_07805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12376_ (.I0(\samples_imag[2][13] ),
    .I1(\samples_imag[3][13] ),
    .S(_03643_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12377_ (.A1(_03665_),
    .A2(\samples_imag[1][13] ),
    .B(_03655_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12378_ (.A1(_03665_),
    .A2(\samples_imag[4][13] ),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12379_ (.A1(_04133_),
    .A2(_04134_),
    .B(_03645_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12380_ (.A1(\samples_imag[5][13] ),
    .A2(_03648_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12381_ (.I0(\samples_imag[6][13] ),
    .I1(\samples_imag[7][13] ),
    .S(_03650_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12382_ (.A1(_03645_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12383_ (.A1(_04136_),
    .A2(_04138_),
    .B(_03655_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12384_ (.A1(_04015_),
    .A2(_04132_),
    .B(_04135_),
    .C(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12385_ (.A1(_03970_),
    .A2(_04038_),
    .B(_04140_),
    .ZN(_07810_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12386_ (.I0(\samples_imag[4][15] ),
    .I1(\samples_imag[5][15] ),
    .I2(\samples_imag[6][15] ),
    .I3(\samples_imag[7][15] ),
    .S0(_03602_),
    .S1(\idx1[1] ),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12387_ (.I(\samples_imag[1][15] ),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12388_ (.I0(\samples_imag[2][15] ),
    .I1(\samples_imag[3][15] ),
    .S(_03602_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12389_ (.I(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12390_ (.A1(_04142_),
    .A2(_03626_),
    .B1(_04144_),
    .B2(\idx1[1] ),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12391_ (.I0(_04141_),
    .I1(_04145_),
    .S(_03601_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12392_ (.A1(\samples_imag[0][15] ),
    .A2(_03620_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12393_ (.A1(_04146_),
    .A2(_04147_),
    .Z(_07820_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12394_ (.I0(\samples_imag[4][12] ),
    .I1(\samples_imag[5][12] ),
    .I2(\samples_imag[6][12] ),
    .I3(\samples_imag[7][12] ),
    .S0(_03650_),
    .S1(_03661_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12395_ (.I(\samples_imag[1][12] ),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12396_ (.I0(\samples_imag[2][12] ),
    .I1(\samples_imag[3][12] ),
    .S(_03649_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12397_ (.I(_04150_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12398_ (.A1(_04149_),
    .A2(_03648_),
    .B1(_04151_),
    .B2(_03645_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12399_ (.I0(_04148_),
    .I1(_04152_),
    .S(_03655_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12400_ (.A1(\samples_imag[0][12] ),
    .A2(_03641_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12401_ (.A1(_04153_),
    .A2(_04154_),
    .Z(_07824_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12402_ (.I(_04079_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12403_ (.A1(\samples_imag[1][11] ),
    .A2(_04094_),
    .B1(_04155_),
    .B2(\samples_imag[4][11] ),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12404_ (.I(_04017_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12405_ (.I(_04020_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12406_ (.A1(\samples_imag[3][11] ),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\samples_imag[5][11] ),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12407_ (.I0(\samples_imag[6][11] ),
    .I1(\samples_imag[7][11] ),
    .S(_03650_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12408_ (.A1(_04011_),
    .A2(_04160_),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12409_ (.A1(_03600_),
    .A2(\samples_imag[2][11] ),
    .B(_03665_),
    .C(_03655_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12410_ (.A1(_04156_),
    .A2(_04159_),
    .A3(_04161_),
    .A4(_04162_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12411_ (.A1(_03727_),
    .A2(_04038_),
    .B(_04163_),
    .ZN(_07829_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12412_ (.I(_04013_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12413_ (.A1(\samples_imag[7][10] ),
    .A2(_04164_),
    .B1(_04094_),
    .B2(\samples_imag[1][10] ),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12414_ (.I(\samples_imag[2][10] ),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12415_ (.I0(\samples_imag[4][10] ),
    .I1(\samples_imag[6][10] ),
    .S(_03644_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12416_ (.A1(_03654_),
    .A2(_04167_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12417_ (.A1(_04166_),
    .A2(_04015_),
    .B(_04168_),
    .C(_03643_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12418_ (.A1(\samples_imag[3][10] ),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\samples_imag[5][10] ),
    .C(_04169_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12419_ (.A1(_03741_),
    .A2(_04038_),
    .B1(_04165_),
    .B2(_04170_),
    .ZN(_07834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12420_ (.I0(\samples_imag[6][9] ),
    .I1(\samples_imag[7][9] ),
    .S(_03642_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12421_ (.A1(\samples_imag[1][9] ),
    .A2(_04094_),
    .B1(_04171_),
    .B2(_04011_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12422_ (.A1(\samples_imag[3][9] ),
    .A2(_04015_),
    .B1(_04097_),
    .B2(\samples_imag[5][9] ),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12423_ (.A1(_03600_),
    .A2(\samples_imag[2][9] ),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12424_ (.A1(_03600_),
    .A2(\samples_imag[4][9] ),
    .B1(_04174_),
    .B2(_03654_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12425_ (.I0(_04173_),
    .I1(_04175_),
    .S(_03665_),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12426_ (.A1(_03751_),
    .A2(_04038_),
    .B1(_04172_),
    .B2(_04176_),
    .ZN(_07839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12427_ (.I0(\samples_imag[6][8] ),
    .I1(\samples_imag[7][8] ),
    .S(_03642_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12428_ (.A1(\samples_imag[1][8] ),
    .A2(_04094_),
    .B1(_04177_),
    .B2(_04011_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12429_ (.A1(\samples_imag[3][8] ),
    .A2(_04015_),
    .B1(_04097_),
    .B2(\samples_imag[5][8] ),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12430_ (.A1(_03599_),
    .A2(\samples_imag[2][8] ),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12431_ (.A1(_03600_),
    .A2(\samples_imag[4][8] ),
    .B1(_04180_),
    .B2(_03654_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12432_ (.I0(_04179_),
    .I1(_04181_),
    .S(_03665_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12433_ (.A1(_03780_),
    .A2(_04038_),
    .B1(_04178_),
    .B2(_04182_),
    .ZN(_07844_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12434_ (.I0(\samples_imag[4][7] ),
    .I1(\samples_imag[5][7] ),
    .I2(\samples_imag[6][7] ),
    .I3(\samples_imag[7][7] ),
    .S0(_03642_),
    .S1(_03661_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12435_ (.I(\samples_imag[1][7] ),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12436_ (.I0(\samples_imag[2][7] ),
    .I1(\samples_imag[3][7] ),
    .S(_03613_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12437_ (.I(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12438_ (.A1(_04184_),
    .A2(_03648_),
    .B1(_04186_),
    .B2(_03661_),
    .C(_04058_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12439_ (.A1(_04058_),
    .A2(_04183_),
    .B(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12440_ (.A1(_03790_),
    .A2(_04038_),
    .B(_04188_),
    .ZN(_07849_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12441_ (.I(_04076_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12442_ (.I0(\samples_imag[5][6] ),
    .I1(\samples_imag[7][6] ),
    .S(_03622_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12443_ (.A1(_04058_),
    .A2(_03650_),
    .A3(_04190_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12444_ (.A1(\samples_imag[2][6] ),
    .A2(_04189_),
    .B(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12445_ (.A1(\samples_imag[3][6] ),
    .A2(_03603_),
    .B1(_03605_),
    .B2(\samples_imag[6][6] ),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12446_ (.A1(_03664_),
    .A2(\samples_imag[1][6] ),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12447_ (.A1(_03664_),
    .A2(\samples_imag[4][6] ),
    .B1(_04194_),
    .B2(_03654_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12448_ (.I0(_04193_),
    .I1(_04195_),
    .S(_03600_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12449_ (.A1(_03797_),
    .A2(_04038_),
    .B1(_04192_),
    .B2(_04196_),
    .ZN(_07854_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12450_ (.I0(\samples_imag[4][5] ),
    .I1(\samples_imag[5][5] ),
    .I2(\samples_imag[6][5] ),
    .I3(\samples_imag[7][5] ),
    .S0(_03649_),
    .S1(_03644_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12451_ (.I(\samples_imag[1][5] ),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12452_ (.I0(\samples_imag[2][5] ),
    .I1(\samples_imag[3][5] ),
    .S(_03613_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12453_ (.I(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12454_ (.A1(_04198_),
    .A2(_03648_),
    .B1(_04200_),
    .B2(_03644_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12455_ (.I0(_04197_),
    .I1(_04201_),
    .S(_03654_),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12456_ (.A1(\samples_imag[0][5] ),
    .A2(_03641_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12457_ (.A1(_04202_),
    .A2(_04203_),
    .Z(_07859_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12458_ (.I0(\samples_imag[4][4] ),
    .I1(\samples_imag[5][4] ),
    .I2(\samples_imag[6][4] ),
    .I3(\samples_imag[7][4] ),
    .S0(_03649_),
    .S1(_03644_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12459_ (.I(\samples_imag[1][4] ),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12460_ (.I0(\samples_imag[2][4] ),
    .I1(\samples_imag[3][4] ),
    .S(_03613_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12461_ (.I(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12462_ (.A1(_04205_),
    .A2(_03648_),
    .B1(_04207_),
    .B2(_03644_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12463_ (.I0(_04204_),
    .I1(_04208_),
    .S(_03654_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12464_ (.A1(\samples_imag[0][4] ),
    .A2(_03641_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12465_ (.A1(_04209_),
    .A2(_04210_),
    .Z(_07864_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12466_ (.I0(\samples_imag[4][3] ),
    .I1(\samples_imag[5][3] ),
    .I2(\samples_imag[6][3] ),
    .I3(\samples_imag[7][3] ),
    .S0(_03642_),
    .S1(_03644_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12467_ (.I(\samples_imag[1][3] ),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12468_ (.I0(\samples_imag[2][3] ),
    .I1(\samples_imag[3][3] ),
    .S(_03613_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12469_ (.I(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12470_ (.A1(_04212_),
    .A2(_03648_),
    .B1(_04214_),
    .B2(_03661_),
    .C(_04058_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12471_ (.A1(_04058_),
    .A2(_04211_),
    .B(_04215_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12472_ (.A1(_03836_),
    .A2(_04010_),
    .B(_04216_),
    .ZN(_07869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12473_ (.I0(\samples_imag[6][2] ),
    .I1(\samples_imag[7][2] ),
    .S(_03642_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12474_ (.A1(\samples_imag[1][2] ),
    .A2(_04094_),
    .B1(_04217_),
    .B2(_04011_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12475_ (.A1(\samples_imag[3][2] ),
    .A2(_04015_),
    .B1(_04097_),
    .B2(\samples_imag[5][2] ),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12476_ (.A1(_03599_),
    .A2(\samples_imag[2][2] ),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12477_ (.A1(_03600_),
    .A2(\samples_imag[4][2] ),
    .B1(_04220_),
    .B2(_03617_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12478_ (.I0(_04219_),
    .I1(_04221_),
    .S(_03665_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12479_ (.A1(_03846_),
    .A2(_04010_),
    .B1(_04218_),
    .B2(_04222_),
    .ZN(_07874_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12480_ (.I(_05868_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12481_ (.I(_05885_),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12482_ (.I(_05899_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12483_ (.I(_05911_),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12484_ (.A1(_00011_),
    .A2(_03896_),
    .Z(_05931_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12485_ (.I(_07903_),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12486_ (.I(_05916_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12487_ (.I(_05950_),
    .ZN(_06039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12488_ (.I(_05953_),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12489_ (.I(_05976_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12490_ (.I(_05979_),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12491_ (.I(_07911_),
    .ZN(_07914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12492_ (.I(_05986_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12493_ (.I(_05958_),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12494_ (.I(_06013_),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12495_ (.I(_06076_),
    .ZN(_06072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12496_ (.I(_06064_),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12497_ (.I(_07917_),
    .ZN(_07921_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12498_ (.I(_06075_),
    .ZN(_06078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12499_ (.I(_06084_),
    .ZN(_06082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12500_ (.I(_06046_),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12501_ (.I(_06097_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12502_ (.I(_06122_),
    .ZN(_06118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12503_ (.I(_06117_),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12504_ (.I(_07893_),
    .ZN(_07935_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12505_ (.I(_06121_),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12506_ (.I(_06133_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12507_ (.I(_06137_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12508_ (.I(_06145_),
    .ZN(_07925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12509_ (.I(_06147_),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12510_ (.I(_06168_),
    .ZN(_06217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12511_ (.I(_07957_),
    .ZN(_07946_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12512_ (.I(_06178_),
    .ZN(_07951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12513_ (.I(_06179_),
    .ZN(_06188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12514_ (.I(_06193_),
    .ZN(_06191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12515_ (.I(_06197_),
    .ZN(_06195_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12516_ (.I(_06207_),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12517_ (.I(_07967_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12518_ (.I(_06228_),
    .ZN(_07962_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12519_ (.I(_06229_),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12520_ (.I(_06243_),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12521_ (.I(_06247_),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12522_ (.I(_06280_),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12523_ (.I(_05912_),
    .ZN(_07897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12524_ (.I(_06294_),
    .ZN(_06291_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12525_ (.I(_07978_),
    .ZN(_06318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12526_ (.I(_05954_),
    .ZN(_07904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12527_ (.I(_06426_),
    .ZN(_06422_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12528_ (.I(_06379_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12529_ (.I(_07993_),
    .ZN(_06354_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12530_ (.I(_08011_),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12531_ (.I(_06336_),
    .ZN(_06366_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12532_ (.I(_06402_),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12533_ (.I(_08009_),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12534_ (.I(_07928_),
    .ZN(_08013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12535_ (.I(_06373_),
    .ZN(_06393_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12536_ (.I(_06433_),
    .ZN(_06428_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12537_ (.I(_08024_),
    .ZN(_08027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12538_ (.I(_06420_),
    .ZN(_06417_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12539_ (.I(_08035_),
    .ZN(_08037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12540_ (.I(_08031_),
    .ZN(_06447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12541_ (.I0(_03845_),
    .I1(_08035_),
    .S(_03817_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12542_ (.A1(_03740_),
    .A2(_04223_),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12543_ (.I(_08032_),
    .ZN(_08045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12544_ (.I(_08058_),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12545_ (.I(_08051_),
    .ZN(_08070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12546_ (.I(_06299_),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12547_ (.I(_06465_),
    .ZN(_06482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12548_ (.I(_06474_),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12549_ (.I(_06475_),
    .ZN(_06484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12550_ (.I(_08081_),
    .ZN(_08079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12551_ (.I(_06524_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12552_ (.I(_06514_),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12553_ (.I(_06549_),
    .ZN(_06572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12554_ (.A1(_03898_),
    .A2(_03714_),
    .Z(_08114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12555_ (.I(_06581_),
    .ZN(_06591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12556_ (.I(_06571_),
    .ZN(_08119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12557_ (.I(_06579_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _12558_ (.I(_03897_),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12559_ (.A1(_04224_),
    .A2(_03739_),
    .Z(_08123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12560_ (.I(_06640_),
    .ZN(_06650_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12561_ (.I(_06615_),
    .ZN(_08137_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12562_ (.I(_06634_),
    .ZN(_08141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12563_ (.I(_06639_),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12564_ (.I(_06630_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12565_ (.A1(_04224_),
    .A2(_03750_),
    .Z(_08144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12566_ (.I(_06670_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12567_ (.I(_06690_),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12568_ (.A1(_04224_),
    .A2(_03771_),
    .Z(_08156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12569_ (.I(_06721_),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12570_ (.I(_06723_),
    .ZN(_08166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12571_ (.I(_06744_),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12572_ (.A1(_04224_),
    .A2(_03789_),
    .Z(_08169_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12573_ (.I(_06801_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12574_ (.I(_06769_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12575_ (.I(_06772_),
    .ZN(_08179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12576_ (.I(_06732_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12577_ (.I(_06800_),
    .ZN(_06850_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12578_ (.A1(_04224_),
    .A2(_03796_),
    .Z(_08184_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12579_ (.I(_06858_),
    .ZN(_06860_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12580_ (.I(_06813_),
    .ZN(_06826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12581_ (.I(_06784_),
    .ZN(_06835_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12582_ (.I(_06802_),
    .ZN(_06852_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12583_ (.A1(_04224_),
    .A2(_03809_),
    .Z(_08199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12584_ (.I(_06872_),
    .ZN(_08202_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12585_ (.I(_06899_),
    .ZN(_08210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12586_ (.A1(_04224_),
    .A2(_03835_),
    .Z(_08215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12587_ (.I(_06944_),
    .ZN(_06946_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12588_ (.I(_06911_),
    .ZN(_06921_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12589_ (.I(_06920_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12590_ (.I(_06891_),
    .ZN(_06930_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12591_ (.I(_06912_),
    .ZN(_06941_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12592_ (.I(_06902_),
    .ZN(_08223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12593_ (.A1(_04224_),
    .A2(_03817_),
    .Z(_08229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12594_ (.I(_06954_),
    .ZN(_06963_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12595_ (.I(_06938_),
    .ZN(_06972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12596_ (.I(_06955_),
    .ZN(_06983_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12597_ (.A1(_04224_),
    .A2(_03845_),
    .Z(_08240_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12598_ (.I(_06994_),
    .ZN(_08248_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12599_ (.I(_07000_),
    .ZN(_08252_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12600_ (.I(_06980_),
    .ZN(_07006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12601_ (.I(_07001_),
    .ZN(_07011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12602_ (.A1(_04224_),
    .A2(_03854_),
    .Z(_08258_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12603_ (.I(_07021_),
    .ZN(_08267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12604_ (.A1(_03897_),
    .A2(_03875_),
    .Z(_08272_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12605_ (.I(_07042_),
    .ZN(_07049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12606_ (.I(_07043_),
    .ZN(_07052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12607_ (.A1(_03897_),
    .A2(_03925_),
    .Z(_08303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12608_ (.A1(_00701_),
    .A2(_00697_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12609_ (.A1(_00588_),
    .A2(_00579_),
    .A3(_00586_),
    .B(_04225_),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12610_ (.A1(_00709_),
    .A2(_00713_),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12611_ (.A1(_00826_),
    .A2(_07095_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12612_ (.A1(_00834_),
    .A2(_04226_),
    .Z(_07107_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12613_ (.I(_00927_),
    .ZN(_07113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12614_ (.I0(_00721_),
    .I1(_07104_),
    .S(_00616_),
    .Z(_07124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12615_ (.I(_00836_),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12616_ (.I(_00648_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12617_ (.I0(_07110_),
    .I1(_04227_),
    .S(_00693_),
    .Z(_07130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12618_ (.I(_00928_),
    .ZN(_07133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12619_ (.A1(_00626_),
    .A2(_07124_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12620_ (.A1(_00687_),
    .A2(_04228_),
    .ZN(_07137_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12621_ (.A1(_00645_),
    .A2(_00836_),
    .B(_00839_),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12622_ (.A1(_00640_),
    .A2(_00649_),
    .A3(_00667_),
    .Z(_07143_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12623_ (.A1(_00645_),
    .A2(_00928_),
    .B(_00932_),
    .ZN(_07146_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12624_ (.A1(_00889_),
    .A2(_00859_),
    .A3(_00862_),
    .Z(_07178_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12625_ (.A1(_00812_),
    .A2(_00809_),
    .Z(_07181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12626_ (.I(_00974_),
    .ZN(_07184_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12627_ (.A1(_07176_),
    .A2(_01001_),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12628_ (.I(_02319_),
    .ZN(_07438_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12629_ (.I(_02896_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12630_ (.A1(_03484_),
    .A2(_03555_),
    .Z(_04229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12631_ (.I(_07645_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12632_ (.A1(_07647_),
    .A2(_07638_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12633_ (.A1(_03556_),
    .A2(_04231_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12634_ (.A1(_04229_),
    .A2(_04230_),
    .B(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12635_ (.I(_04233_),
    .ZN(_07681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12636_ (.A1(_03433_),
    .A2(_03449_),
    .A3(_03483_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12637_ (.A1(_03514_),
    .A2(_03538_),
    .A3(_03554_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12638_ (.A1(\butterfly_count[1] ),
    .A2(_04234_),
    .A3(_04235_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12639_ (.A1(_04234_),
    .A2(_04235_),
    .B(_07639_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12640_ (.A1(_04236_),
    .A2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12641_ (.I(_04238_),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12642_ (.I(_07704_),
    .ZN(_07702_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12643_ (.A1(_07740_),
    .A2(_07745_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12644_ (.A1(_07702_),
    .A2(_05857_),
    .A3(_07691_),
    .A4(_07715_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12645_ (.A1(_07730_),
    .A2(_07760_),
    .A3(_04240_),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12646_ (.A1(_07696_),
    .A2(_07720_),
    .A3(_07725_),
    .A4(_07735_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12647_ (.A1(_07755_),
    .A2(_04239_),
    .A3(_04241_),
    .A4(_04242_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12648_ (.A1(_07706_),
    .A2(_07710_),
    .A3(_07750_),
    .A4(_04243_),
    .Z(_07707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12649_ (.I(_07785_),
    .ZN(_07788_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12650_ (.I(\sample_count[1] ),
    .ZN(_07798_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12651_ (.I(_07687_),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12652_ (.I(_07818_),
    .ZN(_07816_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12653_ (.A1(_07810_),
    .A2(_07820_),
    .A3(_07824_),
    .A4(_07829_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12654_ (.A1(_07839_),
    .A2(_07844_),
    .A3(_07849_),
    .A4(_07874_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12655_ (.A1(_07854_),
    .A2(_07859_),
    .A3(_07864_),
    .A4(_07869_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12656_ (.A1(_04245_),
    .A2(_04246_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12657_ (.A1(_07805_),
    .A2(_07834_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12658_ (.A1(_07818_),
    .A2(_05868_),
    .A3(_04247_),
    .A4(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12659_ (.A1(_04244_),
    .A2(_04249_),
    .Z(_07821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12660_ (.I(_05910_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12661_ (.I(_07895_),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12662_ (.I(_07896_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12663_ (.I(_05952_),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12664_ (.A1(_03897_),
    .A2(_03700_),
    .Z(_05923_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12665_ (.I(_05970_),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12666_ (.I(_07907_),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12667_ (.A1(_03897_),
    .A2(_03779_),
    .Z(_06050_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12668_ (.I(_05991_),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12669_ (.I(_06015_),
    .ZN(_06061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12670_ (.I(_06096_),
    .ZN(_06090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12671_ (.I(_07919_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12672_ (.I(_07930_),
    .ZN(_06044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12673_ (.A1(_03897_),
    .A2(_03827_),
    .Z(_06103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12674_ (.I(_06110_),
    .ZN(_06107_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12675_ (.I(_06071_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12676_ (.I(_07892_),
    .ZN(_07923_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12677_ (.I(_06146_),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12678_ (.I(_06161_),
    .ZN(_06158_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12679_ (.I(_07944_),
    .ZN(_07936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12680_ (.I(_06206_),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12681_ (.A1(_03897_),
    .A2(_03896_),
    .Z(_06213_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12682_ (.I(_07945_),
    .ZN(_07947_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12683_ (.A1(_03897_),
    .A2(_03907_),
    .Z(_06263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12684_ (.I(_07958_),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12685_ (.A1(_03897_),
    .A2(_03915_),
    .Z(_06310_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12686_ (.I(_06293_),
    .ZN(_06290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12687_ (.I(_06274_),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12688_ (.I(_07968_),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12689_ (.I(_06342_),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12690_ (.I(_07979_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12691_ (.I(_06332_),
    .ZN(_06330_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12692_ (.I(_06427_),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12693_ (.I(_06380_),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12694_ (.I(_07994_),
    .ZN(_06037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12695_ (.I(_06369_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12696_ (.A1(_03898_),
    .A2(_03941_),
    .ZN(_08002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12697_ (.I(_06403_),
    .ZN(_06398_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12698_ (.I(_08012_),
    .ZN(_06091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12699_ (.I(_06396_),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12700_ (.I(_06434_),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12701_ (.I(_06421_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12702_ (.I(_08047_),
    .ZN(_08034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12703_ (.A1(_03726_),
    .A2(_03817_),
    .Z(_08038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12704_ (.I(_08043_),
    .ZN(_06448_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12705_ (.I(_08050_),
    .ZN(_08046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12706_ (.I(_08054_),
    .ZN(_08049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12707_ (.I(_08071_),
    .ZN(_08057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12708_ (.I(_07952_),
    .ZN(_06451_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12709_ (.I(_06461_),
    .ZN(_06459_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12710_ (.I(_08059_),
    .ZN(_08068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12711_ (.I(_06468_),
    .ZN(_06253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12712_ (.I(_06486_),
    .ZN(_06483_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12713_ (.I(_06494_),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12714_ (.I(_08080_),
    .ZN(_08087_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12715_ (.A1(_08088_),
    .A2(_06337_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12716_ (.A1(_08098_),
    .A2(_04250_),
    .Z(_08095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12717_ (.A1(_03715_),
    .A2(_03925_),
    .Z(_06502_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12718_ (.I(_06548_),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12719_ (.I(_06536_),
    .ZN(_06538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12720_ (.I(_06570_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12721_ (.I(_06576_),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12722_ (.A1(_03980_),
    .A2(_03979_),
    .Z(_08115_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12723_ (.I(_06633_),
    .ZN(_08120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12724_ (.I(_06638_),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12725_ (.A1(_03980_),
    .A2(_03714_),
    .Z(_08124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12726_ (.I(_06669_),
    .ZN(_06664_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12727_ (.I(_06689_),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12728_ (.A1(_03980_),
    .A2(_03739_),
    .Z(_08145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12729_ (.I(_06720_),
    .ZN(_06716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12730_ (.I(_06743_),
    .ZN(_06741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12731_ (.A1(_03980_),
    .A2(_03750_),
    .Z(_08157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12732_ (.I(_06768_),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12733_ (.I(_06730_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12734_ (.I(_06798_),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12735_ (.A1(_03980_),
    .A2(_03771_),
    .Z(_08170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12736_ (.I(_06824_),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12737_ (.I(_06782_),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12738_ (.I(_06855_),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12739_ (.A1(_03876_),
    .A2(_03789_),
    .Z(_08185_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12740_ (.I(_06818_),
    .ZN(_06827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12741_ (.I(_06871_),
    .ZN(_08187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12742_ (.I(_06839_),
    .ZN(_06836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12743_ (.I(_06898_),
    .ZN(_08194_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12744_ (.A1(_03876_),
    .A2(_03796_),
    .Z(_08200_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12745_ (.I(_06888_),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12746_ (.A1(_03876_),
    .A2(_03809_),
    .Z(_08216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12747_ (.A1(_03876_),
    .A2(_03835_),
    .Z(_08230_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12748_ (.I(_06993_),
    .ZN(_08232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12749_ (.I(_06976_),
    .ZN(_06973_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12750_ (.I(_06945_),
    .ZN(_08237_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12751_ (.A1(_03876_),
    .A2(_03817_),
    .Z(_08241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12752_ (.I(_07020_),
    .ZN(_08255_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12753_ (.A1(_03876_),
    .A2(_03845_),
    .Z(_08259_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12754_ (.A1(_03876_),
    .A2(_03854_),
    .Z(_08273_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12755_ (.I(_07072_),
    .ZN(_08300_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12756_ (.A1(_03876_),
    .A2(_03875_),
    .Z(_08304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12757_ (.I(_08044_),
    .ZN(_08067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12758_ (.I(_08069_),
    .ZN(_08077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12759_ (.I(_08118_),
    .ZN(_06627_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12760_ (.I(_08132_),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12761_ (.I(_08147_),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12762_ (.I(_08159_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12763_ (.I(_08172_),
    .ZN(_06815_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12764_ (.I(_08180_),
    .ZN(_06846_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12765_ (.I(_08245_),
    .ZN(_06998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12766_ (.I(_08284_),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12767_ (.I(_07900_),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12768_ (.I(_07905_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12769_ (.I(_07916_),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12770_ (.I(_07927_),
    .ZN(_06143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12771_ (.I(_07932_),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12772_ (.I(_07940_),
    .ZN(_06203_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12773_ (.I(_07941_),
    .ZN(_06199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12774_ (.I(_07953_),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12775_ (.I(_07955_),
    .ZN(_06271_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12776_ (.I(_08048_),
    .ZN(_08056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12777_ (.I(_08055_),
    .ZN(_08089_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12778_ (.I(_08072_),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12779_ (.I(_08198_),
    .ZN(_06866_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12780_ (.I(_08214_),
    .ZN(_06909_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12781_ (.I(_08228_),
    .ZN(_06952_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12782_ (.I(_07074_),
    .ZN(_07071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12783_ (.I(_08242_),
    .ZN(_07018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12784_ (.I0(\bit_rev_idx[0] ),
    .I1(\sample_count[2] ),
    .S(_03597_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12785_ (.I0(\bit_rev_idx[1] ),
    .I1(\sample_count[1] ),
    .S(_03597_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12786_ (.I0(\bit_rev_idx[2] ),
    .I1(\sample_count[0] ),
    .S(_03597_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12787_ (.I0(_00564_),
    .I1(net83),
    .S(_00565_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12788_ (.A1(_00564_),
    .A2(net83),
    .B1(_04251_),
    .B2(\state[0] ),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12789_ (.I(_04252_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12790_ (.A1(_07686_),
    .A2(_03634_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _12791_ (.I(\state[2] ),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12792_ (.I(\state[1] ),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12793_ (.A1(_04254_),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12794_ (.A1(_03593_),
    .A2(_03991_),
    .A3(_04256_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12795_ (.I0(\butterfly_count[0] ),
    .I1(_04253_),
    .S(_04257_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12796_ (.A1(_07770_),
    .A2(_03634_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12797_ (.I0(\butterfly_count[1] ),
    .I1(_04258_),
    .S(_04257_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12798_ (.A1(_07771_),
    .A2(_03634_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12799_ (.I0(\butterfly_count[2] ),
    .I1(_04259_),
    .S(_04257_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12800_ (.I(\butterfly_in_group[0] ),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12801_ (.I(_03636_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12802_ (.A1(_07685_),
    .A2(_07683_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12803_ (.A1(_07678_),
    .A2(_07682_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12804_ (.I(_07666_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12805_ (.A1(_07674_),
    .A2(_07671_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12806_ (.A1(_04265_),
    .A2(_07670_),
    .B(_07667_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12807_ (.A1(_04266_),
    .A2(_04264_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12808_ (.A1(_04267_),
    .A2(_07663_),
    .B(_07662_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12809_ (.A1(_07689_),
    .A2(_04262_),
    .B(_04263_),
    .C(_04268_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12810_ (.A1(_07683_),
    .A2(_05877_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12811_ (.A1(_04236_),
    .A2(_04237_),
    .B(_04270_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12812_ (.A1(_03419_),
    .A2(_03498_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12813_ (.A1(_03345_),
    .A2(_03364_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12814_ (.A1(_03493_),
    .A2(_03494_),
    .B1(_04272_),
    .B2(_04273_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12815_ (.A1(_03414_),
    .A2(_03486_),
    .B(_03501_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12816_ (.A1(_03501_),
    .A2(_03414_),
    .A3(_03486_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12817_ (.A1(_03372_),
    .A2(_03398_),
    .A3(_03415_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12818_ (.A1(_03345_),
    .A2(_03364_),
    .B(_03392_),
    .C(_04277_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12819_ (.A1(_03392_),
    .A2(_04277_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12820_ (.A1(_04275_),
    .A2(_04276_),
    .A3(_04278_),
    .A4(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _12821_ (.A1(_03345_),
    .A2(_03364_),
    .A3(_03416_),
    .B(_03456_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12822_ (.A1(_03452_),
    .A2(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12823_ (.A1(_03445_),
    .A2(_03447_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12824_ (.A1(_03414_),
    .A2(_03487_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12825_ (.A1(net46),
    .A2(_03426_),
    .B(_04283_),
    .C(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12826_ (.A1(_03421_),
    .A2(_03432_),
    .A3(_04282_),
    .A4(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12827_ (.A1(_03465_),
    .A2(_03467_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12828_ (.A1(_07177_),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12829_ (.A1(_03370_),
    .A2(_03454_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12830_ (.I0(_07630_),
    .I1(_04289_),
    .S(net10),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12831_ (.A1(_07650_),
    .A2(_07639_),
    .A3(_07686_),
    .A4(_07656_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12832_ (.A1(_07647_),
    .A2(_07644_),
    .A3(_07653_),
    .A4(_07659_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12833_ (.A1(_03504_),
    .A2(_04290_),
    .A3(_04291_),
    .A4(_04292_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _12834_ (.A1(_04280_),
    .A2(_04286_),
    .A3(_04288_),
    .A4(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12835_ (.I(_03505_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12836_ (.A1(_04295_),
    .A2(_04275_),
    .A3(_04276_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12837_ (.I(_04296_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12838_ (.A1(_03488_),
    .A2(_03489_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12839_ (.A1(_03433_),
    .A2(_03449_),
    .A3(_03483_),
    .A4(_04298_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12840_ (.A1(_04235_),
    .A2(_04294_),
    .B(_04297_),
    .C(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12841_ (.A1(_04274_),
    .A2(_04300_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12842_ (.A1(_03418_),
    .A2(_03420_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12843_ (.I(_03452_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12844_ (.A1(_04303_),
    .A2(_04281_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12845_ (.A1(_03468_),
    .A2(_03572_),
    .B(_03477_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12846_ (.A1(_07650_),
    .A2(_04305_),
    .B(_07649_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12847_ (.A1(_07177_),
    .A2(_04306_),
    .B(_02196_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12848_ (.A1(_03465_),
    .A2(_03467_),
    .A3(_04307_),
    .Z(_04308_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12849_ (.A1(_03465_),
    .A2(_03467_),
    .B(_04306_),
    .C(_02507_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12850_ (.A1(_04290_),
    .A2(_04308_),
    .A3(_04309_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _12851_ (.A1(_04302_),
    .A2(_04304_),
    .A3(_04283_),
    .A4(_04310_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12852_ (.A1(_04234_),
    .A2(_04235_),
    .B(_04311_),
    .C(_03427_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12853_ (.A1(_03432_),
    .A2(_04312_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12854_ (.A1(_04269_),
    .A2(_04271_),
    .B(_04301_),
    .C(_04313_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12855_ (.A1(_04303_),
    .A2(_04281_),
    .A3(_04310_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12856_ (.A1(_04303_),
    .A2(_04281_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12857_ (.A1(_03445_),
    .A2(_03452_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _12858_ (.A1(_03445_),
    .A2(_04315_),
    .A3(_04316_),
    .B1(_04317_),
    .B2(_04310_),
    .B3(_04281_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12859_ (.A1(_04286_),
    .A2(_04296_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12860_ (.A1(_03345_),
    .A2(_03361_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12861_ (.A1(_03419_),
    .A2(_03498_),
    .B(_03491_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12862_ (.A1(_04272_),
    .A2(_04320_),
    .B(_04321_),
    .C(_03497_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12863_ (.A1(_03516_),
    .A2(_03527_),
    .A3(_04274_),
    .A4(_04322_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12864_ (.A1(_03518_),
    .A2(_03526_),
    .B(_03517_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12865_ (.A1(_03518_),
    .A2(_03526_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12866_ (.A1(_04324_),
    .A2(_04325_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12867_ (.A1(_03534_),
    .A2(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12868_ (.A1(_04310_),
    .A2(_04319_),
    .A3(_04323_),
    .B(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12869_ (.I(_03483_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12870_ (.A1(_03434_),
    .A2(_03436_),
    .B1(_03445_),
    .B2(_04329_),
    .C(_03447_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12871_ (.A1(_03519_),
    .A2(_03534_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12872_ (.A1(_03337_),
    .A2(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12873_ (.I(_03337_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12874_ (.A1(_03335_),
    .A2(_03311_),
    .A3(_03312_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12875_ (.A1(_04333_),
    .A2(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12876_ (.I0(_04332_),
    .I1(_04335_),
    .S(_03526_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12877_ (.A1(_07675_),
    .A2(_07667_),
    .A3(_07671_),
    .A4(_07663_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12878_ (.A1(_07679_),
    .A2(_07678_),
    .B(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12879_ (.A1(_07679_),
    .A2(_07685_),
    .A3(_07683_),
    .A4(_07688_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12880_ (.A1(_04338_),
    .A2(_04268_),
    .B1(_04339_),
    .B2(_04337_),
    .C(_03342_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12881_ (.A1(_04333_),
    .A2(_04334_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12882_ (.A1(_04331_),
    .A2(_04335_),
    .B(_04341_),
    .C(_04340_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12883_ (.A1(_03496_),
    .A2(_03364_),
    .A3(_03416_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12884_ (.A1(_03516_),
    .A2(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12885_ (.A1(_04342_),
    .A2(_04322_),
    .A3(_04302_),
    .A4(_04344_),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12886_ (.A1(_04280_),
    .A2(_04345_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12887_ (.A1(_03547_),
    .A2(_04346_),
    .A3(_04336_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12888_ (.A1(_04318_),
    .A2(_04328_),
    .A3(_04330_),
    .A4(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12889_ (.A1(_03484_),
    .A2(_04298_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _12890_ (.A1(_04287_),
    .A2(_04235_),
    .A3(_04294_),
    .A4(_04327_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12891_ (.A1(_03443_),
    .A2(_03444_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12892_ (.A1(_03501_),
    .A2(_03414_),
    .A3(_03486_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12893_ (.A1(_03504_),
    .A2(_04352_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12894_ (.A1(_04288_),
    .A2(_04306_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12895_ (.A1(_03482_),
    .A2(_03481_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12896_ (.A1(_04290_),
    .A2(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12897_ (.A1(_04351_),
    .A2(_04353_),
    .A3(_04354_),
    .A4(_04356_),
    .Z(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12898_ (.A1(_04349_),
    .A2(_04350_),
    .B1(_04357_),
    .B2(_04229_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12899_ (.A1(_03434_),
    .A2(_03437_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12900_ (.A1(_03440_),
    .A2(_04359_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12901_ (.A1(_03500_),
    .A2(_03530_),
    .A3(_04319_),
    .B(_04360_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12902_ (.A1(_04234_),
    .A2(_04235_),
    .B(_04311_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12903_ (.I0(_04361_),
    .I1(_04360_),
    .S(_04362_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12904_ (.A1(_04304_),
    .A2(_04310_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12905_ (.A1(_03484_),
    .A2(_04298_),
    .B(_03553_),
    .C(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12906_ (.I(_03547_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12907_ (.A1(_03514_),
    .A2(_03538_),
    .A3(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12908_ (.A1(_03553_),
    .A2(_04364_),
    .B(_04367_),
    .C(_03484_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12909_ (.A1(_04365_),
    .A2(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12910_ (.A1(_04363_),
    .A2(_04358_),
    .A3(_04348_),
    .A4(_04369_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12911_ (.I0(_04272_),
    .I1(_03499_),
    .S(_03361_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12912_ (.A1(_03538_),
    .A2(_04274_),
    .A3(_04310_),
    .A4(_04371_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12913_ (.A1(_03484_),
    .A2(_03555_),
    .B(_04319_),
    .C(_04372_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12914_ (.I(_03540_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12915_ (.A1(_03546_),
    .A2(_04373_),
    .B(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12916_ (.A1(_03512_),
    .A2(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12917_ (.A1(_03500_),
    .A2(_03516_),
    .A3(_03530_),
    .A4(_04300_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12918_ (.A1(_03527_),
    .A2(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12919_ (.A1(_04370_),
    .A2(_04314_),
    .A3(_04376_),
    .A4(_04378_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12920_ (.A1(_07688_),
    .A2(_04379_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12921_ (.A1(_04370_),
    .A2(_04314_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12922_ (.A1(_04376_),
    .A2(_04378_),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12923_ (.A1(\butterfly_count[0] ),
    .A2(_04381_),
    .A3(_04382_),
    .B(_04261_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12924_ (.A1(_04260_),
    .A2(_04261_),
    .B1(_04380_),
    .B2(_04383_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _12925_ (.A1(_04314_),
    .A2(_04370_),
    .A3(_04376_),
    .A4(_04378_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12926_ (.A1(_04238_),
    .A2(_04376_),
    .A3(_04378_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12927_ (.A1(_05866_),
    .A2(_04384_),
    .B1(_04381_),
    .B2(_04385_),
    .C(_03636_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12928_ (.A1(\butterfly_in_group[1] ),
    .A2(_03636_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12929_ (.A1(_04387_),
    .A2(_04386_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12930_ (.I(\butterfly_in_group[2] ),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12931_ (.A1(_05865_),
    .A2(_07683_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12932_ (.A1(_04379_),
    .A2(_04389_),
    .Z(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12933_ (.A1(_04233_),
    .A2(_04381_),
    .A3(_04382_),
    .B(_04261_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12934_ (.A1(_04388_),
    .A2(_04261_),
    .B1(_04390_),
    .B2(_04391_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12935_ (.I(_00563_),
    .Z(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12936_ (.I0(net84),
    .I1(\samples_imag[0][0] ),
    .S(_04392_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12937_ (.I0(net85),
    .I1(\samples_imag[6][4] ),
    .S(_04392_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12938_ (.I0(net86),
    .I1(\samples_imag[6][5] ),
    .S(_04392_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12939_ (.I0(net87),
    .I1(\samples_imag[6][6] ),
    .S(_04392_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12940_ (.I0(net88),
    .I1(\samples_imag[6][7] ),
    .S(_04392_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12941_ (.I0(net89),
    .I1(\samples_imag[6][8] ),
    .S(_04392_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12942_ (.I0(net90),
    .I1(\samples_imag[6][9] ),
    .S(_04392_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12943_ (.I0(net91),
    .I1(\samples_imag[6][10] ),
    .S(_04392_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12944_ (.I0(net92),
    .I1(\samples_imag[6][11] ),
    .S(_04392_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _12945_ (.I(_00563_),
    .Z(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12946_ (.I(_04393_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12947_ (.I0(net93),
    .I1(\samples_imag[6][12] ),
    .S(_04394_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12948_ (.I0(net94),
    .I1(\samples_imag[6][13] ),
    .S(_04394_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12949_ (.I0(net95),
    .I1(\samples_imag[0][10] ),
    .S(_04394_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12950_ (.I0(net96),
    .I1(\samples_imag[6][14] ),
    .S(_04394_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12951_ (.I0(net97),
    .I1(\samples_imag[6][15] ),
    .S(_04394_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12952_ (.I0(net98),
    .I1(\samples_imag[7][0] ),
    .S(_04394_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12953_ (.I0(net99),
    .I1(\samples_imag[7][1] ),
    .S(_04394_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12954_ (.I0(net100),
    .I1(\samples_imag[7][2] ),
    .S(_04394_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12955_ (.I0(net101),
    .I1(\samples_imag[7][3] ),
    .S(_04394_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12956_ (.I0(net102),
    .I1(\samples_imag[7][4] ),
    .S(_04394_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12957_ (.I(_04393_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12958_ (.I0(net103),
    .I1(\samples_imag[7][5] ),
    .S(_04395_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12959_ (.I0(net104),
    .I1(\samples_imag[7][6] ),
    .S(_04395_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12960_ (.I0(net105),
    .I1(\samples_imag[7][7] ),
    .S(_04395_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12961_ (.I0(net106),
    .I1(\samples_imag[0][11] ),
    .S(_04395_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12962_ (.I0(net107),
    .I1(\samples_imag[7][8] ),
    .S(_04395_),
    .Z(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12963_ (.I0(net108),
    .I1(\samples_imag[7][9] ),
    .S(_04395_),
    .Z(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12964_ (.I0(net109),
    .I1(\samples_imag[7][10] ),
    .S(_04395_),
    .Z(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12965_ (.I0(net110),
    .I1(\samples_imag[7][11] ),
    .S(_04395_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12966_ (.I0(net111),
    .I1(\samples_imag[7][12] ),
    .S(_04395_),
    .Z(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12967_ (.I0(net112),
    .I1(\samples_imag[7][13] ),
    .S(_04395_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _12968_ (.I(_00563_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12969_ (.I(_04396_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12970_ (.I0(net113),
    .I1(\samples_imag[7][14] ),
    .S(_04397_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12971_ (.I0(net114),
    .I1(\samples_imag[7][15] ),
    .S(_04397_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12972_ (.I0(net115),
    .I1(\samples_imag[0][12] ),
    .S(_04397_),
    .Z(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12973_ (.I0(net116),
    .I1(\samples_imag[0][13] ),
    .S(_04397_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12974_ (.I0(net117),
    .I1(\samples_imag[0][14] ),
    .S(_04397_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12975_ (.I0(net118),
    .I1(\samples_imag[0][15] ),
    .S(_04397_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12976_ (.I0(net119),
    .I1(\samples_imag[1][0] ),
    .S(_04397_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12977_ (.I0(net120),
    .I1(\samples_imag[1][1] ),
    .S(_04397_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12978_ (.I0(net121),
    .I1(\samples_imag[1][2] ),
    .S(_04397_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12979_ (.I0(net122),
    .I1(\samples_imag[1][3] ),
    .S(_04397_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12980_ (.I(_04396_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12981_ (.I0(net123),
    .I1(\samples_imag[0][1] ),
    .S(_04398_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12982_ (.I0(net124),
    .I1(\samples_imag[1][4] ),
    .S(_04398_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12983_ (.I0(net125),
    .I1(\samples_imag[1][5] ),
    .S(_04398_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12984_ (.I0(net126),
    .I1(\samples_imag[1][6] ),
    .S(_04398_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12985_ (.I0(net127),
    .I1(\samples_imag[1][7] ),
    .S(_04398_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12986_ (.I0(net128),
    .I1(\samples_imag[1][8] ),
    .S(_04398_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12987_ (.I0(net129),
    .I1(\samples_imag[1][9] ),
    .S(_04398_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12988_ (.I0(net130),
    .I1(\samples_imag[1][10] ),
    .S(_04398_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12989_ (.I0(net131),
    .I1(\samples_imag[1][11] ),
    .S(_04398_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12990_ (.I0(net132),
    .I1(\samples_imag[1][12] ),
    .S(_04398_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _12991_ (.I(_04396_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12992_ (.I0(net133),
    .I1(\samples_imag[1][13] ),
    .S(_04399_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12993_ (.I0(net134),
    .I1(\samples_imag[0][2] ),
    .S(_04399_),
    .Z(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12994_ (.I0(net135),
    .I1(\samples_imag[1][14] ),
    .S(_04399_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12995_ (.I0(net136),
    .I1(\samples_imag[1][15] ),
    .S(_04399_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12996_ (.I0(net137),
    .I1(\samples_imag[2][0] ),
    .S(_04399_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12997_ (.I0(net138),
    .I1(\samples_imag[2][1] ),
    .S(_04399_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12998_ (.I0(net139),
    .I1(\samples_imag[2][2] ),
    .S(_04399_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12999_ (.I0(net140),
    .I1(\samples_imag[2][3] ),
    .S(_04399_),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13000_ (.I0(net141),
    .I1(\samples_imag[2][4] ),
    .S(_04399_),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13001_ (.I0(net142),
    .I1(\samples_imag[2][5] ),
    .S(_04399_),
    .Z(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13002_ (.I(_04396_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13003_ (.I0(net143),
    .I1(\samples_imag[2][6] ),
    .S(_04400_),
    .Z(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13004_ (.I0(net144),
    .I1(\samples_imag[2][7] ),
    .S(_04400_),
    .Z(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13005_ (.I0(net145),
    .I1(\samples_imag[0][3] ),
    .S(_04400_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13006_ (.I0(net146),
    .I1(\samples_imag[2][8] ),
    .S(_04400_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13007_ (.I0(net147),
    .I1(\samples_imag[2][9] ),
    .S(_04400_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13008_ (.I0(net148),
    .I1(\samples_imag[2][10] ),
    .S(_04400_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13009_ (.I0(net149),
    .I1(\samples_imag[2][11] ),
    .S(_04400_),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13010_ (.I0(net150),
    .I1(\samples_imag[2][12] ),
    .S(_04400_),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13011_ (.I0(net151),
    .I1(\samples_imag[2][13] ),
    .S(_04400_),
    .Z(_00099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13012_ (.I0(net152),
    .I1(\samples_imag[2][14] ),
    .S(_04400_),
    .Z(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13013_ (.I(_04396_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13014_ (.I0(net153),
    .I1(\samples_imag[2][15] ),
    .S(_04401_),
    .Z(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13015_ (.I0(net154),
    .I1(\samples_imag[3][0] ),
    .S(_04401_),
    .Z(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13016_ (.I0(net155),
    .I1(\samples_imag[3][1] ),
    .S(_04401_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13017_ (.I0(net156),
    .I1(\samples_imag[0][4] ),
    .S(_04401_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13018_ (.I0(net157),
    .I1(\samples_imag[3][2] ),
    .S(_04401_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13019_ (.I0(net158),
    .I1(\samples_imag[3][3] ),
    .S(_04401_),
    .Z(_00106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13020_ (.I0(net159),
    .I1(\samples_imag[3][4] ),
    .S(_04401_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13021_ (.I0(net160),
    .I1(\samples_imag[3][5] ),
    .S(_04401_),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13022_ (.I0(net161),
    .I1(\samples_imag[3][6] ),
    .S(_04401_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13023_ (.I0(net162),
    .I1(\samples_imag[3][7] ),
    .S(_04401_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13024_ (.I(_04396_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13025_ (.I0(net163),
    .I1(\samples_imag[3][8] ),
    .S(_04402_),
    .Z(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13026_ (.I0(net164),
    .I1(\samples_imag[3][9] ),
    .S(_04402_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13027_ (.I0(net165),
    .I1(\samples_imag[3][10] ),
    .S(_04402_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13028_ (.I0(net166),
    .I1(\samples_imag[3][11] ),
    .S(_04402_),
    .Z(_00114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13029_ (.I0(net167),
    .I1(\samples_imag[0][5] ),
    .S(_04402_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13030_ (.I0(net168),
    .I1(\samples_imag[3][12] ),
    .S(_04402_),
    .Z(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13031_ (.I0(net169),
    .I1(\samples_imag[3][13] ),
    .S(_04402_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13032_ (.I0(net170),
    .I1(\samples_imag[3][14] ),
    .S(_04402_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13033_ (.I0(net171),
    .I1(\samples_imag[3][15] ),
    .S(_04402_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13034_ (.I0(net172),
    .I1(\samples_imag[4][0] ),
    .S(_04402_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13035_ (.I(_04396_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13036_ (.I0(net173),
    .I1(\samples_imag[4][1] ),
    .S(_04403_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13037_ (.I0(net174),
    .I1(\samples_imag[4][2] ),
    .S(_04403_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13038_ (.I0(net175),
    .I1(\samples_imag[4][3] ),
    .S(_04403_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13039_ (.I0(net176),
    .I1(\samples_imag[4][4] ),
    .S(_04403_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13040_ (.I0(net177),
    .I1(\samples_imag[4][5] ),
    .S(_04403_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13041_ (.I0(net178),
    .I1(\samples_imag[0][6] ),
    .S(_04403_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13042_ (.I0(net179),
    .I1(\samples_imag[4][6] ),
    .S(_04403_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13043_ (.I0(net180),
    .I1(\samples_imag[4][7] ),
    .S(_04403_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13044_ (.I0(net181),
    .I1(\samples_imag[4][8] ),
    .S(_04403_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13045_ (.I0(net182),
    .I1(\samples_imag[4][9] ),
    .S(_04403_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13046_ (.I(_04396_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13047_ (.I0(net183),
    .I1(\samples_imag[4][10] ),
    .S(_04404_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13048_ (.I0(net184),
    .I1(\samples_imag[4][11] ),
    .S(_04404_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13049_ (.I0(net185),
    .I1(\samples_imag[4][12] ),
    .S(_04404_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13050_ (.I0(net186),
    .I1(\samples_imag[4][13] ),
    .S(_04404_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13051_ (.I0(net187),
    .I1(\samples_imag[4][14] ),
    .S(_04404_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13052_ (.I0(net188),
    .I1(\samples_imag[4][15] ),
    .S(_04404_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13053_ (.I0(net189),
    .I1(\samples_imag[0][7] ),
    .S(_04404_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13054_ (.I0(net190),
    .I1(\samples_imag[5][0] ),
    .S(_04404_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13055_ (.I0(net191),
    .I1(\samples_imag[5][1] ),
    .S(_04404_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13056_ (.I0(net192),
    .I1(\samples_imag[5][2] ),
    .S(_04404_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13057_ (.I(_04396_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13058_ (.I0(net193),
    .I1(\samples_imag[5][3] ),
    .S(_04405_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13059_ (.I0(net194),
    .I1(\samples_imag[5][4] ),
    .S(_04405_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13060_ (.I0(net195),
    .I1(\samples_imag[5][5] ),
    .S(_04405_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13061_ (.I0(net196),
    .I1(\samples_imag[5][6] ),
    .S(_04405_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13062_ (.I0(net197),
    .I1(\samples_imag[5][7] ),
    .S(_04405_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13063_ (.I0(net198),
    .I1(\samples_imag[5][8] ),
    .S(_04405_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13064_ (.I0(net199),
    .I1(\samples_imag[5][9] ),
    .S(_04405_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13065_ (.I0(net200),
    .I1(\samples_imag[0][8] ),
    .S(_04405_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13066_ (.I0(net201),
    .I1(\samples_imag[5][10] ),
    .S(_04405_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13067_ (.I0(net202),
    .I1(\samples_imag[5][11] ),
    .S(_04405_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13068_ (.I(_04396_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13069_ (.I0(net203),
    .I1(\samples_imag[5][12] ),
    .S(_04406_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13070_ (.I0(net204),
    .I1(\samples_imag[5][13] ),
    .S(_04406_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13071_ (.I0(net205),
    .I1(\samples_imag[5][14] ),
    .S(_04406_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13072_ (.I0(net206),
    .I1(\samples_imag[5][15] ),
    .S(_04406_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13073_ (.I0(net207),
    .I1(\samples_imag[6][0] ),
    .S(_04406_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13074_ (.I0(net208),
    .I1(\samples_imag[6][1] ),
    .S(_04406_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13075_ (.I0(net209),
    .I1(\samples_imag[6][2] ),
    .S(_04406_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13076_ (.I0(net210),
    .I1(\samples_imag[6][3] ),
    .S(_04406_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13077_ (.I0(net211),
    .I1(\samples_imag[0][9] ),
    .S(_04406_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13078_ (.I0(net212),
    .I1(\samples_real[0][0] ),
    .S(_04406_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13079_ (.I(_00563_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13080_ (.I(_04407_),
    .Z(_04408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13081_ (.I0(net213),
    .I1(\samples_real[6][4] ),
    .S(_04408_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13082_ (.I0(net214),
    .I1(\samples_real[6][5] ),
    .S(_04408_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13083_ (.I0(net215),
    .I1(\samples_real[6][6] ),
    .S(_04408_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13084_ (.I0(net216),
    .I1(\samples_real[6][7] ),
    .S(_04408_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13085_ (.I0(net217),
    .I1(\samples_real[6][8] ),
    .S(_04408_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13086_ (.I0(net218),
    .I1(\samples_real[6][9] ),
    .S(_04408_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13087_ (.I0(net219),
    .I1(\samples_real[6][10] ),
    .S(_04408_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13088_ (.I0(net220),
    .I1(\samples_real[6][11] ),
    .S(_04408_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13089_ (.I0(net221),
    .I1(\samples_real[6][12] ),
    .S(_04408_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13090_ (.I0(net222),
    .I1(\samples_real[6][13] ),
    .S(_04408_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13091_ (.I(_04407_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13092_ (.I0(net223),
    .I1(\samples_real[0][10] ),
    .S(_04409_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13093_ (.I0(net224),
    .I1(\samples_real[6][14] ),
    .S(_04409_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13094_ (.I0(net225),
    .I1(\samples_real[6][15] ),
    .S(_04409_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13095_ (.I0(net226),
    .I1(\samples_real[7][0] ),
    .S(_04409_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13096_ (.I0(net227),
    .I1(\samples_real[7][1] ),
    .S(_04409_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13097_ (.I0(net228),
    .I1(\samples_real[7][2] ),
    .S(_04409_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13098_ (.I0(net229),
    .I1(\samples_real[7][3] ),
    .S(_04409_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13099_ (.I0(net230),
    .I1(\samples_real[7][4] ),
    .S(_04409_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13100_ (.I0(net231),
    .I1(\samples_real[7][5] ),
    .S(_04409_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13101_ (.I0(net232),
    .I1(\samples_real[7][6] ),
    .S(_04409_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13102_ (.I(_04407_),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13103_ (.I0(net233),
    .I1(\samples_real[7][7] ),
    .S(_04410_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13104_ (.I0(net234),
    .I1(\samples_real[0][11] ),
    .S(_04410_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13105_ (.I0(net235),
    .I1(\samples_real[7][8] ),
    .S(_04410_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13106_ (.I0(net236),
    .I1(\samples_real[7][9] ),
    .S(_04410_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13107_ (.I0(net237),
    .I1(\samples_real[7][10] ),
    .S(_04410_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13108_ (.I0(net238),
    .I1(\samples_real[7][11] ),
    .S(_04410_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13109_ (.I0(net239),
    .I1(\samples_real[7][12] ),
    .S(_04410_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13110_ (.I0(net240),
    .I1(\samples_real[7][13] ),
    .S(_04410_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13111_ (.I0(net241),
    .I1(\samples_real[7][14] ),
    .S(_04410_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13112_ (.I0(net242),
    .I1(\samples_real[7][15] ),
    .S(_04410_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13113_ (.I(_04407_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13114_ (.I0(net243),
    .I1(\samples_real[0][12] ),
    .S(_04411_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13115_ (.I0(net244),
    .I1(\samples_real[0][13] ),
    .S(_04411_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13116_ (.I0(net245),
    .I1(\samples_real[0][14] ),
    .S(_04411_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13117_ (.I0(net246),
    .I1(\samples_real[0][15] ),
    .S(_04411_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13118_ (.I0(net247),
    .I1(\samples_real[1][0] ),
    .S(_04411_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13119_ (.I0(net248),
    .I1(\samples_real[1][1] ),
    .S(_04411_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13120_ (.I0(net249),
    .I1(\samples_real[1][2] ),
    .S(_04411_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13121_ (.I0(net250),
    .I1(\samples_real[1][3] ),
    .S(_04411_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13122_ (.I0(net251),
    .I1(\samples_real[0][1] ),
    .S(_04411_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13123_ (.I0(net252),
    .I1(\samples_real[1][4] ),
    .S(_04411_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _13124_ (.I(_04407_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13125_ (.I0(net253),
    .I1(\samples_real[1][5] ),
    .S(_04412_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13126_ (.I0(net254),
    .I1(\samples_real[1][6] ),
    .S(_04412_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13127_ (.I0(net255),
    .I1(\samples_real[1][7] ),
    .S(_04412_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13128_ (.I0(net256),
    .I1(\samples_real[1][8] ),
    .S(_04412_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13129_ (.I0(net257),
    .I1(\samples_real[1][9] ),
    .S(_04412_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13130_ (.I0(net258),
    .I1(\samples_real[1][10] ),
    .S(_04412_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13131_ (.I0(net259),
    .I1(\samples_real[1][11] ),
    .S(_04412_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13132_ (.I0(net260),
    .I1(\samples_real[1][12] ),
    .S(_04412_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13133_ (.I0(net261),
    .I1(\samples_real[1][13] ),
    .S(_04412_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13134_ (.I0(net262),
    .I1(\samples_real[0][2] ),
    .S(_04412_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13135_ (.I(_04407_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13136_ (.I0(net263),
    .I1(\samples_real[1][14] ),
    .S(_04413_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13137_ (.I0(net264),
    .I1(\samples_real[1][15] ),
    .S(_04413_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13138_ (.I0(net265),
    .I1(\samples_real[2][0] ),
    .S(_04413_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13139_ (.I0(net266),
    .I1(\samples_real[2][1] ),
    .S(_04413_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13140_ (.I0(net267),
    .I1(\samples_real[2][2] ),
    .S(_04413_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13141_ (.I0(net268),
    .I1(\samples_real[2][3] ),
    .S(_04413_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13142_ (.I0(net269),
    .I1(\samples_real[2][4] ),
    .S(_04413_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13143_ (.I0(net270),
    .I1(\samples_real[2][5] ),
    .S(_04413_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13144_ (.I0(net271),
    .I1(\samples_real[2][6] ),
    .S(_04413_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13145_ (.I0(net272),
    .I1(\samples_real[2][7] ),
    .S(_04413_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13146_ (.I(_04407_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13147_ (.I0(net273),
    .I1(\samples_real[0][3] ),
    .S(_04414_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13148_ (.I0(net274),
    .I1(\samples_real[2][8] ),
    .S(_04414_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13149_ (.I0(net275),
    .I1(\samples_real[2][9] ),
    .S(_04414_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13150_ (.I0(net276),
    .I1(\samples_real[2][10] ),
    .S(_04414_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13151_ (.I0(net277),
    .I1(\samples_real[2][11] ),
    .S(_04414_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13152_ (.I0(net278),
    .I1(\samples_real[2][12] ),
    .S(_04414_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13153_ (.I0(net279),
    .I1(\samples_real[2][13] ),
    .S(_04414_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13154_ (.I0(net280),
    .I1(\samples_real[2][14] ),
    .S(_04414_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13155_ (.I0(net281),
    .I1(\samples_real[2][15] ),
    .S(_04414_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13156_ (.I0(net282),
    .I1(\samples_real[3][0] ),
    .S(_04414_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13157_ (.I(_04407_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13158_ (.I0(net283),
    .I1(\samples_real[3][1] ),
    .S(_04415_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13159_ (.I0(net284),
    .I1(\samples_real[0][4] ),
    .S(_04415_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13160_ (.I0(net285),
    .I1(\samples_real[3][2] ),
    .S(_04415_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13161_ (.I0(net286),
    .I1(\samples_real[3][3] ),
    .S(_04415_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13162_ (.I0(net287),
    .I1(\samples_real[3][4] ),
    .S(_04415_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13163_ (.I0(net288),
    .I1(\samples_real[3][5] ),
    .S(_04415_),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13164_ (.I0(net289),
    .I1(\samples_real[3][6] ),
    .S(_04415_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13165_ (.I0(net290),
    .I1(\samples_real[3][7] ),
    .S(_04415_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13166_ (.I0(net291),
    .I1(\samples_real[3][8] ),
    .S(_04415_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13167_ (.I0(net292),
    .I1(\samples_real[3][9] ),
    .S(_04415_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13168_ (.I(_04407_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13169_ (.I0(net293),
    .I1(\samples_real[3][10] ),
    .S(_04416_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13170_ (.I0(net294),
    .I1(\samples_real[3][11] ),
    .S(_04416_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13171_ (.I0(net295),
    .I1(\samples_real[0][5] ),
    .S(_04416_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13172_ (.I0(net296),
    .I1(\samples_real[3][12] ),
    .S(_04416_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13173_ (.I0(net297),
    .I1(\samples_real[3][13] ),
    .S(_04416_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13174_ (.I0(net298),
    .I1(\samples_real[3][14] ),
    .S(_04416_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13175_ (.I0(net299),
    .I1(\samples_real[3][15] ),
    .S(_04416_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13176_ (.I0(net300),
    .I1(\samples_real[4][0] ),
    .S(_04416_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13177_ (.I0(net301),
    .I1(\samples_real[4][1] ),
    .S(_04416_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13178_ (.I0(net302),
    .I1(\samples_real[4][2] ),
    .S(_04416_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13179_ (.I(_04407_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13180_ (.I0(net303),
    .I1(\samples_real[4][3] ),
    .S(_04417_),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13181_ (.I0(net304),
    .I1(\samples_real[4][4] ),
    .S(_04417_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13182_ (.I0(net305),
    .I1(\samples_real[4][5] ),
    .S(_04417_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13183_ (.I0(net306),
    .I1(\samples_real[0][6] ),
    .S(_04417_),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13184_ (.I0(net307),
    .I1(\samples_real[4][6] ),
    .S(_04417_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13185_ (.I0(net308),
    .I1(\samples_real[4][7] ),
    .S(_04417_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13186_ (.I0(net309),
    .I1(\samples_real[4][8] ),
    .S(_04417_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13187_ (.I0(net310),
    .I1(\samples_real[4][9] ),
    .S(_04417_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13188_ (.I0(net311),
    .I1(\samples_real[4][10] ),
    .S(_04417_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13189_ (.I0(net312),
    .I1(\samples_real[4][11] ),
    .S(_04417_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13190_ (.I(_00563_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13191_ (.I0(net313),
    .I1(\samples_real[4][12] ),
    .S(_04418_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13192_ (.I0(net314),
    .I1(\samples_real[4][13] ),
    .S(_04418_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13193_ (.I0(net315),
    .I1(\samples_real[4][14] ),
    .S(_04418_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13194_ (.I0(net316),
    .I1(\samples_real[4][15] ),
    .S(_04418_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13195_ (.I0(net317),
    .I1(\samples_real[0][7] ),
    .S(_04418_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13196_ (.I0(net318),
    .I1(\samples_real[5][0] ),
    .S(_04418_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13197_ (.I0(net319),
    .I1(\samples_real[5][1] ),
    .S(_04418_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13198_ (.I0(net320),
    .I1(\samples_real[5][2] ),
    .S(_04418_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13199_ (.I0(net321),
    .I1(\samples_real[5][3] ),
    .S(_04418_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13200_ (.I0(net322),
    .I1(\samples_real[5][4] ),
    .S(_04418_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13201_ (.I(_00563_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13202_ (.I0(net323),
    .I1(\samples_real[5][5] ),
    .S(_04419_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13203_ (.I0(net324),
    .I1(\samples_real[5][6] ),
    .S(_04419_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13204_ (.I0(net325),
    .I1(\samples_real[5][7] ),
    .S(_04419_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13205_ (.I0(net326),
    .I1(\samples_real[5][8] ),
    .S(_04419_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13206_ (.I0(net327),
    .I1(\samples_real[5][9] ),
    .S(_04419_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13207_ (.I0(net328),
    .I1(\samples_real[0][8] ),
    .S(_04419_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13208_ (.I0(net329),
    .I1(\samples_real[5][10] ),
    .S(_04419_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13209_ (.I0(net330),
    .I1(\samples_real[5][11] ),
    .S(_04419_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13210_ (.I0(net331),
    .I1(\samples_real[5][12] ),
    .S(_04419_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13211_ (.I0(net332),
    .I1(\samples_real[5][13] ),
    .S(_04419_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13212_ (.I0(net333),
    .I1(\samples_real[5][14] ),
    .S(_04393_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13213_ (.I0(net334),
    .I1(\samples_real[5][15] ),
    .S(_04393_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13214_ (.I0(net335),
    .I1(\samples_real[6][0] ),
    .S(_04393_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13215_ (.I0(net336),
    .I1(\samples_real[6][1] ),
    .S(_04393_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13216_ (.I0(net337),
    .I1(\samples_real[6][2] ),
    .S(_04393_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13217_ (.I0(net338),
    .I1(\samples_real[6][3] ),
    .S(_04393_),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13218_ (.I0(net339),
    .I1(\samples_real[0][9] ),
    .S(_04393_),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13219_ (.A1(_03591_),
    .A2(_04392_),
    .B(net340),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13220_ (.I0(_04254_),
    .I1(net340),
    .S(_00565_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13221_ (.A1(\state[0] ),
    .A2(_04421_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13222_ (.A1(net340),
    .A2(_03592_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13223_ (.A1(\state[2] ),
    .A2(_04420_),
    .B(_04422_),
    .C(_04423_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13224_ (.I(net341),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13225_ (.I0(net341),
    .I1(_04393_),
    .S(net82),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13226_ (.I(_04425_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13227_ (.A1(_00564_),
    .A2(_04424_),
    .B1(_04426_),
    .B2(\state[0] ),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13228_ (.I0(\group[0] ),
    .I1(_04379_),
    .S(_04261_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13229_ (.I0(\group[1] ),
    .I1(_03556_),
    .S(_04261_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13230_ (.I0(\group[2] ),
    .I1(net10),
    .S(_04261_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13231_ (.I0(_03643_),
    .I1(_00013_),
    .S(_04261_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13232_ (.I0(_03645_),
    .I1(_00014_),
    .S(_04261_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13233_ (.A1(\group[0] ),
    .A2(_07783_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13234_ (.A1(\group[1] ),
    .A2(_07777_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13235_ (.A1(_04427_),
    .A2(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13236_ (.A1(_03670_),
    .A2(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13237_ (.A1(\group[2] ),
    .A2(_02507_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13238_ (.A1(_04430_),
    .A2(_04431_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13239_ (.A1(_03669_),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13240_ (.A1(\butterfly_in_group[2] ),
    .A2(_07886_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _13241_ (.A1(_07889_),
    .A2(_07891_),
    .A3(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13242_ (.A1(_04433_),
    .A2(_04435_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13243_ (.I(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13244_ (.I0(_04058_),
    .I1(_04437_),
    .S(_04261_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13245_ (.I0(_03730_),
    .I1(_00015_),
    .S(_03636_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13246_ (.I(_05880_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13247_ (.I0(_03673_),
    .I1(_04438_),
    .S(_03636_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _13248_ (.A1(_05879_),
    .A2(_07680_),
    .A3(_04436_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13249_ (.I0(_03731_),
    .I1(_04439_),
    .S(_03636_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13250_ (.I(_07803_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13251_ (.A1(\state[2] ),
    .A2(_04440_),
    .A3(_07797_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13252_ (.A1(_03595_),
    .A2(_07789_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13253_ (.A1(\state[0] ),
    .A2(_04256_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13254_ (.A1(_04254_),
    .A2(net80),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13255_ (.A1(_00566_),
    .A2(_04442_),
    .A3(_04443_),
    .A4(_04444_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13256_ (.I0(\sample_count[0] ),
    .I1(_04441_),
    .S(_04445_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13257_ (.A1(\state[2] ),
    .A2(_04440_),
    .A3(_07800_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13258_ (.I0(\sample_count[1] ),
    .I1(_04446_),
    .S(_04445_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13259_ (.A1(\state[2] ),
    .A2(_07804_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13260_ (.I0(\sample_count[2] ),
    .I1(_04447_),
    .S(_04445_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13261_ (.I(_07817_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13262_ (.A1(\temp_imag[0] ),
    .A2(_07820_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13263_ (.I(_07812_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13264_ (.I(_07831_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13265_ (.I(_07841_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13266_ (.I(_07851_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13267_ (.I(_07861_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13268_ (.I(_07871_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13269_ (.I(_07880_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13270_ (.A1(_04456_),
    .A2(_07815_),
    .B(_07881_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13271_ (.I(_07877_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13272_ (.A1(_07876_),
    .A2(_04457_),
    .B(_04458_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13273_ (.A1(_04455_),
    .A2(_04459_),
    .B(_07872_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13274_ (.I(_07867_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13275_ (.A1(_07866_),
    .A2(_04460_),
    .B(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13276_ (.A1(_04454_),
    .A2(_04462_),
    .B(_07862_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13277_ (.I(_07857_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13278_ (.A1(_07856_),
    .A2(_04463_),
    .B(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13279_ (.A1(_04453_),
    .A2(_04465_),
    .B(_07852_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13280_ (.I(_07847_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13281_ (.A1(_07846_),
    .A2(_04466_),
    .B(_04467_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13282_ (.A1(_04452_),
    .A2(_04468_),
    .B(_07842_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13283_ (.I(_07837_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13284_ (.A1(_07836_),
    .A2(_04469_),
    .B(_04470_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13285_ (.A1(_04451_),
    .A2(_04471_),
    .B(_07832_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13286_ (.I(_07827_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13287_ (.A1(_07826_),
    .A2(_04472_),
    .B(_04473_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13288_ (.A1(_04450_),
    .A2(_04474_),
    .B(_07813_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13289_ (.I(_07808_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13290_ (.A1(_07807_),
    .A2(_04475_),
    .B(_04476_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13291_ (.A1(_04449_),
    .A2(_04477_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13292_ (.A1(_07876_),
    .A2(_05870_),
    .B(_04458_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13293_ (.A1(_04455_),
    .A2(_04479_),
    .B(_07872_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13294_ (.A1(_07866_),
    .A2(_04480_),
    .B(_04461_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13295_ (.A1(_04454_),
    .A2(_04481_),
    .B(_07862_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13296_ (.A1(_07856_),
    .A2(_04482_),
    .B(_04464_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13297_ (.A1(_04453_),
    .A2(_04483_),
    .B(_07852_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13298_ (.A1(_07846_),
    .A2(_04484_),
    .B(_04467_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13299_ (.A1(_04452_),
    .A2(_04485_),
    .B(_07842_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13300_ (.A1(_07836_),
    .A2(_04486_),
    .B(_04470_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13301_ (.A1(_04451_),
    .A2(_04487_),
    .B(_07832_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13302_ (.A1(_07826_),
    .A2(_04488_),
    .B(_04473_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13303_ (.A1(_04450_),
    .A2(_04489_),
    .B(_07813_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13304_ (.A1(_07807_),
    .A2(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13305_ (.A1(_04450_),
    .A2(_04474_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13306_ (.A1(_04452_),
    .A2(_04468_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13307_ (.A1(_07856_),
    .A2(_04482_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13308_ (.A1(_04454_),
    .A2(_04462_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13309_ (.A1(_04455_),
    .A2(_04459_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13310_ (.A1(_07876_),
    .A2(_05870_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13311_ (.A1(_07866_),
    .A2(_04480_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13312_ (.A1(_05871_),
    .A2(_04448_),
    .A3(_04497_),
    .A4(_04498_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13313_ (.A1(_04494_),
    .A2(_04495_),
    .A3(_04496_),
    .A4(_04499_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13314_ (.A1(_07846_),
    .A2(_04484_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13315_ (.A1(_04453_),
    .A2(_04465_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13316_ (.A1(_07836_),
    .A2(_04486_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13317_ (.A1(_04500_),
    .A2(_04501_),
    .A3(_04502_),
    .A4(_04503_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13318_ (.A1(_07826_),
    .A2(_04488_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13319_ (.A1(_04451_),
    .A2(_04471_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13320_ (.A1(_04493_),
    .A2(_04504_),
    .A3(_04505_),
    .A4(_04506_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13321_ (.A1(_04491_),
    .A2(_04492_),
    .A3(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13322_ (.A1(\temp_imag[0] ),
    .A2(_07822_),
    .A3(_04508_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13323_ (.A1(_04478_),
    .A2(_04509_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13324_ (.A1(_04448_),
    .A2(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13325_ (.A1(\butterfly_count[2] ),
    .A2(_03990_),
    .B(_03594_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13326_ (.A1(_04256_),
    .A2(_04444_),
    .A3(_04512_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13327_ (.I(\sample_count[2] ),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13328_ (.A1(_04514_),
    .A2(_07799_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13329_ (.A1(_04254_),
    .A2(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13330_ (.A1(\bit_rev_idx[1] ),
    .A2(\bit_rev_idx[0] ),
    .A3(\bit_rev_idx[2] ),
    .B(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13331_ (.A1(_04513_),
    .A2(_04517_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13332_ (.A1(_04010_),
    .A2(_04518_),
    .Z(_04519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13333_ (.A1(\samples_imag[0][0] ),
    .A2(_03641_),
    .B1(_04511_),
    .B2(_04519_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13334_ (.I(_07811_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13335_ (.I(_07825_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13336_ (.I(_07835_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13337_ (.I(_07845_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13338_ (.I(_07855_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13339_ (.I(_07865_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13340_ (.I(_07875_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13341_ (.A1(_07880_),
    .A2(_05873_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13342_ (.A1(_07879_),
    .A2(_04528_),
    .B(_07876_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13343_ (.A1(_04527_),
    .A2(_04529_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13344_ (.A1(_07871_),
    .A2(_04530_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13345_ (.A1(_07870_),
    .A2(_04531_),
    .B(_07866_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13346_ (.A1(_04526_),
    .A2(_04532_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13347_ (.A1(_07861_),
    .A2(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13348_ (.A1(_07860_),
    .A2(_04534_),
    .B(_07856_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13349_ (.A1(_04525_),
    .A2(_04535_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13350_ (.A1(_07851_),
    .A2(_04536_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13351_ (.A1(_07850_),
    .A2(_04537_),
    .B(_07846_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13352_ (.A1(_04524_),
    .A2(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13353_ (.A1(_07841_),
    .A2(_04539_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13354_ (.A1(_07840_),
    .A2(_04540_),
    .B(_07836_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13355_ (.A1(_04523_),
    .A2(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13356_ (.A1(_07831_),
    .A2(_04542_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13357_ (.A1(_07830_),
    .A2(_04543_),
    .B(_07826_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13358_ (.A1(_04522_),
    .A2(_04544_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13359_ (.A1(_07812_),
    .A2(_04545_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13360_ (.A1(_04521_),
    .A2(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13361_ (.A1(_07807_),
    .A2(_04547_),
    .B(_07806_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13362_ (.A1(_04449_),
    .A2(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _13363_ (.A1(\temp_imag[0] ),
    .A2(_07823_),
    .A3(_04549_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _13364_ (.I(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13365_ (.A1(_07817_),
    .A2(_04551_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13366_ (.A1(_03728_),
    .A2(_04518_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _13367_ (.A1(_03728_),
    .A2(_04520_),
    .B1(_04552_),
    .B2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13368_ (.A1(_03596_),
    .A2(_04554_),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13369_ (.A1(_04255_),
    .A2(net48),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13370_ (.I0(\samples_imag[0][0] ),
    .I1(_04556_),
    .S(_04518_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13371_ (.A1(_04555_),
    .A2(_04557_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13372_ (.A1(_07876_),
    .A2(_05874_),
    .B(_07875_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13373_ (.I(_07870_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13374_ (.A1(_04455_),
    .A2(_04558_),
    .B(_04559_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13375_ (.A1(_07866_),
    .A2(_04560_),
    .B(_07865_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13376_ (.I(_07860_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13377_ (.A1(_04454_),
    .A2(_04561_),
    .B(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13378_ (.A1(_07856_),
    .A2(_04563_),
    .B(_07855_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13379_ (.I(_07850_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13380_ (.A1(_04453_),
    .A2(_04564_),
    .B(_04565_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13381_ (.A1(_07846_),
    .A2(_04566_),
    .B(_07845_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13382_ (.I(_07840_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13383_ (.A1(_04452_),
    .A2(_04567_),
    .B(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13384_ (.A1(_07836_),
    .A2(_04569_),
    .Z(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13385_ (.A1(_04551_),
    .A2(_04570_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13386_ (.I(_04510_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13387_ (.A1(_04503_),
    .A2(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13388_ (.I(_04008_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13389_ (.I0(\samples_imag[0][10] ),
    .I1(_04573_),
    .S(_04574_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13390_ (.I0(_04571_),
    .I1(_04575_),
    .S(_03905_),
    .Z(_04576_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13391_ (.I(_03594_),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13392_ (.I(_04577_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13393_ (.I0(net49),
    .I1(_04576_),
    .S(_04578_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13394_ (.I(_04518_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13395_ (.I0(\samples_imag[0][10] ),
    .I1(_04579_),
    .S(_04580_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13396_ (.A1(_07831_),
    .A2(_04542_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _13397_ (.I(_04550_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13398_ (.A1(_07831_),
    .A2(_04542_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13399_ (.A1(_04581_),
    .A2(_04582_),
    .A3(_04583_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13400_ (.A1(_04506_),
    .A2(_04572_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13401_ (.I0(\samples_imag[0][11] ),
    .I1(_04585_),
    .S(_04574_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13402_ (.I0(_04584_),
    .I1(_04586_),
    .S(_03905_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13403_ (.I0(net50),
    .I1(_04587_),
    .S(_04578_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13404_ (.I0(\samples_imag[0][11] ),
    .I1(_04588_),
    .S(_04580_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13405_ (.A1(_07836_),
    .A2(_04569_),
    .B(_07835_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13406_ (.I(_07830_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13407_ (.A1(_04451_),
    .A2(_04589_),
    .B(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13408_ (.A1(_07826_),
    .A2(_04591_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13409_ (.A1(_07826_),
    .A2(_04591_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13410_ (.A1(_04582_),
    .A2(_04592_),
    .A3(_04593_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13411_ (.A1(_04505_),
    .A2(_04572_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13412_ (.I0(\samples_imag[0][12] ),
    .I1(_04595_),
    .S(_04574_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13413_ (.I0(_04594_),
    .I1(_04596_),
    .S(_03905_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13414_ (.I(_04577_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13415_ (.I0(net51),
    .I1(_04597_),
    .S(_04598_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13416_ (.I0(\samples_imag[0][12] ),
    .I1(_04599_),
    .S(_04580_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13417_ (.A1(_07812_),
    .A2(_04545_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13418_ (.A1(_04546_),
    .A2(_04582_),
    .A3(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13419_ (.A1(_04492_),
    .A2(_04572_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13420_ (.I0(\samples_imag[0][13] ),
    .I1(_04602_),
    .S(_04574_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13421_ (.I0(_04601_),
    .I1(_04603_),
    .S(_03905_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13422_ (.I0(net52),
    .I1(_04604_),
    .S(_04598_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13423_ (.I0(\samples_imag[0][13] ),
    .I1(_04605_),
    .S(_04580_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13424_ (.A1(_04522_),
    .A2(_04593_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13425_ (.A1(_07812_),
    .A2(_04606_),
    .B(_07811_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13426_ (.A1(_07807_),
    .A2(_04607_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13427_ (.A1(_04551_),
    .A2(_04608_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13428_ (.A1(_04491_),
    .A2(_04572_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13429_ (.I0(\samples_imag[0][14] ),
    .I1(_04610_),
    .S(_04574_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13430_ (.I0(_04609_),
    .I1(_04611_),
    .S(_03905_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13431_ (.I0(net53),
    .I1(_04612_),
    .S(_04598_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13432_ (.I0(\samples_imag[0][14] ),
    .I1(_04613_),
    .S(_04580_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13433_ (.I(_04509_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13434_ (.A1(_04478_),
    .A2(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13435_ (.I0(\samples_imag[0][15] ),
    .I1(_04615_),
    .S(_04574_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13436_ (.I0(_04549_),
    .I1(_04616_),
    .S(_03905_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13437_ (.I0(net54),
    .I1(_04617_),
    .S(_04598_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13438_ (.I0(\samples_imag[0][15] ),
    .I1(_04618_),
    .S(_04580_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13439_ (.I(_05875_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13440_ (.A1(_04619_),
    .A2(_04582_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13441_ (.A1(_05871_),
    .A2(_04572_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13442_ (.I0(\samples_imag[0][1] ),
    .I1(_04621_),
    .S(_04574_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13443_ (.I0(_04620_),
    .I1(_04622_),
    .S(_03905_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13444_ (.I0(net55),
    .I1(_04623_),
    .S(_04598_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13445_ (.I0(\samples_imag[0][1] ),
    .I1(_04624_),
    .S(_04580_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13446_ (.A1(_07876_),
    .A2(_05874_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13447_ (.A1(_04551_),
    .A2(_04625_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13448_ (.A1(_04497_),
    .A2(_04572_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13449_ (.I0(\samples_imag[0][2] ),
    .I1(_04627_),
    .S(_04574_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13450_ (.I0(_04626_),
    .I1(_04628_),
    .S(_03905_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13451_ (.I0(net56),
    .I1(_04629_),
    .S(_04598_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13452_ (.I0(\samples_imag[0][2] ),
    .I1(_04630_),
    .S(_04580_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13453_ (.A1(_04455_),
    .A2(_04530_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13454_ (.A1(_04582_),
    .A2(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13455_ (.A1(_04496_),
    .A2(_04572_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13456_ (.I0(\samples_imag[0][3] ),
    .I1(_04633_),
    .S(_04574_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13457_ (.I(_03712_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13458_ (.I0(_04632_),
    .I1(_04634_),
    .S(_04635_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13459_ (.I0(net57),
    .I1(_04636_),
    .S(_04598_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13460_ (.I0(\samples_imag[0][3] ),
    .I1(_04637_),
    .S(_04580_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13461_ (.A1(_07866_),
    .A2(_04560_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13462_ (.A1(_04582_),
    .A2(_04638_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13463_ (.A1(_04498_),
    .A2(_04572_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13464_ (.I0(\samples_imag[0][4] ),
    .I1(_04640_),
    .S(_04574_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13465_ (.I0(_04639_),
    .I1(_04641_),
    .S(_04635_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13466_ (.I0(net58),
    .I1(_04642_),
    .S(_04598_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13467_ (.I0(\samples_imag[0][4] ),
    .I1(_04643_),
    .S(_04580_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13468_ (.A1(_07861_),
    .A2(_04533_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13469_ (.A1(_07861_),
    .A2(_04533_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13470_ (.A1(_04644_),
    .A2(_04582_),
    .A3(_04645_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13471_ (.A1(_04495_),
    .A2(_04572_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13472_ (.I(_04008_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13473_ (.I0(\samples_imag[0][5] ),
    .I1(_04647_),
    .S(_04648_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13474_ (.I0(_04646_),
    .I1(_04649_),
    .S(_04635_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13475_ (.I0(net59),
    .I1(_04650_),
    .S(_04598_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13476_ (.I(_04518_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13477_ (.I0(\samples_imag[0][5] ),
    .I1(_04651_),
    .S(_04652_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13478_ (.A1(_07856_),
    .A2(_04563_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13479_ (.A1(_04582_),
    .A2(_04653_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13480_ (.A1(_04494_),
    .A2(_04510_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13481_ (.I0(\samples_imag[0][6] ),
    .I1(_04655_),
    .S(_04648_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13482_ (.I0(_04654_),
    .I1(_04656_),
    .S(_04635_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13483_ (.I0(net60),
    .I1(_04657_),
    .S(_04598_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13484_ (.I0(\samples_imag[0][6] ),
    .I1(_04658_),
    .S(_04652_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13485_ (.A1(_07851_),
    .A2(_04536_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13486_ (.A1(_07851_),
    .A2(_04536_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13487_ (.A1(_04659_),
    .A2(_04582_),
    .A3(_04660_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13488_ (.A1(_04502_),
    .A2(_04510_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13489_ (.I0(\samples_imag[0][7] ),
    .I1(_04662_),
    .S(_04648_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13490_ (.I0(_04661_),
    .I1(_04663_),
    .S(_04635_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13491_ (.I(_04577_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13492_ (.I0(net61),
    .I1(_04664_),
    .S(_04665_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13493_ (.I0(\samples_imag[0][7] ),
    .I1(_04666_),
    .S(_04652_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13494_ (.A1(_07846_),
    .A2(_04566_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13495_ (.A1(_04582_),
    .A2(_04667_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13496_ (.A1(_04501_),
    .A2(_04510_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13497_ (.I0(\samples_imag[0][8] ),
    .I1(_04669_),
    .S(_04648_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13498_ (.I0(_04668_),
    .I1(_04670_),
    .S(_04635_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13499_ (.I0(net62),
    .I1(_04671_),
    .S(_04665_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13500_ (.I0(\samples_imag[0][8] ),
    .I1(_04672_),
    .S(_04652_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13501_ (.A1(_07841_),
    .A2(_04539_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13502_ (.A1(_07841_),
    .A2(_04539_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13503_ (.A1(_04673_),
    .A2(_04550_),
    .A3(_04674_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13504_ (.A1(_04493_),
    .A2(_04510_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13505_ (.I0(\samples_imag[0][9] ),
    .I1(_04676_),
    .S(_04648_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13506_ (.I0(_04675_),
    .I1(_04677_),
    .S(_04635_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13507_ (.I0(net63),
    .I1(_04678_),
    .S(_04665_),
    .Z(_04679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13508_ (.I0(\samples_imag[0][9] ),
    .I1(_04679_),
    .S(_04652_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13509_ (.I(\bit_rev_idx[0] ),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13510_ (.A1(\bit_rev_idx[1] ),
    .A2(_04680_),
    .A3(\bit_rev_idx[2] ),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13511_ (.A1(\state[2] ),
    .A2(_04515_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13512_ (.A1(_04513_),
    .A2(_04682_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13513_ (.A1(_04516_),
    .A2(_04681_),
    .B(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13514_ (.I(_04684_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13515_ (.I(_04685_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13516_ (.A1(_03735_),
    .A2(_03754_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13517_ (.I(_04687_),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13518_ (.A1(_04511_),
    .A2(_04684_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13519_ (.I0(\samples_imag[1][0] ),
    .I1(_04689_),
    .S(_04094_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13520_ (.A1(_07817_),
    .A2(_03755_),
    .A3(_04551_),
    .A4(_04685_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13521_ (.A1(_04688_),
    .A2(_04690_),
    .B(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13522_ (.A1(_04556_),
    .A2(_04686_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13523_ (.A1(_03647_),
    .A2(_04686_),
    .B1(_04692_),
    .B2(_04255_),
    .C(_04693_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13524_ (.I0(\samples_imag[1][10] ),
    .I1(_04573_),
    .S(_04094_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13525_ (.I0(_04571_),
    .I1(_04694_),
    .S(_04688_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13526_ (.I0(net49),
    .I1(_04695_),
    .S(_04665_),
    .Z(_04696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13527_ (.I0(\samples_imag[1][10] ),
    .I1(_04696_),
    .S(_04686_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13528_ (.I0(\samples_imag[1][11] ),
    .I1(_04585_),
    .S(_04094_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13529_ (.I0(_04584_),
    .I1(_04697_),
    .S(_04688_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13530_ (.I0(net50),
    .I1(_04698_),
    .S(_04665_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13531_ (.I0(\samples_imag[1][11] ),
    .I1(_04699_),
    .S(_04686_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13532_ (.I(_04021_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13533_ (.I0(\samples_imag[1][12] ),
    .I1(_04595_),
    .S(_04700_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13534_ (.I0(_04594_),
    .I1(_04701_),
    .S(_04688_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13535_ (.I0(net51),
    .I1(_04702_),
    .S(_04665_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13536_ (.I0(\samples_imag[1][12] ),
    .I1(_04703_),
    .S(_04686_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13537_ (.I0(\samples_imag[1][13] ),
    .I1(_04602_),
    .S(_04700_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13538_ (.I0(_04601_),
    .I1(_04704_),
    .S(_04688_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13539_ (.I0(net52),
    .I1(_04705_),
    .S(_04665_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13540_ (.I0(\samples_imag[1][13] ),
    .I1(_04706_),
    .S(_04686_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13541_ (.I0(\samples_imag[1][14] ),
    .I1(_04610_),
    .S(_04700_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13542_ (.I0(_04609_),
    .I1(_04707_),
    .S(_04688_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13543_ (.I0(net53),
    .I1(_04708_),
    .S(_04665_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13544_ (.I0(\samples_imag[1][14] ),
    .I1(_04709_),
    .S(_04686_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13545_ (.I0(\samples_imag[1][15] ),
    .I1(_04615_),
    .S(_04700_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13546_ (.I0(_04549_),
    .I1(_04710_),
    .S(_04688_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13547_ (.I0(net54),
    .I1(_04711_),
    .S(_04665_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13548_ (.I0(\samples_imag[1][15] ),
    .I1(_04712_),
    .S(_04686_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13549_ (.I0(\samples_imag[1][1] ),
    .I1(_04621_),
    .S(_04700_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13550_ (.I0(_04620_),
    .I1(_04713_),
    .S(_04688_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13551_ (.I0(net55),
    .I1(_04714_),
    .S(_04665_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13552_ (.I(_04685_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13553_ (.I0(\samples_imag[1][1] ),
    .I1(_04715_),
    .S(_04716_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13554_ (.I0(\samples_imag[1][2] ),
    .I1(_04627_),
    .S(_04700_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13555_ (.I0(_04626_),
    .I1(_04717_),
    .S(_04688_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13556_ (.I(_04577_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13557_ (.I0(net56),
    .I1(_04718_),
    .S(_04719_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13558_ (.I0(\samples_imag[1][2] ),
    .I1(_04720_),
    .S(_04716_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13559_ (.I0(\samples_imag[1][3] ),
    .I1(_04633_),
    .S(_04700_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13560_ (.I(_04687_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13561_ (.I0(_04632_),
    .I1(_04721_),
    .S(_04722_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13562_ (.I0(net57),
    .I1(_04723_),
    .S(_04719_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13563_ (.I0(\samples_imag[1][3] ),
    .I1(_04724_),
    .S(_04716_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13564_ (.I0(\samples_imag[1][4] ),
    .I1(_04640_),
    .S(_04700_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13565_ (.I0(_04639_),
    .I1(_04725_),
    .S(_04722_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13566_ (.I0(net58),
    .I1(_04726_),
    .S(_04719_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13567_ (.I0(\samples_imag[1][4] ),
    .I1(_04727_),
    .S(_04716_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13568_ (.I0(\samples_imag[1][5] ),
    .I1(_04647_),
    .S(_04700_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13569_ (.I0(_04646_),
    .I1(_04728_),
    .S(_04722_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13570_ (.I0(net59),
    .I1(_04729_),
    .S(_04719_),
    .Z(_04730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13571_ (.I0(\samples_imag[1][5] ),
    .I1(_04730_),
    .S(_04716_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13572_ (.I0(\samples_imag[1][6] ),
    .I1(_04655_),
    .S(_04700_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13573_ (.I0(_04654_),
    .I1(_04731_),
    .S(_04722_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13574_ (.I0(net60),
    .I1(_04732_),
    .S(_04719_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13575_ (.I0(\samples_imag[1][6] ),
    .I1(_04733_),
    .S(_04716_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13576_ (.I(_04021_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13577_ (.I0(\samples_imag[1][7] ),
    .I1(_04662_),
    .S(_04734_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13578_ (.I0(_04661_),
    .I1(_04735_),
    .S(_04722_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13579_ (.I0(net61),
    .I1(_04736_),
    .S(_04719_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13580_ (.I0(\samples_imag[1][7] ),
    .I1(_04737_),
    .S(_04716_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13581_ (.I0(\samples_imag[1][8] ),
    .I1(_04669_),
    .S(_04734_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13582_ (.I0(_04668_),
    .I1(_04738_),
    .S(_04722_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13583_ (.I0(net62),
    .I1(_04739_),
    .S(_04719_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13584_ (.I0(\samples_imag[1][8] ),
    .I1(_04740_),
    .S(_04716_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13585_ (.I0(\samples_imag[1][9] ),
    .I1(_04676_),
    .S(_04734_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13586_ (.I0(_04675_),
    .I1(_04741_),
    .S(_04722_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13587_ (.I0(net63),
    .I1(_04742_),
    .S(_04719_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13588_ (.I0(\samples_imag[1][9] ),
    .I1(_04743_),
    .S(_04716_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13589_ (.I(\bit_rev_idx[1] ),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13590_ (.A1(_04744_),
    .A2(\bit_rev_idx[0] ),
    .A3(\bit_rev_idx[2] ),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13591_ (.A1(_04516_),
    .A2(_04745_),
    .B(_04683_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13592_ (.A1(_04511_),
    .A2(_04746_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13593_ (.I0(\samples_imag[2][0] ),
    .I1(_04747_),
    .S(_04189_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13594_ (.A1(_07817_),
    .A2(_04551_),
    .A3(_04746_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13595_ (.I0(_04748_),
    .I1(_04749_),
    .S(_03762_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13596_ (.A1(_03596_),
    .A2(_04750_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13597_ (.I0(\samples_imag[2][0] ),
    .I1(_04556_),
    .S(_04746_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13598_ (.A1(_04751_),
    .A2(_04752_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13599_ (.I0(\samples_imag[2][10] ),
    .I1(_04573_),
    .S(_04189_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13600_ (.A1(_03673_),
    .A2(_03696_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13601_ (.I(_04754_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13602_ (.I0(_04571_),
    .I1(_04753_),
    .S(_04755_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13603_ (.I0(net49),
    .I1(_04756_),
    .S(_04719_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13604_ (.I(_04746_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13605_ (.I0(\samples_imag[2][10] ),
    .I1(_04757_),
    .S(_04758_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13606_ (.I0(\samples_imag[2][11] ),
    .I1(_04585_),
    .S(_04189_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13607_ (.I0(_04584_),
    .I1(_04759_),
    .S(_04755_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13608_ (.I0(net50),
    .I1(_04760_),
    .S(_04719_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13609_ (.I0(\samples_imag[2][11] ),
    .I1(_04761_),
    .S(_04758_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13610_ (.I0(\samples_imag[2][12] ),
    .I1(_04595_),
    .S(_04189_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13611_ (.I0(_04594_),
    .I1(_04762_),
    .S(_04755_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13612_ (.I(_04577_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13613_ (.I0(net51),
    .I1(_04763_),
    .S(_04764_),
    .Z(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13614_ (.I0(\samples_imag[2][12] ),
    .I1(_04765_),
    .S(_04758_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13615_ (.I0(\samples_imag[2][13] ),
    .I1(_04602_),
    .S(_04189_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13616_ (.I0(_04601_),
    .I1(_04766_),
    .S(_04755_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13617_ (.I0(net52),
    .I1(_04767_),
    .S(_04764_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13618_ (.I0(\samples_imag[2][13] ),
    .I1(_04768_),
    .S(_04758_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13619_ (.I0(\samples_imag[2][14] ),
    .I1(_04610_),
    .S(_04189_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13620_ (.I0(_04609_),
    .I1(_04769_),
    .S(_04755_),
    .Z(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13621_ (.I0(net53),
    .I1(_04770_),
    .S(_04764_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13622_ (.I0(\samples_imag[2][14] ),
    .I1(_04771_),
    .S(_04758_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13623_ (.I0(\samples_imag[2][15] ),
    .I1(_04615_),
    .S(_04189_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13624_ (.I0(_04549_),
    .I1(_04772_),
    .S(_04755_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13625_ (.I0(net54),
    .I1(_04773_),
    .S(_04764_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13626_ (.I0(\samples_imag[2][15] ),
    .I1(_04774_),
    .S(_04758_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13627_ (.I0(\samples_imag[2][1] ),
    .I1(_04621_),
    .S(_04189_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13628_ (.I0(_04620_),
    .I1(_04775_),
    .S(_04755_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13629_ (.I0(net55),
    .I1(_04776_),
    .S(_04764_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13630_ (.I0(\samples_imag[2][1] ),
    .I1(_04777_),
    .S(_04758_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13631_ (.I(_04076_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13632_ (.I0(\samples_imag[2][2] ),
    .I1(_04627_),
    .S(_04778_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13633_ (.I0(_04626_),
    .I1(_04779_),
    .S(_04755_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13634_ (.I0(net56),
    .I1(_04780_),
    .S(_04764_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13635_ (.I0(\samples_imag[2][2] ),
    .I1(_04781_),
    .S(_04758_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13636_ (.I0(\samples_imag[2][3] ),
    .I1(_04633_),
    .S(_04778_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13637_ (.I0(_04632_),
    .I1(_04782_),
    .S(_04755_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13638_ (.I0(net57),
    .I1(_04783_),
    .S(_04764_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13639_ (.I0(\samples_imag[2][3] ),
    .I1(_04784_),
    .S(_04758_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13640_ (.I0(\samples_imag[2][4] ),
    .I1(_04640_),
    .S(_04778_),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13641_ (.I0(_04639_),
    .I1(_04785_),
    .S(_04755_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13642_ (.I0(net58),
    .I1(_04786_),
    .S(_04764_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13643_ (.I0(\samples_imag[2][4] ),
    .I1(_04787_),
    .S(_04758_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13644_ (.I0(\samples_imag[2][5] ),
    .I1(_04647_),
    .S(_04778_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13645_ (.I(_04754_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13646_ (.I0(_04646_),
    .I1(_04788_),
    .S(_04789_),
    .Z(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13647_ (.I0(net59),
    .I1(_04790_),
    .S(_04764_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13648_ (.I(_04746_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13649_ (.I0(\samples_imag[2][5] ),
    .I1(_04791_),
    .S(_04792_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13650_ (.I0(\samples_imag[2][6] ),
    .I1(_04655_),
    .S(_04778_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13651_ (.I0(_04654_),
    .I1(_04793_),
    .S(_04789_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13652_ (.I0(net60),
    .I1(_04794_),
    .S(_04764_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13653_ (.I0(\samples_imag[2][6] ),
    .I1(_04795_),
    .S(_04792_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13654_ (.I0(\samples_imag[2][7] ),
    .I1(_04662_),
    .S(_04778_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13655_ (.I0(_04661_),
    .I1(_04796_),
    .S(_04789_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13656_ (.I(_04577_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13657_ (.I0(net61),
    .I1(_04797_),
    .S(_04798_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13658_ (.I0(\samples_imag[2][7] ),
    .I1(_04799_),
    .S(_04792_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13659_ (.I0(\samples_imag[2][8] ),
    .I1(_04669_),
    .S(_04778_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13660_ (.I0(_04668_),
    .I1(_04800_),
    .S(_04789_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13661_ (.I0(net62),
    .I1(_04801_),
    .S(_04798_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13662_ (.I0(\samples_imag[2][8] ),
    .I1(_04802_),
    .S(_04792_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13663_ (.I0(\samples_imag[2][9] ),
    .I1(_04676_),
    .S(_04778_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13664_ (.I0(_04675_),
    .I1(_04803_),
    .S(_04789_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13665_ (.I0(net63),
    .I1(_04804_),
    .S(_04798_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13666_ (.I0(\samples_imag[2][9] ),
    .I1(_04805_),
    .S(_04792_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13667_ (.A1(\bit_rev_idx[1] ),
    .A2(\bit_rev_idx[0] ),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13668_ (.A1(\bit_rev_idx[2] ),
    .A2(_04806_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13669_ (.A1(_04516_),
    .A2(_04807_),
    .B(_04683_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13670_ (.A1(_04511_),
    .A2(_04808_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13671_ (.I0(\samples_imag[3][0] ),
    .I1(_04809_),
    .S(_04157_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13672_ (.A1(_07817_),
    .A2(_04551_),
    .A3(_04808_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13673_ (.I0(_04810_),
    .I1(_04811_),
    .S(_03806_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13674_ (.A1(_03596_),
    .A2(_04812_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13675_ (.I0(\samples_imag[3][0] ),
    .I1(_04556_),
    .S(_04808_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13676_ (.A1(_04813_),
    .A2(_04814_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13677_ (.I0(\samples_imag[3][10] ),
    .I1(_04573_),
    .S(_04157_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13678_ (.A1(_03731_),
    .A2(_03804_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13679_ (.I(_04816_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13680_ (.I0(_04571_),
    .I1(_04815_),
    .S(_04817_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13681_ (.I0(net49),
    .I1(_04818_),
    .S(_04798_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13682_ (.I(_04808_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13683_ (.I0(\samples_imag[3][10] ),
    .I1(_04819_),
    .S(_04820_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13684_ (.I0(\samples_imag[3][11] ),
    .I1(_04585_),
    .S(_04157_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13685_ (.I0(_04584_),
    .I1(_04821_),
    .S(_04817_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13686_ (.I0(net50),
    .I1(_04822_),
    .S(_04798_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13687_ (.I0(\samples_imag[3][11] ),
    .I1(_04823_),
    .S(_04820_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13688_ (.I0(\samples_imag[3][12] ),
    .I1(_04595_),
    .S(_04157_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13689_ (.I0(_04594_),
    .I1(_04824_),
    .S(_04817_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13690_ (.I0(net51),
    .I1(_04825_),
    .S(_04798_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13691_ (.I0(\samples_imag[3][12] ),
    .I1(_04826_),
    .S(_04820_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13692_ (.I0(\samples_imag[3][13] ),
    .I1(_04602_),
    .S(_04157_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13693_ (.I0(_04601_),
    .I1(_04827_),
    .S(_04817_),
    .Z(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13694_ (.I0(net52),
    .I1(_04828_),
    .S(_04798_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13695_ (.I0(\samples_imag[3][13] ),
    .I1(_04829_),
    .S(_04820_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13696_ (.I0(\samples_imag[3][14] ),
    .I1(_04610_),
    .S(_04157_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13697_ (.I0(_04609_),
    .I1(_04830_),
    .S(_04817_),
    .Z(_04831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13698_ (.I0(net53),
    .I1(_04831_),
    .S(_04798_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13699_ (.I0(\samples_imag[3][14] ),
    .I1(_04832_),
    .S(_04820_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13700_ (.I0(\samples_imag[3][15] ),
    .I1(_04615_),
    .S(_04157_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13701_ (.I0(_04549_),
    .I1(_04833_),
    .S(_04817_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13702_ (.I0(net54),
    .I1(_04834_),
    .S(_04798_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13703_ (.I0(\samples_imag[3][15] ),
    .I1(_04835_),
    .S(_04820_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13704_ (.I(_04017_),
    .Z(_04836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13705_ (.I0(\samples_imag[3][1] ),
    .I1(_04621_),
    .S(_04836_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13706_ (.I0(_04620_),
    .I1(_04837_),
    .S(_04817_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13707_ (.I0(net55),
    .I1(_04838_),
    .S(_04798_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13708_ (.I0(\samples_imag[3][1] ),
    .I1(_04839_),
    .S(_04820_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13709_ (.I0(\samples_imag[3][2] ),
    .I1(_04627_),
    .S(_04836_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13710_ (.I0(_04626_),
    .I1(_04840_),
    .S(_04817_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13711_ (.I(_04577_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13712_ (.I0(net56),
    .I1(_04841_),
    .S(_04842_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13713_ (.I0(\samples_imag[3][2] ),
    .I1(_04843_),
    .S(_04820_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13714_ (.I0(\samples_imag[3][3] ),
    .I1(_04633_),
    .S(_04836_),
    .Z(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13715_ (.I0(_04632_),
    .I1(_04844_),
    .S(_04817_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13716_ (.I0(net57),
    .I1(_04845_),
    .S(_04842_),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13717_ (.I0(\samples_imag[3][3] ),
    .I1(_04846_),
    .S(_04820_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13718_ (.I0(\samples_imag[3][4] ),
    .I1(_04640_),
    .S(_04836_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13719_ (.I0(_04639_),
    .I1(_04847_),
    .S(_04817_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13720_ (.I0(net58),
    .I1(_04848_),
    .S(_04842_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13721_ (.I0(\samples_imag[3][4] ),
    .I1(_04849_),
    .S(_04820_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13722_ (.I0(\samples_imag[3][5] ),
    .I1(_04647_),
    .S(_04836_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13723_ (.I(_04816_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13724_ (.I0(_04646_),
    .I1(_04850_),
    .S(_04851_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13725_ (.I0(net59),
    .I1(_04852_),
    .S(_04842_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13726_ (.I(_04808_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13727_ (.I0(\samples_imag[3][5] ),
    .I1(_04853_),
    .S(_04854_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13728_ (.I0(\samples_imag[3][6] ),
    .I1(_04655_),
    .S(_04836_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13729_ (.I0(_04654_),
    .I1(_04855_),
    .S(_04851_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13730_ (.I0(net60),
    .I1(_04856_),
    .S(_04842_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13731_ (.I0(\samples_imag[3][6] ),
    .I1(_04857_),
    .S(_04854_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13732_ (.I0(\samples_imag[3][7] ),
    .I1(_04662_),
    .S(_04836_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13733_ (.I0(_04661_),
    .I1(_04858_),
    .S(_04851_),
    .Z(_04859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13734_ (.I0(net61),
    .I1(_04859_),
    .S(_04842_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13735_ (.I0(\samples_imag[3][7] ),
    .I1(_04860_),
    .S(_04854_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13736_ (.I0(\samples_imag[3][8] ),
    .I1(_04669_),
    .S(_04836_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13737_ (.I0(_04668_),
    .I1(_04861_),
    .S(_04851_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13738_ (.I0(net62),
    .I1(_04862_),
    .S(_04842_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13739_ (.I0(\samples_imag[3][8] ),
    .I1(_04863_),
    .S(_04854_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13740_ (.I0(\samples_imag[3][9] ),
    .I1(_04676_),
    .S(_04836_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13741_ (.I0(_04675_),
    .I1(_04864_),
    .S(_04851_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13742_ (.I0(net63),
    .I1(_04865_),
    .S(_04842_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13743_ (.I0(\samples_imag[3][9] ),
    .I1(_04866_),
    .S(_04854_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13744_ (.I(\bit_rev_idx[2] ),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13745_ (.A1(\bit_rev_idx[1] ),
    .A2(\bit_rev_idx[0] ),
    .A3(_04867_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13746_ (.A1(_04516_),
    .A2(_04868_),
    .B(_04683_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13747_ (.A1(_04511_),
    .A2(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13748_ (.I0(\samples_imag[4][0] ),
    .I1(_04870_),
    .S(_04155_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13749_ (.A1(_07817_),
    .A2(_04551_),
    .A3(_04869_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13750_ (.I0(_04871_),
    .I1(_04872_),
    .S(_03760_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13751_ (.A1(_03596_),
    .A2(_04873_),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13752_ (.I0(\samples_imag[4][0] ),
    .I1(_04556_),
    .S(_04869_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13753_ (.A1(_04874_),
    .A2(_04875_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13754_ (.I0(\samples_imag[4][10] ),
    .I1(_04573_),
    .S(_04155_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13755_ (.A1(_03737_),
    .A2(_03758_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13756_ (.I(_04877_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13757_ (.I0(_04571_),
    .I1(_04876_),
    .S(_04878_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13758_ (.I0(net49),
    .I1(_04879_),
    .S(_04842_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13759_ (.I(_04869_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13760_ (.I0(\samples_imag[4][10] ),
    .I1(_04880_),
    .S(_04881_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13761_ (.I0(\samples_imag[4][11] ),
    .I1(_04585_),
    .S(_04155_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13762_ (.I0(_04584_),
    .I1(_04882_),
    .S(_04878_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13763_ (.I0(net50),
    .I1(_04883_),
    .S(_04842_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13764_ (.I0(\samples_imag[4][11] ),
    .I1(_04884_),
    .S(_04881_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13765_ (.I0(\samples_imag[4][12] ),
    .I1(_04595_),
    .S(_04155_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13766_ (.I0(_04594_),
    .I1(_04885_),
    .S(_04878_),
    .Z(_04886_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13767_ (.I(_04577_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13768_ (.I0(net51),
    .I1(_04886_),
    .S(_04887_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13769_ (.I0(\samples_imag[4][12] ),
    .I1(_04888_),
    .S(_04881_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13770_ (.I0(\samples_imag[4][13] ),
    .I1(_04602_),
    .S(_04155_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13771_ (.I0(_04601_),
    .I1(_04889_),
    .S(_04878_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13772_ (.I0(net52),
    .I1(_04890_),
    .S(_04887_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13773_ (.I0(\samples_imag[4][13] ),
    .I1(_04891_),
    .S(_04881_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13774_ (.I0(\samples_imag[4][14] ),
    .I1(_04610_),
    .S(_04155_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13775_ (.I0(_04609_),
    .I1(_04892_),
    .S(_04878_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13776_ (.I0(net53),
    .I1(_04893_),
    .S(_04887_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13777_ (.I0(\samples_imag[4][14] ),
    .I1(_04894_),
    .S(_04881_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13778_ (.I0(\samples_imag[4][15] ),
    .I1(_04615_),
    .S(_04155_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13779_ (.I0(_04549_),
    .I1(_04895_),
    .S(_04878_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13780_ (.I0(net54),
    .I1(_04896_),
    .S(_04887_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13781_ (.I0(\samples_imag[4][15] ),
    .I1(_04897_),
    .S(_04881_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13782_ (.I0(\samples_imag[4][1] ),
    .I1(_04621_),
    .S(_04155_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13783_ (.I0(_04620_),
    .I1(_04898_),
    .S(_04878_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13784_ (.I0(net55),
    .I1(_04899_),
    .S(_04887_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13785_ (.I0(\samples_imag[4][1] ),
    .I1(_04900_),
    .S(_04881_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13786_ (.I(_04079_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13787_ (.I0(\samples_imag[4][2] ),
    .I1(_04627_),
    .S(_04901_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13788_ (.I0(_04626_),
    .I1(_04902_),
    .S(_04878_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13789_ (.I0(net56),
    .I1(_04903_),
    .S(_04887_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13790_ (.I0(\samples_imag[4][2] ),
    .I1(_04904_),
    .S(_04881_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13791_ (.I0(\samples_imag[4][3] ),
    .I1(_04633_),
    .S(_04901_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13792_ (.I0(_04632_),
    .I1(_04905_),
    .S(_04878_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13793_ (.I0(net57),
    .I1(_04906_),
    .S(_04887_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13794_ (.I0(\samples_imag[4][3] ),
    .I1(_04907_),
    .S(_04881_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13795_ (.I0(\samples_imag[4][4] ),
    .I1(_04640_),
    .S(_04901_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13796_ (.I0(_04639_),
    .I1(_04908_),
    .S(_04878_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13797_ (.I0(net58),
    .I1(_04909_),
    .S(_04887_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13798_ (.I0(\samples_imag[4][4] ),
    .I1(_04910_),
    .S(_04881_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13799_ (.I0(\samples_imag[4][5] ),
    .I1(_04647_),
    .S(_04901_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13800_ (.I(_04877_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13801_ (.I0(_04646_),
    .I1(_04911_),
    .S(_04912_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13802_ (.I0(net59),
    .I1(_04913_),
    .S(_04887_),
    .Z(_04914_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13803_ (.I(_04869_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13804_ (.I0(\samples_imag[4][5] ),
    .I1(_04914_),
    .S(_04915_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13805_ (.I0(\samples_imag[4][6] ),
    .I1(_04655_),
    .S(_04901_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13806_ (.I0(_04654_),
    .I1(_04916_),
    .S(_04912_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13807_ (.I0(net60),
    .I1(_04917_),
    .S(_04887_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13808_ (.I0(\samples_imag[4][6] ),
    .I1(_04918_),
    .S(_04915_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13809_ (.I0(\samples_imag[4][7] ),
    .I1(_04662_),
    .S(_04901_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13810_ (.I0(_04661_),
    .I1(_04919_),
    .S(_04912_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13811_ (.I(_03594_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13812_ (.I(_04921_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13813_ (.I0(net61),
    .I1(_04920_),
    .S(_04922_),
    .Z(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13814_ (.I0(\samples_imag[4][7] ),
    .I1(_04923_),
    .S(_04915_),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13815_ (.I0(\samples_imag[4][8] ),
    .I1(_04669_),
    .S(_04901_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13816_ (.I0(_04668_),
    .I1(_04924_),
    .S(_04912_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13817_ (.I0(net62),
    .I1(_04925_),
    .S(_04922_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13818_ (.I0(\samples_imag[4][8] ),
    .I1(_04926_),
    .S(_04915_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13819_ (.I0(\samples_imag[4][9] ),
    .I1(_04676_),
    .S(_04901_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13820_ (.I0(_04675_),
    .I1(_04927_),
    .S(_04912_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13821_ (.I0(net63),
    .I1(_04928_),
    .S(_04922_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13822_ (.I0(\samples_imag[4][9] ),
    .I1(_04929_),
    .S(_04915_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13823_ (.A1(\bit_rev_idx[1] ),
    .A2(_04680_),
    .A3(_04867_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13824_ (.A1(_04516_),
    .A2(_04930_),
    .B(_04683_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13825_ (.A1(_04511_),
    .A2(_04931_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13826_ (.I0(\samples_imag[5][0] ),
    .I1(_04932_),
    .S(_04158_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13827_ (.A1(_07817_),
    .A2(_04551_),
    .A3(_04931_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13828_ (.I0(_04933_),
    .I1(_04934_),
    .S(_03820_),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13829_ (.A1(_03596_),
    .A2(_04935_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13830_ (.I0(\samples_imag[5][0] ),
    .I1(_04556_),
    .S(_04931_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13831_ (.A1(_04936_),
    .A2(_04937_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13832_ (.I0(\samples_imag[5][10] ),
    .I1(_04573_),
    .S(_04158_),
    .Z(_04938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13833_ (.A1(_03737_),
    .A2(_03767_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13834_ (.I(_04939_),
    .Z(_04940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13835_ (.I0(_04571_),
    .I1(_04938_),
    .S(_04940_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13836_ (.I0(net49),
    .I1(_04941_),
    .S(_04922_),
    .Z(_04942_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13837_ (.I(_04931_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13838_ (.I0(\samples_imag[5][10] ),
    .I1(_04942_),
    .S(_04943_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13839_ (.I0(\samples_imag[5][11] ),
    .I1(_04585_),
    .S(_04158_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13840_ (.I0(_04584_),
    .I1(_04944_),
    .S(_04940_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13841_ (.I0(net50),
    .I1(_04945_),
    .S(_04922_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13842_ (.I0(\samples_imag[5][11] ),
    .I1(_04946_),
    .S(_04943_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13843_ (.I0(\samples_imag[5][12] ),
    .I1(_04595_),
    .S(_04158_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13844_ (.I0(_04594_),
    .I1(_04947_),
    .S(_04940_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13845_ (.I0(net51),
    .I1(_04948_),
    .S(_04922_),
    .Z(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13846_ (.I0(\samples_imag[5][12] ),
    .I1(_04949_),
    .S(_04943_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13847_ (.I0(\samples_imag[5][13] ),
    .I1(_04602_),
    .S(_04158_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13848_ (.I0(_04601_),
    .I1(_04950_),
    .S(_04940_),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13849_ (.I0(net52),
    .I1(_04951_),
    .S(_04922_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13850_ (.I0(\samples_imag[5][13] ),
    .I1(_04952_),
    .S(_04943_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13851_ (.I0(\samples_imag[5][14] ),
    .I1(_04610_),
    .S(_04158_),
    .Z(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13852_ (.I0(_04609_),
    .I1(_04953_),
    .S(_04940_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13853_ (.I0(net53),
    .I1(_04954_),
    .S(_04922_),
    .Z(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13854_ (.I0(\samples_imag[5][14] ),
    .I1(_04955_),
    .S(_04943_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13855_ (.I0(\samples_imag[5][15] ),
    .I1(_04615_),
    .S(_04158_),
    .Z(_04956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13856_ (.I0(_04549_),
    .I1(_04956_),
    .S(_04940_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13857_ (.I0(net54),
    .I1(_04957_),
    .S(_04922_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13858_ (.I0(\samples_imag[5][15] ),
    .I1(_04958_),
    .S(_04943_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13859_ (.I(_04020_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13860_ (.I0(\samples_imag[5][1] ),
    .I1(_04621_),
    .S(_04959_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13861_ (.I0(_04620_),
    .I1(_04960_),
    .S(_04940_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13862_ (.I0(net55),
    .I1(_04961_),
    .S(_04922_),
    .Z(_04962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13863_ (.I0(\samples_imag[5][1] ),
    .I1(_04962_),
    .S(_04943_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13864_ (.I0(\samples_imag[5][2] ),
    .I1(_04627_),
    .S(_04959_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13865_ (.I0(_04626_),
    .I1(_04963_),
    .S(_04940_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13866_ (.I(_04921_),
    .Z(_04965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13867_ (.I0(net56),
    .I1(_04964_),
    .S(_04965_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13868_ (.I0(\samples_imag[5][2] ),
    .I1(_04966_),
    .S(_04943_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13869_ (.I0(\samples_imag[5][3] ),
    .I1(_04633_),
    .S(_04959_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13870_ (.I0(_04632_),
    .I1(_04967_),
    .S(_04940_),
    .Z(_04968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13871_ (.I0(net57),
    .I1(_04968_),
    .S(_04965_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13872_ (.I0(\samples_imag[5][3] ),
    .I1(_04969_),
    .S(_04943_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13873_ (.I0(\samples_imag[5][4] ),
    .I1(_04640_),
    .S(_04959_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13874_ (.I0(_04639_),
    .I1(_04970_),
    .S(_04940_),
    .Z(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13875_ (.I0(net58),
    .I1(_04971_),
    .S(_04965_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13876_ (.I0(\samples_imag[5][4] ),
    .I1(_04972_),
    .S(_04943_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13877_ (.I0(\samples_imag[5][5] ),
    .I1(_04647_),
    .S(_04959_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13878_ (.I(_04939_),
    .Z(_04974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13879_ (.I0(_04646_),
    .I1(_04973_),
    .S(_04974_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13880_ (.I0(net59),
    .I1(_04975_),
    .S(_04965_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13881_ (.I(_04931_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13882_ (.I0(\samples_imag[5][5] ),
    .I1(_04976_),
    .S(_04977_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13883_ (.I0(\samples_imag[5][6] ),
    .I1(_04655_),
    .S(_04959_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13884_ (.I0(_04654_),
    .I1(_04978_),
    .S(_04974_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13885_ (.I0(net60),
    .I1(_04979_),
    .S(_04965_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13886_ (.I0(\samples_imag[5][6] ),
    .I1(_04980_),
    .S(_04977_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13887_ (.I0(\samples_imag[5][7] ),
    .I1(_04662_),
    .S(_04959_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13888_ (.I0(_04661_),
    .I1(_04981_),
    .S(_04974_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13889_ (.I0(net61),
    .I1(_04982_),
    .S(_04965_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13890_ (.I0(\samples_imag[5][7] ),
    .I1(_04983_),
    .S(_04977_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13891_ (.I0(\samples_imag[5][8] ),
    .I1(_04669_),
    .S(_04959_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13892_ (.I0(_04668_),
    .I1(_04984_),
    .S(_04974_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13893_ (.I0(net62),
    .I1(_04985_),
    .S(_04965_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13894_ (.I0(\samples_imag[5][8] ),
    .I1(_04986_),
    .S(_04977_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13895_ (.I0(\samples_imag[5][9] ),
    .I1(_04676_),
    .S(_04959_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13896_ (.I0(_04675_),
    .I1(_04987_),
    .S(_04974_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13897_ (.I0(net63),
    .I1(_04988_),
    .S(_04965_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13898_ (.I0(\samples_imag[5][9] ),
    .I1(_04989_),
    .S(_04977_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13899_ (.A1(_04744_),
    .A2(\bit_rev_idx[0] ),
    .A3(_04867_),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13900_ (.A1(_04516_),
    .A2(_04990_),
    .B(_04683_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13901_ (.A1(_07817_),
    .A2(_04551_),
    .A3(_04991_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13902_ (.A1(_04511_),
    .A2(_04991_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13903_ (.I0(\samples_imag[6][0] ),
    .I1(_04993_),
    .S(_04041_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13904_ (.A1(_03685_),
    .A2(_03707_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13905_ (.I(_04995_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13906_ (.I0(_04992_),
    .I1(_04994_),
    .S(_04996_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13907_ (.A1(_03596_),
    .A2(_04997_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13908_ (.I0(\samples_imag[6][0] ),
    .I1(_04556_),
    .S(_04991_),
    .Z(_04999_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13909_ (.A1(_04998_),
    .A2(_04999_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13910_ (.I0(\samples_imag[6][10] ),
    .I1(_04573_),
    .S(_04041_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13911_ (.I0(_04571_),
    .I1(_05000_),
    .S(_04996_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13912_ (.I0(net49),
    .I1(_05001_),
    .S(_04965_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13913_ (.I(_04991_),
    .Z(_05003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13914_ (.I0(\samples_imag[6][10] ),
    .I1(_05002_),
    .S(_05003_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13915_ (.I0(\samples_imag[6][11] ),
    .I1(_04585_),
    .S(_04041_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13916_ (.I0(_04584_),
    .I1(_05004_),
    .S(_04996_),
    .Z(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13917_ (.I0(net50),
    .I1(_05005_),
    .S(_04965_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13918_ (.I0(\samples_imag[6][11] ),
    .I1(_05006_),
    .S(_05003_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13919_ (.I0(\samples_imag[6][12] ),
    .I1(_04595_),
    .S(_04041_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13920_ (.I0(_04594_),
    .I1(_05007_),
    .S(_04996_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13921_ (.I(_04921_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13922_ (.I0(net51),
    .I1(_05008_),
    .S(_05009_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13923_ (.I0(\samples_imag[6][12] ),
    .I1(_05010_),
    .S(_05003_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13924_ (.I0(\samples_imag[6][13] ),
    .I1(_04602_),
    .S(_04041_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13925_ (.I0(_04601_),
    .I1(_05011_),
    .S(_04996_),
    .Z(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13926_ (.I0(net52),
    .I1(_05012_),
    .S(_05009_),
    .Z(_05013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13927_ (.I0(\samples_imag[6][13] ),
    .I1(_05013_),
    .S(_05003_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13928_ (.I0(\samples_imag[6][14] ),
    .I1(_04610_),
    .S(_04041_),
    .Z(_05014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13929_ (.I0(_04609_),
    .I1(_05014_),
    .S(_04996_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13930_ (.I0(net53),
    .I1(_05015_),
    .S(_05009_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13931_ (.I0(\samples_imag[6][14] ),
    .I1(_05016_),
    .S(_05003_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13932_ (.I0(\samples_imag[6][15] ),
    .I1(_04615_),
    .S(_04041_),
    .Z(_05017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13933_ (.I0(_04549_),
    .I1(_05017_),
    .S(_04996_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13934_ (.I0(net54),
    .I1(_05018_),
    .S(_05009_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13935_ (.I0(\samples_imag[6][15] ),
    .I1(_05019_),
    .S(_05003_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13936_ (.I(_04040_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13937_ (.I0(\samples_imag[6][1] ),
    .I1(_04621_),
    .S(_05020_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13938_ (.I0(_04620_),
    .I1(_05021_),
    .S(_04996_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13939_ (.I0(net55),
    .I1(_05022_),
    .S(_05009_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13940_ (.I0(\samples_imag[6][1] ),
    .I1(_05023_),
    .S(_05003_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13941_ (.I0(\samples_imag[6][2] ),
    .I1(_04627_),
    .S(_05020_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13942_ (.I0(_04626_),
    .I1(_05024_),
    .S(_04996_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13943_ (.I0(net56),
    .I1(_05025_),
    .S(_05009_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13944_ (.I0(\samples_imag[6][2] ),
    .I1(_05026_),
    .S(_05003_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13945_ (.I0(\samples_imag[6][3] ),
    .I1(_04633_),
    .S(_05020_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13946_ (.I(_04995_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13947_ (.I0(_04632_),
    .I1(_05027_),
    .S(_05028_),
    .Z(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13948_ (.I0(net57),
    .I1(_05029_),
    .S(_05009_),
    .Z(_05030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13949_ (.I0(\samples_imag[6][3] ),
    .I1(_05030_),
    .S(_05003_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13950_ (.I0(\samples_imag[6][4] ),
    .I1(_04640_),
    .S(_05020_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13951_ (.I0(_04639_),
    .I1(_05031_),
    .S(_05028_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13952_ (.I0(net58),
    .I1(_05032_),
    .S(_05009_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13953_ (.I0(\samples_imag[6][4] ),
    .I1(_05033_),
    .S(_05003_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13954_ (.I0(\samples_imag[6][5] ),
    .I1(_04647_),
    .S(_05020_),
    .Z(_05034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13955_ (.I0(_04646_),
    .I1(_05034_),
    .S(_05028_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13956_ (.I0(net59),
    .I1(_05035_),
    .S(_05009_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13957_ (.I(_04991_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13958_ (.I0(\samples_imag[6][5] ),
    .I1(_05036_),
    .S(_05037_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13959_ (.I0(\samples_imag[6][6] ),
    .I1(_04655_),
    .S(_05020_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13960_ (.I0(_04654_),
    .I1(_05038_),
    .S(_05028_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13961_ (.I0(net60),
    .I1(_05039_),
    .S(_05009_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13962_ (.I0(\samples_imag[6][6] ),
    .I1(_05040_),
    .S(_05037_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13963_ (.I0(\samples_imag[6][7] ),
    .I1(_04662_),
    .S(_05020_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13964_ (.I0(_04661_),
    .I1(_05041_),
    .S(_05028_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13965_ (.I(_04921_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13966_ (.I0(net61),
    .I1(_05042_),
    .S(_05043_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13967_ (.I0(\samples_imag[6][7] ),
    .I1(_05044_),
    .S(_05037_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13968_ (.I0(\samples_imag[6][8] ),
    .I1(_04669_),
    .S(_05020_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13969_ (.I0(_04668_),
    .I1(_05045_),
    .S(_05028_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13970_ (.I0(net62),
    .I1(_05046_),
    .S(_05043_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13971_ (.I0(\samples_imag[6][8] ),
    .I1(_05047_),
    .S(_05037_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13972_ (.I0(\samples_imag[6][9] ),
    .I1(_04676_),
    .S(_05020_),
    .Z(_05048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13973_ (.I0(_04675_),
    .I1(_05048_),
    .S(_05028_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13974_ (.I0(net63),
    .I1(_05049_),
    .S(_05043_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13975_ (.I0(\samples_imag[6][9] ),
    .I1(_05050_),
    .S(_05037_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13976_ (.A1(_03643_),
    .A2(_04011_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13977_ (.A1(_04867_),
    .A2(_04806_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13978_ (.A1(net80),
    .A2(_05052_),
    .B(_04515_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13979_ (.A1(_04254_),
    .A2(_05053_),
    .B(_04513_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13980_ (.A1(_05051_),
    .A2(_05054_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13981_ (.A1(\samples_imag[7][0] ),
    .A2(_05051_),
    .B1(_04511_),
    .B2(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13982_ (.A1(_03729_),
    .A2(_03707_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13983_ (.I(_05057_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13984_ (.A1(_05058_),
    .A2(_05054_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _13985_ (.A1(_03753_),
    .A2(_05056_),
    .B1(_05059_),
    .B2(_04552_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13986_ (.A1(_03596_),
    .A2(_05060_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13987_ (.I0(_04556_),
    .I1(\samples_imag[7][0] ),
    .S(_05054_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13988_ (.A1(_05061_),
    .A2(_05062_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13989_ (.I0(\samples_imag[7][10] ),
    .I1(_04573_),
    .S(_04164_),
    .Z(_05063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13990_ (.I0(_04571_),
    .I1(_05063_),
    .S(_05058_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _13991_ (.I(_03594_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13992_ (.I0(net49),
    .I1(_05064_),
    .S(_05065_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _13993_ (.I(_05054_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13994_ (.I0(_05066_),
    .I1(\samples_imag[7][10] ),
    .S(_05067_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13995_ (.I0(\samples_imag[7][11] ),
    .I1(_04585_),
    .S(_04164_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13996_ (.I0(_04584_),
    .I1(_05068_),
    .S(_05058_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13997_ (.I0(net50),
    .I1(_05069_),
    .S(_05065_),
    .Z(_05070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13998_ (.I0(_05070_),
    .I1(\samples_imag[7][11] ),
    .S(_05067_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13999_ (.I0(\samples_imag[7][12] ),
    .I1(_04595_),
    .S(_04164_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14000_ (.I0(_04594_),
    .I1(_05071_),
    .S(_05058_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14001_ (.I(_04577_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14002_ (.I0(net51),
    .I1(_05072_),
    .S(_05073_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14003_ (.I0(_05074_),
    .I1(\samples_imag[7][12] ),
    .S(_05067_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14004_ (.I0(\samples_imag[7][13] ),
    .I1(_04602_),
    .S(_04164_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14005_ (.I0(_04601_),
    .I1(_05075_),
    .S(_05058_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14006_ (.I0(net52),
    .I1(_05076_),
    .S(_05073_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14007_ (.I0(_05077_),
    .I1(\samples_imag[7][13] ),
    .S(_05067_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14008_ (.I0(\samples_imag[7][14] ),
    .I1(_04610_),
    .S(_04164_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14009_ (.I0(_04609_),
    .I1(_05078_),
    .S(_05058_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14010_ (.I0(net53),
    .I1(_05079_),
    .S(_05073_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14011_ (.I0(_05080_),
    .I1(\samples_imag[7][14] ),
    .S(_05067_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14012_ (.I0(\samples_imag[7][15] ),
    .I1(_04615_),
    .S(_04164_),
    .Z(_05081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14013_ (.I0(_04549_),
    .I1(_05081_),
    .S(_05058_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14014_ (.I0(net54),
    .I1(_05082_),
    .S(_05073_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14015_ (.I0(_05083_),
    .I1(\samples_imag[7][15] ),
    .S(_05067_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14016_ (.I0(\samples_imag[7][1] ),
    .I1(_04621_),
    .S(_04164_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14017_ (.I0(_04620_),
    .I1(_05084_),
    .S(_05058_),
    .Z(_05085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14018_ (.I0(net55),
    .I1(_05085_),
    .S(_05073_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14019_ (.I0(_05086_),
    .I1(\samples_imag[7][1] ),
    .S(_05067_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14020_ (.I0(\samples_imag[7][2] ),
    .I1(_04627_),
    .S(_04164_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14021_ (.I0(_04626_),
    .I1(_05087_),
    .S(_05058_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14022_ (.I0(net56),
    .I1(_05088_),
    .S(_05073_),
    .Z(_05089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14023_ (.I0(_05089_),
    .I1(\samples_imag[7][2] ),
    .S(_05067_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14024_ (.I0(\samples_imag[7][3] ),
    .I1(_04633_),
    .S(_04164_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14025_ (.I0(_04632_),
    .I1(_05090_),
    .S(_05058_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14026_ (.I0(net57),
    .I1(_05091_),
    .S(_05073_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14027_ (.I0(_05092_),
    .I1(\samples_imag[7][3] ),
    .S(_05067_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14028_ (.I(_04013_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14029_ (.I0(\samples_imag[7][4] ),
    .I1(_04640_),
    .S(_05093_),
    .Z(_05094_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14030_ (.I(_05057_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14031_ (.I0(_04639_),
    .I1(_05094_),
    .S(_05095_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14032_ (.I0(net58),
    .I1(_05096_),
    .S(_05073_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14033_ (.I0(_05097_),
    .I1(\samples_imag[7][4] ),
    .S(_05067_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14034_ (.I0(\samples_imag[7][5] ),
    .I1(_04647_),
    .S(_05093_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14035_ (.I0(_04646_),
    .I1(_05098_),
    .S(_05095_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14036_ (.I0(net59),
    .I1(_05099_),
    .S(_05073_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14037_ (.I(_05054_),
    .Z(_05101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14038_ (.I0(_05100_),
    .I1(\samples_imag[7][5] ),
    .S(_05101_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14039_ (.I0(\samples_imag[7][6] ),
    .I1(_04655_),
    .S(_05093_),
    .Z(_05102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14040_ (.I0(_04654_),
    .I1(_05102_),
    .S(_05095_),
    .Z(_05103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14041_ (.I0(net60),
    .I1(_05103_),
    .S(_05073_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14042_ (.I0(_05104_),
    .I1(\samples_imag[7][6] ),
    .S(_05101_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14043_ (.I0(\samples_imag[7][7] ),
    .I1(_04662_),
    .S(_05093_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14044_ (.I0(_04661_),
    .I1(_05105_),
    .S(_05095_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14045_ (.I(_04577_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14046_ (.I0(net61),
    .I1(_05106_),
    .S(_05107_),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14047_ (.I0(_05108_),
    .I1(\samples_imag[7][7] ),
    .S(_05101_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14048_ (.I0(\samples_imag[7][8] ),
    .I1(_04669_),
    .S(_05093_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14049_ (.I0(_04668_),
    .I1(_05109_),
    .S(_05095_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14050_ (.I0(net62),
    .I1(_05110_),
    .S(_05107_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14051_ (.I0(_05111_),
    .I1(\samples_imag[7][8] ),
    .S(_05101_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14052_ (.I0(\samples_imag[7][9] ),
    .I1(_04676_),
    .S(_05093_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14053_ (.I0(_04675_),
    .I1(_05112_),
    .S(_05095_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14054_ (.I0(net63),
    .I1(_05113_),
    .S(_05107_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14055_ (.I0(_05114_),
    .I1(\samples_imag[7][9] ),
    .S(_05101_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14056_ (.I(_07703_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14057_ (.A1(\temp_real[0] ),
    .A2(_04037_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14058_ (.I(_07698_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14059_ (.I(_07717_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14060_ (.I(_07727_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14061_ (.I(_07737_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14062_ (.I(_07747_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14063_ (.I(_07757_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14064_ (.I(_07766_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14065_ (.A1(_05123_),
    .A2(_07701_),
    .B(_07767_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14066_ (.I(_07763_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14067_ (.A1(_07762_),
    .A2(_05124_),
    .B(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14068_ (.A1(_05122_),
    .A2(_05126_),
    .B(_07758_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14069_ (.I(_07753_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14070_ (.A1(_07752_),
    .A2(_05127_),
    .B(_05128_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14071_ (.A1(_05121_),
    .A2(_05129_),
    .B(_07748_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14072_ (.I(_07743_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14073_ (.A1(_07742_),
    .A2(_05130_),
    .B(_05131_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14074_ (.A1(_05120_),
    .A2(_05132_),
    .B(_07738_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14075_ (.I(_07733_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14076_ (.A1(_07732_),
    .A2(_05133_),
    .B(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14077_ (.A1(_05119_),
    .A2(_05135_),
    .B(_07728_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14078_ (.I(_07723_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14079_ (.A1(_07722_),
    .A2(_05136_),
    .B(_05137_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14080_ (.A1(_05118_),
    .A2(_05138_),
    .B(_07718_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14081_ (.I(_07713_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14082_ (.A1(_07712_),
    .A2(_05139_),
    .B(_05140_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14083_ (.A1(_05117_),
    .A2(_05141_),
    .B(_07699_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14084_ (.I(_07694_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14085_ (.A1(_07693_),
    .A2(_05142_),
    .B(_05143_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14086_ (.A1(_05116_),
    .A2(_05144_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14087_ (.A1(_07762_),
    .A2(_05855_),
    .B(_05125_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14088_ (.A1(_05122_),
    .A2(_05146_),
    .B(_07758_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14089_ (.A1(_07752_),
    .A2(_05147_),
    .B(_05128_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14090_ (.A1(_05121_),
    .A2(_05148_),
    .B(_07748_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14091_ (.A1(_07742_),
    .A2(_05149_),
    .B(_05131_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14092_ (.A1(_05120_),
    .A2(_05150_),
    .B(_07738_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14093_ (.A1(_07732_),
    .A2(_05151_),
    .B(_05134_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14094_ (.A1(_05119_),
    .A2(_05152_),
    .B(_07728_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14095_ (.A1(_07722_),
    .A2(_05153_),
    .B(_05137_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14096_ (.A1(_05118_),
    .A2(_05154_),
    .B(_07718_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14097_ (.A1(_07712_),
    .A2(_05155_),
    .B(_05140_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14098_ (.A1(_05117_),
    .A2(_05156_),
    .B(_07699_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14099_ (.A1(_07693_),
    .A2(_05157_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14100_ (.A1(_05117_),
    .A2(_05141_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14101_ (.A1(_05119_),
    .A2(_05135_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14102_ (.A1(_07712_),
    .A2(_05155_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14103_ (.A1(_05118_),
    .A2(_05138_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14104_ (.A1(_07722_),
    .A2(_05153_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14105_ (.A1(_07742_),
    .A2(_05149_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14106_ (.A1(_05121_),
    .A2(_05129_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14107_ (.A1(_05122_),
    .A2(_05126_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14108_ (.A1(_07762_),
    .A2(_05855_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14109_ (.A1(_07752_),
    .A2(_05147_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14110_ (.A1(_05856_),
    .A2(_05115_),
    .A3(_05167_),
    .A4(_05168_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14111_ (.A1(_05164_),
    .A2(_05165_),
    .A3(_05166_),
    .A4(_05169_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14112_ (.A1(_07732_),
    .A2(_05151_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14113_ (.A1(_05120_),
    .A2(_05132_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14114_ (.A1(_05163_),
    .A2(_05170_),
    .A3(_05171_),
    .A4(_05172_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14115_ (.A1(_05160_),
    .A2(_05161_),
    .A3(_05162_),
    .A4(_05173_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14116_ (.A1(_05158_),
    .A2(_05159_),
    .A3(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14117_ (.A1(\temp_real[0] ),
    .A2(_07708_),
    .A3(_05175_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14118_ (.A1(_05145_),
    .A2(_05176_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14119_ (.A1(_05115_),
    .A2(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14120_ (.A1(\samples_real[0][0] ),
    .A2(_03641_),
    .B1(_04519_),
    .B2(_05178_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14121_ (.I(_07697_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14122_ (.I(_07711_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14123_ (.I(_07721_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14124_ (.I(_07731_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14125_ (.I(_07741_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14126_ (.I(_07751_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14127_ (.I(_07761_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14128_ (.A1(_07766_),
    .A2(_05858_),
    .Z(_05187_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14129_ (.A1(_07765_),
    .A2(_05187_),
    .B(_07762_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14130_ (.A1(_05186_),
    .A2(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14131_ (.A1(_07757_),
    .A2(_05189_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14132_ (.A1(_07756_),
    .A2(_05190_),
    .B(_07752_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14133_ (.A1(_05185_),
    .A2(_05191_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14134_ (.A1(_07747_),
    .A2(_05192_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14135_ (.A1(_07746_),
    .A2(_05193_),
    .B(_07742_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14136_ (.A1(_05184_),
    .A2(_05194_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14137_ (.A1(_07737_),
    .A2(_05195_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14138_ (.A1(_07736_),
    .A2(_05196_),
    .B(_07732_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14139_ (.A1(_05183_),
    .A2(_05197_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14140_ (.A1(_07727_),
    .A2(_05198_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14141_ (.A1(_07726_),
    .A2(_05199_),
    .B(_07722_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14142_ (.A1(_05182_),
    .A2(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14143_ (.A1(_07717_),
    .A2(_05201_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14144_ (.A1(_07716_),
    .A2(_05202_),
    .B(_07712_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14145_ (.A1(_05181_),
    .A2(_05203_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14146_ (.A1(_07698_),
    .A2(_05204_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14147_ (.A1(_05180_),
    .A2(_05205_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14148_ (.A1(_07693_),
    .A2(_05206_),
    .B(_07692_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _14149_ (.A1(_05116_),
    .A2(_05207_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14150_ (.A1(\temp_real[0] ),
    .A2(_07709_),
    .A3(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _14151_ (.I(_05209_),
    .Z(_05210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14152_ (.A1(_07703_),
    .A2(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14153_ (.A1(_03728_),
    .A2(_05179_),
    .B1(_05211_),
    .B2(_04553_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14154_ (.A1(_03596_),
    .A2(_05212_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14155_ (.A1(_04255_),
    .A2(net64),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14156_ (.I0(\samples_real[0][0] ),
    .I1(_05214_),
    .S(_04518_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14157_ (.A1(_05213_),
    .A2(_05215_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14158_ (.A1(_07762_),
    .A2(_05859_),
    .B(_07761_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14159_ (.I(_07756_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14160_ (.A1(_05122_),
    .A2(_05216_),
    .B(_05217_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14161_ (.A1(_07752_),
    .A2(_05218_),
    .B(_07751_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14162_ (.I(_07746_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14163_ (.A1(_05121_),
    .A2(_05219_),
    .B(_05220_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14164_ (.A1(_07742_),
    .A2(_05221_),
    .B(_07741_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14165_ (.I(_07736_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14166_ (.A1(_05120_),
    .A2(_05222_),
    .B(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14167_ (.A1(_07732_),
    .A2(_05224_),
    .B(_07731_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14168_ (.I(_07726_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14169_ (.A1(_05119_),
    .A2(_05225_),
    .B(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14170_ (.A1(_07722_),
    .A2(_05227_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14171_ (.A1(_05210_),
    .A2(_05228_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14172_ (.I(_05177_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14173_ (.A1(_05163_),
    .A2(_05230_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14174_ (.I0(\samples_real[0][10] ),
    .I1(_05231_),
    .S(_04648_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14175_ (.I0(_05229_),
    .I1(_05232_),
    .S(_04635_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14176_ (.I0(net65),
    .I1(_05233_),
    .S(_05043_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14177_ (.I0(\samples_real[0][10] ),
    .I1(_05234_),
    .S(_04652_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14178_ (.A1(_07717_),
    .A2(_05201_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _14179_ (.I(_05209_),
    .Z(_05236_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14180_ (.A1(_07717_),
    .A2(_05201_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14181_ (.A1(_05235_),
    .A2(_05236_),
    .A3(_05237_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14182_ (.A1(_05162_),
    .A2(_05230_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14183_ (.I0(\samples_real[0][11] ),
    .I1(_05239_),
    .S(_04648_),
    .Z(_05240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14184_ (.I0(_05238_),
    .I1(_05240_),
    .S(_04635_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14185_ (.I0(net66),
    .I1(_05241_),
    .S(_05043_),
    .Z(_05242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14186_ (.I0(\samples_real[0][11] ),
    .I1(_05242_),
    .S(_04652_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14187_ (.A1(_07722_),
    .A2(_05227_),
    .B(_07721_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14188_ (.I(_07716_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14189_ (.A1(_05118_),
    .A2(_05243_),
    .B(_05244_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14190_ (.A1(_07712_),
    .A2(_05245_),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14191_ (.A1(_07712_),
    .A2(_05245_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14192_ (.A1(_05236_),
    .A2(_05246_),
    .A3(_05247_),
    .Z(_05248_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14193_ (.A1(_05161_),
    .A2(_05230_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14194_ (.I0(\samples_real[0][12] ),
    .I1(_05249_),
    .S(_04648_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14195_ (.I0(_05248_),
    .I1(_05250_),
    .S(_04635_),
    .Z(_05251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14196_ (.I0(net67),
    .I1(_05251_),
    .S(_05043_),
    .Z(_05252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14197_ (.I0(\samples_real[0][12] ),
    .I1(_05252_),
    .S(_04652_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14198_ (.A1(_07698_),
    .A2(_05204_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14199_ (.A1(_05205_),
    .A2(_05236_),
    .A3(_05253_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14200_ (.A1(_05159_),
    .A2(_05230_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14201_ (.I0(\samples_real[0][13] ),
    .I1(_05255_),
    .S(_04648_),
    .Z(_05256_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14202_ (.I(_03712_),
    .Z(_05257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14203_ (.I0(_05254_),
    .I1(_05256_),
    .S(_05257_),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14204_ (.I0(net68),
    .I1(_05258_),
    .S(_05043_),
    .Z(_05259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14205_ (.I0(\samples_real[0][13] ),
    .I1(_05259_),
    .S(_04652_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14206_ (.A1(_05181_),
    .A2(_05247_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14207_ (.A1(_07698_),
    .A2(_05260_),
    .B(_07697_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14208_ (.A1(_07693_),
    .A2(_05261_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14209_ (.A1(_05210_),
    .A2(_05262_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14210_ (.A1(_05158_),
    .A2(_05230_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14211_ (.I0(\samples_real[0][14] ),
    .I1(_05264_),
    .S(_04648_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14212_ (.I0(_05263_),
    .I1(_05265_),
    .S(_05257_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14213_ (.I0(net69),
    .I1(_05266_),
    .S(_05043_),
    .Z(_05267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14214_ (.I0(\samples_real[0][14] ),
    .I1(_05267_),
    .S(_04652_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14215_ (.I(_05145_),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14216_ (.A1(_05268_),
    .A2(_05176_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14217_ (.I(_04008_),
    .Z(_05270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14218_ (.I0(\samples_real[0][15] ),
    .I1(_05269_),
    .S(_05270_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14219_ (.I0(_05208_),
    .I1(_05271_),
    .S(_05257_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14220_ (.I0(net70),
    .I1(_05272_),
    .S(_05043_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14221_ (.I(_04518_),
    .Z(_05274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14222_ (.I0(\samples_real[0][15] ),
    .I1(_05273_),
    .S(_05274_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14223_ (.I(_05860_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14224_ (.A1(_05275_),
    .A2(_05236_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14225_ (.A1(_05856_),
    .A2(_05230_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14226_ (.I0(\samples_real[0][1] ),
    .I1(_05277_),
    .S(_05270_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14227_ (.I0(_05276_),
    .I1(_05278_),
    .S(_05257_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14228_ (.I0(net71),
    .I1(_05279_),
    .S(_05043_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14229_ (.I0(\samples_real[0][1] ),
    .I1(_05280_),
    .S(_05274_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14230_ (.A1(_07762_),
    .A2(_05859_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14231_ (.A1(_05210_),
    .A2(_05281_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14232_ (.A1(_05167_),
    .A2(_05230_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14233_ (.I0(\samples_real[0][2] ),
    .I1(_05283_),
    .S(_05270_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14234_ (.I0(_05282_),
    .I1(_05284_),
    .S(_05257_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14235_ (.I(_04921_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14236_ (.I0(net72),
    .I1(_05285_),
    .S(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14237_ (.I0(\samples_real[0][2] ),
    .I1(_05287_),
    .S(_05274_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14238_ (.A1(_05122_),
    .A2(_05189_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14239_ (.A1(_05236_),
    .A2(_05288_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14240_ (.A1(_05166_),
    .A2(_05230_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14241_ (.I0(\samples_real[0][3] ),
    .I1(_05290_),
    .S(_05270_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14242_ (.I0(_05289_),
    .I1(_05291_),
    .S(_05257_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14243_ (.I0(net73),
    .I1(_05292_),
    .S(_05286_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14244_ (.I0(\samples_real[0][3] ),
    .I1(_05293_),
    .S(_05274_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14245_ (.A1(_07752_),
    .A2(_05218_),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14246_ (.A1(_05236_),
    .A2(_05294_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14247_ (.A1(_05168_),
    .A2(_05230_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14248_ (.I0(\samples_real[0][4] ),
    .I1(_05296_),
    .S(_05270_),
    .Z(_05297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14249_ (.I0(_05295_),
    .I1(_05297_),
    .S(_05257_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14250_ (.I0(net74),
    .I1(_05298_),
    .S(_05286_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14251_ (.I0(\samples_real[0][4] ),
    .I1(_05299_),
    .S(_05274_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14252_ (.A1(_07747_),
    .A2(_05192_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14253_ (.A1(_07747_),
    .A2(_05192_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14254_ (.A1(_05300_),
    .A2(_05236_),
    .A3(_05301_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14255_ (.A1(_05165_),
    .A2(_05230_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14256_ (.I0(\samples_real[0][5] ),
    .I1(_05303_),
    .S(_05270_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14257_ (.I0(_05302_),
    .I1(_05304_),
    .S(_05257_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14258_ (.I0(net75),
    .I1(_05305_),
    .S(_05286_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14259_ (.I0(\samples_real[0][5] ),
    .I1(_05306_),
    .S(_05274_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14260_ (.A1(_07742_),
    .A2(_05221_),
    .Z(_05307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14261_ (.A1(_05236_),
    .A2(_05307_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14262_ (.A1(_05164_),
    .A2(_05177_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14263_ (.I0(\samples_real[0][6] ),
    .I1(_05309_),
    .S(_05270_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14264_ (.I0(_05308_),
    .I1(_05310_),
    .S(_05257_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14265_ (.I0(net76),
    .I1(_05311_),
    .S(_05286_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14266_ (.I0(\samples_real[0][6] ),
    .I1(_05312_),
    .S(_05274_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14267_ (.A1(_07737_),
    .A2(_05195_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14268_ (.A1(_07737_),
    .A2(_05195_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14269_ (.A1(_05313_),
    .A2(_05236_),
    .A3(_05314_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14270_ (.A1(_05172_),
    .A2(_05177_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14271_ (.I0(\samples_real[0][7] ),
    .I1(_05316_),
    .S(_05270_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14272_ (.I0(_05315_),
    .I1(_05317_),
    .S(_05257_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14273_ (.I0(net77),
    .I1(_05318_),
    .S(_05286_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14274_ (.I0(\samples_real[0][7] ),
    .I1(_05319_),
    .S(_05274_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14275_ (.A1(_07732_),
    .A2(_05224_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14276_ (.A1(_05236_),
    .A2(_05320_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14277_ (.A1(_05171_),
    .A2(_05177_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14278_ (.I0(\samples_real[0][8] ),
    .I1(_05322_),
    .S(_05270_),
    .Z(_05323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14279_ (.I0(_05321_),
    .I1(_05323_),
    .S(_03712_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14280_ (.I0(net78),
    .I1(_05324_),
    .S(_05286_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14281_ (.I0(\samples_real[0][8] ),
    .I1(_05325_),
    .S(_05274_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14282_ (.A1(_07727_),
    .A2(_05198_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14283_ (.A1(_07727_),
    .A2(_05198_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14284_ (.A1(_05326_),
    .A2(_05209_),
    .A3(_05327_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14285_ (.A1(_05160_),
    .A2(_05177_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14286_ (.I0(\samples_real[0][9] ),
    .I1(_05329_),
    .S(_05270_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14287_ (.I0(_05328_),
    .I1(_05330_),
    .S(_03712_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14288_ (.I0(net79),
    .I1(_05331_),
    .S(_05286_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14289_ (.I0(\samples_real[0][9] ),
    .I1(_05332_),
    .S(_05274_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14290_ (.A1(_04685_),
    .A2(_05178_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14291_ (.I0(\samples_real[1][0] ),
    .I1(_05333_),
    .S(_04094_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14292_ (.A1(_07703_),
    .A2(_03755_),
    .A3(_04685_),
    .A4(_05210_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14293_ (.A1(_04688_),
    .A2(_05334_),
    .B(_05335_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14294_ (.A1(_04686_),
    .A2(_05214_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _14295_ (.A1(_03614_),
    .A2(_04686_),
    .B1(_05336_),
    .B2(_04255_),
    .C(_05337_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14296_ (.I0(\samples_real[1][10] ),
    .I1(_05231_),
    .S(_04734_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14297_ (.I0(_05229_),
    .I1(_05338_),
    .S(_04722_),
    .Z(_05339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14298_ (.I0(net65),
    .I1(_05339_),
    .S(_05286_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14299_ (.I0(\samples_real[1][10] ),
    .I1(_05340_),
    .S(_04716_),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14300_ (.I0(\samples_real[1][11] ),
    .I1(_05239_),
    .S(_04734_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14301_ (.I0(_05238_),
    .I1(_05341_),
    .S(_04722_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14302_ (.I0(net66),
    .I1(_05342_),
    .S(_05286_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14303_ (.I(_04685_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14304_ (.I0(\samples_real[1][11] ),
    .I1(_05343_),
    .S(_05344_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14305_ (.I0(\samples_real[1][12] ),
    .I1(_05249_),
    .S(_04734_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14306_ (.I0(_05248_),
    .I1(_05345_),
    .S(_04722_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14307_ (.I(_04921_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14308_ (.I0(net67),
    .I1(_05346_),
    .S(_05347_),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14309_ (.I0(\samples_real[1][12] ),
    .I1(_05348_),
    .S(_05344_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14310_ (.I0(\samples_real[1][13] ),
    .I1(_05255_),
    .S(_04734_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14311_ (.I(_04687_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14312_ (.I0(_05254_),
    .I1(_05349_),
    .S(_05350_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14313_ (.I0(net68),
    .I1(_05351_),
    .S(_05347_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14314_ (.I0(\samples_real[1][13] ),
    .I1(_05352_),
    .S(_05344_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14315_ (.I0(\samples_real[1][14] ),
    .I1(_05264_),
    .S(_04734_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14316_ (.I0(_05263_),
    .I1(_05353_),
    .S(_05350_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14317_ (.I0(net69),
    .I1(_05354_),
    .S(_05347_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14318_ (.I0(\samples_real[1][14] ),
    .I1(_05355_),
    .S(_05344_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14319_ (.I0(\samples_real[1][15] ),
    .I1(_05269_),
    .S(_04734_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14320_ (.I0(_05208_),
    .I1(_05356_),
    .S(_05350_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14321_ (.I0(net70),
    .I1(_05357_),
    .S(_05347_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14322_ (.I0(\samples_real[1][15] ),
    .I1(_05358_),
    .S(_05344_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14323_ (.I0(\samples_real[1][1] ),
    .I1(_05277_),
    .S(_04734_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14324_ (.I0(_05276_),
    .I1(_05359_),
    .S(_05350_),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14325_ (.I0(net71),
    .I1(_05360_),
    .S(_05347_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14326_ (.I0(\samples_real[1][1] ),
    .I1(_05361_),
    .S(_05344_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14327_ (.I0(\samples_real[1][2] ),
    .I1(_05283_),
    .S(_04022_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14328_ (.I0(_05282_),
    .I1(_05362_),
    .S(_05350_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14329_ (.I0(net72),
    .I1(_05363_),
    .S(_05347_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14330_ (.I0(\samples_real[1][2] ),
    .I1(_05364_),
    .S(_05344_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14331_ (.I0(\samples_real[1][3] ),
    .I1(_05290_),
    .S(_04022_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14332_ (.I0(_05289_),
    .I1(_05365_),
    .S(_05350_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14333_ (.I0(net73),
    .I1(_05366_),
    .S(_05347_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14334_ (.I0(\samples_real[1][3] ),
    .I1(_05367_),
    .S(_05344_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14335_ (.I0(\samples_real[1][4] ),
    .I1(_05296_),
    .S(_04022_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14336_ (.I0(_05295_),
    .I1(_05368_),
    .S(_05350_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14337_ (.I0(net74),
    .I1(_05369_),
    .S(_05347_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14338_ (.I0(\samples_real[1][4] ),
    .I1(_05370_),
    .S(_05344_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14339_ (.I0(\samples_real[1][5] ),
    .I1(_05303_),
    .S(_04022_),
    .Z(_05371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14340_ (.I0(_05302_),
    .I1(_05371_),
    .S(_05350_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14341_ (.I0(net75),
    .I1(_05372_),
    .S(_05347_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14342_ (.I0(\samples_real[1][5] ),
    .I1(_05373_),
    .S(_05344_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14343_ (.I0(\samples_real[1][6] ),
    .I1(_05309_),
    .S(_04022_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14344_ (.I0(_05308_),
    .I1(_05374_),
    .S(_05350_),
    .Z(_05375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14345_ (.I0(net76),
    .I1(_05375_),
    .S(_05347_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14346_ (.I0(\samples_real[1][6] ),
    .I1(_05376_),
    .S(_04685_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14347_ (.I0(\samples_real[1][7] ),
    .I1(_05316_),
    .S(_04022_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14348_ (.I0(_05315_),
    .I1(_05377_),
    .S(_05350_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14349_ (.I(_04921_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14350_ (.I0(net77),
    .I1(_05378_),
    .S(_05379_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14351_ (.I0(\samples_real[1][7] ),
    .I1(_05380_),
    .S(_04685_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14352_ (.I0(\samples_real[1][8] ),
    .I1(_05322_),
    .S(_04022_),
    .Z(_05381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14353_ (.I0(_05321_),
    .I1(_05381_),
    .S(_04687_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14354_ (.I0(net78),
    .I1(_05382_),
    .S(_05379_),
    .Z(_05383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14355_ (.I0(\samples_real[1][8] ),
    .I1(_05383_),
    .S(_04685_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14356_ (.I0(\samples_real[1][9] ),
    .I1(_05329_),
    .S(_04022_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14357_ (.I0(_05328_),
    .I1(_05384_),
    .S(_04687_),
    .Z(_05385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14358_ (.I0(net79),
    .I1(_05385_),
    .S(_05379_),
    .Z(_05386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14359_ (.I0(\samples_real[1][9] ),
    .I1(_05386_),
    .S(_04685_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14360_ (.A1(_04746_),
    .A2(_05178_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14361_ (.I0(\samples_real[2][0] ),
    .I1(_05387_),
    .S(_04189_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14362_ (.A1(_07703_),
    .A2(_04746_),
    .A3(_05210_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14363_ (.I0(_05388_),
    .I1(_05389_),
    .S(_03762_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14364_ (.A1(_03596_),
    .A2(_05390_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14365_ (.I0(\samples_real[2][0] ),
    .I1(_05214_),
    .S(_04746_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14366_ (.A1(_05391_),
    .A2(_05392_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14367_ (.I0(\samples_real[2][10] ),
    .I1(_05231_),
    .S(_04778_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14368_ (.I0(_05229_),
    .I1(_05393_),
    .S(_04789_),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14369_ (.I0(net65),
    .I1(_05394_),
    .S(_05379_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14370_ (.I0(\samples_real[2][10] ),
    .I1(_05395_),
    .S(_04792_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14371_ (.I0(\samples_real[2][11] ),
    .I1(_05239_),
    .S(_04778_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14372_ (.I0(_05238_),
    .I1(_05396_),
    .S(_04789_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14373_ (.I0(net66),
    .I1(_05397_),
    .S(_05379_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14374_ (.I0(\samples_real[2][11] ),
    .I1(_05398_),
    .S(_04792_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14375_ (.I(_04076_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14376_ (.I0(\samples_real[2][12] ),
    .I1(_05249_),
    .S(_05399_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14377_ (.I0(_05248_),
    .I1(_05400_),
    .S(_04789_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14378_ (.I0(net67),
    .I1(_05401_),
    .S(_05379_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14379_ (.I0(\samples_real[2][12] ),
    .I1(_05402_),
    .S(_04792_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14380_ (.I0(\samples_real[2][13] ),
    .I1(_05255_),
    .S(_05399_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14381_ (.I0(_05254_),
    .I1(_05403_),
    .S(_04789_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14382_ (.I0(net68),
    .I1(_05404_),
    .S(_05379_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14383_ (.I0(\samples_real[2][13] ),
    .I1(_05405_),
    .S(_04792_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14384_ (.I0(\samples_real[2][14] ),
    .I1(_05264_),
    .S(_05399_),
    .Z(_05406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14385_ (.I0(_05263_),
    .I1(_05406_),
    .S(_04789_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14386_ (.I0(net69),
    .I1(_05407_),
    .S(_05379_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14387_ (.I0(\samples_real[2][14] ),
    .I1(_05408_),
    .S(_04792_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14388_ (.I0(\samples_real[2][15] ),
    .I1(_05269_),
    .S(_05399_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14389_ (.I(_04754_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14390_ (.I0(_05208_),
    .I1(_05409_),
    .S(_05410_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14391_ (.I0(net70),
    .I1(_05411_),
    .S(_05379_),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14392_ (.I(_04746_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14393_ (.I0(\samples_real[2][15] ),
    .I1(_05412_),
    .S(_05413_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14394_ (.I0(\samples_real[2][1] ),
    .I1(_05277_),
    .S(_05399_),
    .Z(_05414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14395_ (.I0(_05276_),
    .I1(_05414_),
    .S(_05410_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14396_ (.I0(net71),
    .I1(_05415_),
    .S(_05379_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14397_ (.I0(\samples_real[2][1] ),
    .I1(_05416_),
    .S(_05413_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14398_ (.I0(\samples_real[2][2] ),
    .I1(_05283_),
    .S(_05399_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14399_ (.I0(_05282_),
    .I1(_05417_),
    .S(_05410_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14400_ (.I(_04921_),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14401_ (.I0(net72),
    .I1(_05418_),
    .S(_05419_),
    .Z(_05420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14402_ (.I0(\samples_real[2][2] ),
    .I1(_05420_),
    .S(_05413_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14403_ (.I0(\samples_real[2][3] ),
    .I1(_05290_),
    .S(_05399_),
    .Z(_05421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14404_ (.I0(_05289_),
    .I1(_05421_),
    .S(_05410_),
    .Z(_05422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14405_ (.I0(net73),
    .I1(_05422_),
    .S(_05419_),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14406_ (.I0(\samples_real[2][3] ),
    .I1(_05423_),
    .S(_05413_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14407_ (.I0(\samples_real[2][4] ),
    .I1(_05296_),
    .S(_05399_),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14408_ (.I0(_05295_),
    .I1(_05424_),
    .S(_05410_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14409_ (.I0(net74),
    .I1(_05425_),
    .S(_05419_),
    .Z(_05426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14410_ (.I0(\samples_real[2][4] ),
    .I1(_05426_),
    .S(_05413_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14411_ (.I0(\samples_real[2][5] ),
    .I1(_05303_),
    .S(_05399_),
    .Z(_05427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14412_ (.I0(_05302_),
    .I1(_05427_),
    .S(_05410_),
    .Z(_05428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14413_ (.I0(net75),
    .I1(_05428_),
    .S(_05419_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14414_ (.I0(\samples_real[2][5] ),
    .I1(_05429_),
    .S(_05413_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14415_ (.I0(\samples_real[2][6] ),
    .I1(_05309_),
    .S(_05399_),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14416_ (.I0(_05308_),
    .I1(_05430_),
    .S(_05410_),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14417_ (.I0(net76),
    .I1(_05431_),
    .S(_05419_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14418_ (.I0(\samples_real[2][6] ),
    .I1(_05432_),
    .S(_05413_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14419_ (.I0(\samples_real[2][7] ),
    .I1(_05316_),
    .S(_04076_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14420_ (.I0(_05315_),
    .I1(_05433_),
    .S(_05410_),
    .Z(_05434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14421_ (.I0(net77),
    .I1(_05434_),
    .S(_05419_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14422_ (.I0(\samples_real[2][7] ),
    .I1(_05435_),
    .S(_05413_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14423_ (.I0(\samples_real[2][8] ),
    .I1(_05322_),
    .S(_04076_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14424_ (.I0(_05321_),
    .I1(_05436_),
    .S(_05410_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14425_ (.I0(net78),
    .I1(_05437_),
    .S(_05419_),
    .Z(_05438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14426_ (.I0(\samples_real[2][8] ),
    .I1(_05438_),
    .S(_05413_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14427_ (.I0(\samples_real[2][9] ),
    .I1(_05329_),
    .S(_04076_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14428_ (.I0(_05328_),
    .I1(_05439_),
    .S(_05410_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14429_ (.I0(net79),
    .I1(_05440_),
    .S(_05419_),
    .Z(_05441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14430_ (.I0(\samples_real[2][9] ),
    .I1(_05441_),
    .S(_05413_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14431_ (.A1(_04808_),
    .A2(_05178_),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14432_ (.I0(\samples_real[3][0] ),
    .I1(_05442_),
    .S(_04157_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14433_ (.A1(_07703_),
    .A2(_04808_),
    .A3(_05210_),
    .Z(_05444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14434_ (.I0(_05443_),
    .I1(_05444_),
    .S(_03806_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14435_ (.A1(_05065_),
    .A2(_05445_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14436_ (.I0(\samples_real[3][0] ),
    .I1(_05214_),
    .S(_04808_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14437_ (.A1(_05446_),
    .A2(_05447_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14438_ (.I0(\samples_real[3][10] ),
    .I1(_05231_),
    .S(_04836_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14439_ (.I0(_05229_),
    .I1(_05448_),
    .S(_04851_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14440_ (.I0(net65),
    .I1(_05449_),
    .S(_05419_),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14441_ (.I0(\samples_real[3][10] ),
    .I1(_05450_),
    .S(_04854_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14442_ (.I(_04017_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14443_ (.I0(\samples_real[3][11] ),
    .I1(_05239_),
    .S(_05451_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14444_ (.I0(_05238_),
    .I1(_05452_),
    .S(_04851_),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14445_ (.I0(net66),
    .I1(_05453_),
    .S(_05419_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14446_ (.I0(\samples_real[3][11] ),
    .I1(_05454_),
    .S(_04854_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14447_ (.I0(\samples_real[3][12] ),
    .I1(_05249_),
    .S(_05451_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14448_ (.I0(_05248_),
    .I1(_05455_),
    .S(_04851_),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14449_ (.I(_04921_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14450_ (.I0(net67),
    .I1(_05456_),
    .S(_05457_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14451_ (.I0(\samples_real[3][12] ),
    .I1(_05458_),
    .S(_04854_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14452_ (.I0(\samples_real[3][13] ),
    .I1(_05255_),
    .S(_05451_),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14453_ (.I0(_05254_),
    .I1(_05459_),
    .S(_04851_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14454_ (.I0(net68),
    .I1(_05460_),
    .S(_05457_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14455_ (.I0(\samples_real[3][13] ),
    .I1(_05461_),
    .S(_04854_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14456_ (.I0(\samples_real[3][14] ),
    .I1(_05264_),
    .S(_05451_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14457_ (.I0(_05263_),
    .I1(_05462_),
    .S(_04851_),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14458_ (.I0(net69),
    .I1(_05463_),
    .S(_05457_),
    .Z(_05464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14459_ (.I0(\samples_real[3][14] ),
    .I1(_05464_),
    .S(_04854_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14460_ (.I0(\samples_real[3][15] ),
    .I1(_05269_),
    .S(_05451_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14461_ (.I(_04816_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14462_ (.I0(_05208_),
    .I1(_05465_),
    .S(_05466_),
    .Z(_05467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14463_ (.I0(net70),
    .I1(_05467_),
    .S(_05457_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14464_ (.I(_04808_),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14465_ (.I0(\samples_real[3][15] ),
    .I1(_05468_),
    .S(_05469_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14466_ (.I0(\samples_real[3][1] ),
    .I1(_05277_),
    .S(_05451_),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14467_ (.I0(_05276_),
    .I1(_05470_),
    .S(_05466_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14468_ (.I0(net71),
    .I1(_05471_),
    .S(_05457_),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14469_ (.I0(\samples_real[3][1] ),
    .I1(_05472_),
    .S(_05469_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14470_ (.I0(\samples_real[3][2] ),
    .I1(_05283_),
    .S(_05451_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14471_ (.I0(_05282_),
    .I1(_05473_),
    .S(_05466_),
    .Z(_05474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14472_ (.I0(net72),
    .I1(_05474_),
    .S(_05457_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14473_ (.I0(\samples_real[3][2] ),
    .I1(_05475_),
    .S(_05469_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14474_ (.I0(\samples_real[3][3] ),
    .I1(_05290_),
    .S(_05451_),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14475_ (.I0(_05289_),
    .I1(_05476_),
    .S(_05466_),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14476_ (.I0(net73),
    .I1(_05477_),
    .S(_05457_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14477_ (.I0(\samples_real[3][3] ),
    .I1(_05478_),
    .S(_05469_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14478_ (.I0(\samples_real[3][4] ),
    .I1(_05296_),
    .S(_05451_),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14479_ (.I0(_05295_),
    .I1(_05479_),
    .S(_05466_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14480_ (.I0(net74),
    .I1(_05480_),
    .S(_05457_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14481_ (.I0(\samples_real[3][4] ),
    .I1(_05481_),
    .S(_05469_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14482_ (.I0(\samples_real[3][5] ),
    .I1(_05303_),
    .S(_05451_),
    .Z(_05482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14483_ (.I0(_05302_),
    .I1(_05482_),
    .S(_05466_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14484_ (.I0(net75),
    .I1(_05483_),
    .S(_05457_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14485_ (.I0(\samples_real[3][5] ),
    .I1(_05484_),
    .S(_05469_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14486_ (.I0(\samples_real[3][6] ),
    .I1(_05309_),
    .S(_04017_),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14487_ (.I0(_05308_),
    .I1(_05485_),
    .S(_05466_),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14488_ (.I0(net76),
    .I1(_05486_),
    .S(_05457_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14489_ (.I0(\samples_real[3][6] ),
    .I1(_05487_),
    .S(_05469_),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14490_ (.I0(\samples_real[3][7] ),
    .I1(_05316_),
    .S(_04017_),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14491_ (.I0(_05315_),
    .I1(_05488_),
    .S(_05466_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14492_ (.I(_04921_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14493_ (.I0(net77),
    .I1(_05489_),
    .S(_05490_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14494_ (.I0(\samples_real[3][7] ),
    .I1(_05491_),
    .S(_05469_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14495_ (.I0(\samples_real[3][8] ),
    .I1(_05322_),
    .S(_04017_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14496_ (.I0(_05321_),
    .I1(_05492_),
    .S(_05466_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14497_ (.I0(net78),
    .I1(_05493_),
    .S(_05490_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14498_ (.I0(\samples_real[3][8] ),
    .I1(_05494_),
    .S(_05469_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14499_ (.I0(\samples_real[3][9] ),
    .I1(_05329_),
    .S(_04017_),
    .Z(_05495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14500_ (.I0(_05328_),
    .I1(_05495_),
    .S(_05466_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14501_ (.I0(net79),
    .I1(_05496_),
    .S(_05490_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14502_ (.I0(\samples_real[3][9] ),
    .I1(_05497_),
    .S(_05469_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14503_ (.A1(_04869_),
    .A2(_05178_),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14504_ (.I0(\samples_real[4][0] ),
    .I1(_05498_),
    .S(_04155_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14505_ (.A1(_07703_),
    .A2(_04869_),
    .A3(_05210_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14506_ (.I0(_05499_),
    .I1(_05500_),
    .S(_03760_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14507_ (.A1(_05065_),
    .A2(_05501_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14508_ (.I0(\samples_real[4][0] ),
    .I1(_05214_),
    .S(_04869_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14509_ (.A1(_05502_),
    .A2(_05503_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14510_ (.I0(\samples_real[4][10] ),
    .I1(_05231_),
    .S(_04901_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14511_ (.I0(_05229_),
    .I1(_05504_),
    .S(_04912_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14512_ (.I0(net65),
    .I1(_05505_),
    .S(_05490_),
    .Z(_05506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14513_ (.I0(\samples_real[4][10] ),
    .I1(_05506_),
    .S(_04915_),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14514_ (.I0(\samples_real[4][11] ),
    .I1(_05239_),
    .S(_04901_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14515_ (.I0(_05238_),
    .I1(_05507_),
    .S(_04912_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14516_ (.I0(net66),
    .I1(_05508_),
    .S(_05490_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14517_ (.I0(\samples_real[4][11] ),
    .I1(_05509_),
    .S(_04915_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14518_ (.I(_04079_),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14519_ (.I0(\samples_real[4][12] ),
    .I1(_05249_),
    .S(_05510_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14520_ (.I0(_05248_),
    .I1(_05511_),
    .S(_04912_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14521_ (.I0(net67),
    .I1(_05512_),
    .S(_05490_),
    .Z(_05513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14522_ (.I0(\samples_real[4][12] ),
    .I1(_05513_),
    .S(_04915_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14523_ (.I0(\samples_real[4][13] ),
    .I1(_05255_),
    .S(_05510_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14524_ (.I0(_05254_),
    .I1(_05514_),
    .S(_04912_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14525_ (.I0(net68),
    .I1(_05515_),
    .S(_05490_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14526_ (.I0(\samples_real[4][13] ),
    .I1(_05516_),
    .S(_04915_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14527_ (.I0(\samples_real[4][14] ),
    .I1(_05264_),
    .S(_05510_),
    .Z(_05517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14528_ (.I0(_05263_),
    .I1(_05517_),
    .S(_04912_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14529_ (.I0(net69),
    .I1(_05518_),
    .S(_05490_),
    .Z(_05519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14530_ (.I0(\samples_real[4][14] ),
    .I1(_05519_),
    .S(_04915_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14531_ (.I0(\samples_real[4][15] ),
    .I1(_05269_),
    .S(_05510_),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14532_ (.I(_04877_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14533_ (.I0(_05208_),
    .I1(_05520_),
    .S(_05521_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14534_ (.I0(net70),
    .I1(_05522_),
    .S(_05490_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14535_ (.I(_04869_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14536_ (.I0(\samples_real[4][15] ),
    .I1(_05523_),
    .S(_05524_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14537_ (.I0(\samples_real[4][1] ),
    .I1(_05277_),
    .S(_05510_),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14538_ (.I0(_05276_),
    .I1(_05525_),
    .S(_05521_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14539_ (.I0(net71),
    .I1(_05526_),
    .S(_05490_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14540_ (.I0(\samples_real[4][1] ),
    .I1(_05527_),
    .S(_05524_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14541_ (.I0(\samples_real[4][2] ),
    .I1(_05283_),
    .S(_05510_),
    .Z(_05528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14542_ (.I0(_05282_),
    .I1(_05528_),
    .S(_05521_),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14543_ (.I(_03594_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14544_ (.I0(net72),
    .I1(_05529_),
    .S(_05530_),
    .Z(_05531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14545_ (.I0(\samples_real[4][2] ),
    .I1(_05531_),
    .S(_05524_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14546_ (.I0(\samples_real[4][3] ),
    .I1(_05290_),
    .S(_05510_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14547_ (.I0(_05289_),
    .I1(_05532_),
    .S(_05521_),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14548_ (.I0(net73),
    .I1(_05533_),
    .S(_05530_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14549_ (.I0(\samples_real[4][3] ),
    .I1(_05534_),
    .S(_05524_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14550_ (.I0(\samples_real[4][4] ),
    .I1(_05296_),
    .S(_05510_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14551_ (.I0(_05295_),
    .I1(_05535_),
    .S(_05521_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14552_ (.I0(net74),
    .I1(_05536_),
    .S(_05530_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14553_ (.I0(\samples_real[4][4] ),
    .I1(_05537_),
    .S(_05524_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14554_ (.I0(\samples_real[4][5] ),
    .I1(_05303_),
    .S(_05510_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14555_ (.I0(_05302_),
    .I1(_05538_),
    .S(_05521_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14556_ (.I0(net75),
    .I1(_05539_),
    .S(_05530_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14557_ (.I0(\samples_real[4][5] ),
    .I1(_05540_),
    .S(_05524_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14558_ (.I0(\samples_real[4][6] ),
    .I1(_05309_),
    .S(_05510_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14559_ (.I0(_05308_),
    .I1(_05541_),
    .S(_05521_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14560_ (.I0(net76),
    .I1(_05542_),
    .S(_05530_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14561_ (.I0(\samples_real[4][6] ),
    .I1(_05543_),
    .S(_05524_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14562_ (.I0(\samples_real[4][7] ),
    .I1(_05316_),
    .S(_04079_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14563_ (.I0(_05315_),
    .I1(_05544_),
    .S(_05521_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14564_ (.I0(net77),
    .I1(_05545_),
    .S(_05530_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14565_ (.I0(\samples_real[4][7] ),
    .I1(_05546_),
    .S(_05524_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14566_ (.I0(\samples_real[4][8] ),
    .I1(_05322_),
    .S(_04079_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14567_ (.I0(_05321_),
    .I1(_05547_),
    .S(_05521_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14568_ (.I0(net78),
    .I1(_05548_),
    .S(_05530_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14569_ (.I0(\samples_real[4][8] ),
    .I1(_05549_),
    .S(_05524_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14570_ (.I0(\samples_real[4][9] ),
    .I1(_05329_),
    .S(_04079_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14571_ (.I0(_05328_),
    .I1(_05550_),
    .S(_05521_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14572_ (.I0(net79),
    .I1(_05551_),
    .S(_05530_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14573_ (.I0(\samples_real[4][9] ),
    .I1(_05552_),
    .S(_05524_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14574_ (.A1(_04931_),
    .A2(_05178_),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14575_ (.I0(\samples_real[5][0] ),
    .I1(_05553_),
    .S(_04158_),
    .Z(_05554_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14576_ (.A1(_07703_),
    .A2(_04931_),
    .A3(_05210_),
    .Z(_05555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14577_ (.I0(_05554_),
    .I1(_05555_),
    .S(_03820_),
    .Z(_05556_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14578_ (.A1(_05065_),
    .A2(_05556_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14579_ (.I0(\samples_real[5][0] ),
    .I1(_05214_),
    .S(_04931_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14580_ (.A1(_05557_),
    .A2(_05558_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14581_ (.I0(\samples_real[5][10] ),
    .I1(_05231_),
    .S(_04959_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14582_ (.I0(_05229_),
    .I1(_05559_),
    .S(_04974_),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14583_ (.I0(net65),
    .I1(_05560_),
    .S(_05530_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14584_ (.I0(\samples_real[5][10] ),
    .I1(_05561_),
    .S(_04977_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14585_ (.I(_04020_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14586_ (.I0(\samples_real[5][11] ),
    .I1(_05239_),
    .S(_05562_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14587_ (.I0(_05238_),
    .I1(_05563_),
    .S(_04974_),
    .Z(_05564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14588_ (.I0(net66),
    .I1(_05564_),
    .S(_05530_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14589_ (.I0(\samples_real[5][11] ),
    .I1(_05565_),
    .S(_04977_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14590_ (.I0(\samples_real[5][12] ),
    .I1(_05249_),
    .S(_05562_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14591_ (.I0(_05248_),
    .I1(_05566_),
    .S(_04974_),
    .Z(_05567_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14592_ (.I(_03594_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14593_ (.I0(net67),
    .I1(_05567_),
    .S(_05568_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14594_ (.I0(\samples_real[5][12] ),
    .I1(_05569_),
    .S(_04977_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14595_ (.I0(\samples_real[5][13] ),
    .I1(_05255_),
    .S(_05562_),
    .Z(_05570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14596_ (.I0(_05254_),
    .I1(_05570_),
    .S(_04974_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14597_ (.I0(net68),
    .I1(_05571_),
    .S(_05568_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14598_ (.I0(\samples_real[5][13] ),
    .I1(_05572_),
    .S(_04977_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14599_ (.I0(\samples_real[5][14] ),
    .I1(_05264_),
    .S(_05562_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14600_ (.I0(_05263_),
    .I1(_05573_),
    .S(_04974_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14601_ (.I0(net69),
    .I1(_05574_),
    .S(_05568_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14602_ (.I0(\samples_real[5][14] ),
    .I1(_05575_),
    .S(_04977_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14603_ (.I0(\samples_real[5][15] ),
    .I1(_05269_),
    .S(_05562_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14604_ (.I(_04939_),
    .Z(_05577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14605_ (.I0(_05208_),
    .I1(_05576_),
    .S(_05577_),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14606_ (.I0(net70),
    .I1(_05578_),
    .S(_05568_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14607_ (.I(_04931_),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14608_ (.I0(\samples_real[5][15] ),
    .I1(_05579_),
    .S(_05580_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14609_ (.I0(\samples_real[5][1] ),
    .I1(_05277_),
    .S(_05562_),
    .Z(_05581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14610_ (.I0(_05276_),
    .I1(_05581_),
    .S(_05577_),
    .Z(_05582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14611_ (.I0(net71),
    .I1(_05582_),
    .S(_05568_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14612_ (.I0(\samples_real[5][1] ),
    .I1(_05583_),
    .S(_05580_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14613_ (.I0(\samples_real[5][2] ),
    .I1(_05283_),
    .S(_05562_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14614_ (.I0(_05282_),
    .I1(_05584_),
    .S(_05577_),
    .Z(_05585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14615_ (.I0(net72),
    .I1(_05585_),
    .S(_05568_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14616_ (.I0(\samples_real[5][2] ),
    .I1(_05586_),
    .S(_05580_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14617_ (.I0(\samples_real[5][3] ),
    .I1(_05290_),
    .S(_05562_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14618_ (.I0(_05289_),
    .I1(_05587_),
    .S(_05577_),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14619_ (.I0(net73),
    .I1(_05588_),
    .S(_05568_),
    .Z(_05589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14620_ (.I0(\samples_real[5][3] ),
    .I1(_05589_),
    .S(_05580_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14621_ (.I0(\samples_real[5][4] ),
    .I1(_05296_),
    .S(_05562_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14622_ (.I0(_05295_),
    .I1(_05590_),
    .S(_05577_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14623_ (.I0(net74),
    .I1(_05591_),
    .S(_05568_),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14624_ (.I0(\samples_real[5][4] ),
    .I1(_05592_),
    .S(_05580_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14625_ (.I0(\samples_real[5][5] ),
    .I1(_05303_),
    .S(_05562_),
    .Z(_05593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14626_ (.I0(_05302_),
    .I1(_05593_),
    .S(_05577_),
    .Z(_05594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14627_ (.I0(net75),
    .I1(_05594_),
    .S(_05568_),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14628_ (.I0(\samples_real[5][5] ),
    .I1(_05595_),
    .S(_05580_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14629_ (.I0(\samples_real[5][6] ),
    .I1(_05309_),
    .S(_04020_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14630_ (.I0(_05308_),
    .I1(_05596_),
    .S(_05577_),
    .Z(_05597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14631_ (.I0(net76),
    .I1(_05597_),
    .S(_05568_),
    .Z(_05598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14632_ (.I0(\samples_real[5][6] ),
    .I1(_05598_),
    .S(_05580_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14633_ (.I0(\samples_real[5][7] ),
    .I1(_05316_),
    .S(_04020_),
    .Z(_05599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14634_ (.I0(_05315_),
    .I1(_05599_),
    .S(_05577_),
    .Z(_05600_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14635_ (.I(_03594_),
    .Z(_05601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14636_ (.I0(net77),
    .I1(_05600_),
    .S(_05601_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14637_ (.I0(\samples_real[5][7] ),
    .I1(_05602_),
    .S(_05580_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14638_ (.I0(\samples_real[5][8] ),
    .I1(_05322_),
    .S(_04020_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14639_ (.I0(_05321_),
    .I1(_05603_),
    .S(_05577_),
    .Z(_05604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14640_ (.I0(net78),
    .I1(_05604_),
    .S(_05601_),
    .Z(_05605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14641_ (.I0(\samples_real[5][8] ),
    .I1(_05605_),
    .S(_05580_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14642_ (.I0(\samples_real[5][9] ),
    .I1(_05329_),
    .S(_04020_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14643_ (.I0(_05328_),
    .I1(_05606_),
    .S(_05577_),
    .Z(_05607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14644_ (.I0(net79),
    .I1(_05607_),
    .S(_05601_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14645_ (.I0(\samples_real[5][9] ),
    .I1(_05608_),
    .S(_05580_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14646_ (.A1(_07703_),
    .A2(_04991_),
    .A3(_05210_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14647_ (.A1(_04991_),
    .A2(_05178_),
    .Z(_05610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14648_ (.I0(\samples_real[6][0] ),
    .I1(_05610_),
    .S(_04041_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14649_ (.I0(_05609_),
    .I1(_05611_),
    .S(_04996_),
    .Z(_05612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14650_ (.A1(_05065_),
    .A2(_05612_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14651_ (.I0(\samples_real[6][0] ),
    .I1(_05214_),
    .S(_04991_),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14652_ (.A1(_05613_),
    .A2(_05614_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14653_ (.I0(\samples_real[6][10] ),
    .I1(_05231_),
    .S(_05020_),
    .Z(_05615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14654_ (.I0(_05229_),
    .I1(_05615_),
    .S(_05028_),
    .Z(_05616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14655_ (.I0(net65),
    .I1(_05616_),
    .S(_05601_),
    .Z(_05617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14656_ (.I0(\samples_real[6][10] ),
    .I1(_05617_),
    .S(_05037_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14657_ (.I(_04040_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14658_ (.I0(\samples_real[6][11] ),
    .I1(_05239_),
    .S(_05618_),
    .Z(_05619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14659_ (.I0(_05238_),
    .I1(_05619_),
    .S(_05028_),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14660_ (.I0(net66),
    .I1(_05620_),
    .S(_05601_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14661_ (.I0(\samples_real[6][11] ),
    .I1(_05621_),
    .S(_05037_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14662_ (.I0(\samples_real[6][12] ),
    .I1(_05249_),
    .S(_05618_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14663_ (.I0(_05248_),
    .I1(_05622_),
    .S(_05028_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14664_ (.I0(net67),
    .I1(_05623_),
    .S(_05601_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14665_ (.I0(\samples_real[6][12] ),
    .I1(_05624_),
    .S(_05037_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14666_ (.I0(\samples_real[6][13] ),
    .I1(_05255_),
    .S(_05618_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14667_ (.I(_04995_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14668_ (.I0(_05254_),
    .I1(_05625_),
    .S(_05626_),
    .Z(_05627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14669_ (.I0(net68),
    .I1(_05627_),
    .S(_05601_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14670_ (.I0(\samples_real[6][13] ),
    .I1(_05628_),
    .S(_05037_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14671_ (.I0(\samples_real[6][14] ),
    .I1(_05264_),
    .S(_05618_),
    .Z(_05629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14672_ (.I0(_05263_),
    .I1(_05629_),
    .S(_05626_),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14673_ (.I0(net69),
    .I1(_05630_),
    .S(_05601_),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14674_ (.I0(\samples_real[6][14] ),
    .I1(_05631_),
    .S(_05037_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14675_ (.I0(\samples_real[6][15] ),
    .I1(_05269_),
    .S(_05618_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14676_ (.I0(_05208_),
    .I1(_05632_),
    .S(_05626_),
    .Z(_05633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14677_ (.I0(net70),
    .I1(_05633_),
    .S(_05601_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _14678_ (.I(_04991_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14679_ (.I0(\samples_real[6][15] ),
    .I1(_05634_),
    .S(_05635_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14680_ (.I0(\samples_real[6][1] ),
    .I1(_05277_),
    .S(_05618_),
    .Z(_05636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14681_ (.I0(_05276_),
    .I1(_05636_),
    .S(_05626_),
    .Z(_05637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14682_ (.I0(net71),
    .I1(_05637_),
    .S(_05601_),
    .Z(_05638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14683_ (.I0(\samples_real[6][1] ),
    .I1(_05638_),
    .S(_05635_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14684_ (.I0(\samples_real[6][2] ),
    .I1(_05283_),
    .S(_05618_),
    .Z(_05639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14685_ (.I0(_05282_),
    .I1(_05639_),
    .S(_05626_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14686_ (.I0(net72),
    .I1(_05640_),
    .S(_03595_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14687_ (.I0(\samples_real[6][2] ),
    .I1(_05641_),
    .S(_05635_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14688_ (.I0(\samples_real[6][3] ),
    .I1(_05290_),
    .S(_05618_),
    .Z(_05642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14689_ (.I0(_05289_),
    .I1(_05642_),
    .S(_05626_),
    .Z(_05643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14690_ (.I0(net73),
    .I1(_05643_),
    .S(_03595_),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14691_ (.I0(\samples_real[6][3] ),
    .I1(_05644_),
    .S(_05635_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14692_ (.I0(\samples_real[6][4] ),
    .I1(_05296_),
    .S(_05618_),
    .Z(_05645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14693_ (.I0(_05295_),
    .I1(_05645_),
    .S(_05626_),
    .Z(_05646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14694_ (.I0(net74),
    .I1(_05646_),
    .S(_03595_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14695_ (.I0(\samples_real[6][4] ),
    .I1(_05647_),
    .S(_05635_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14696_ (.I0(\samples_real[6][5] ),
    .I1(_05303_),
    .S(_05618_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14697_ (.I0(_05302_),
    .I1(_05648_),
    .S(_05626_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14698_ (.I0(net75),
    .I1(_05649_),
    .S(_03595_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14699_ (.I0(\samples_real[6][5] ),
    .I1(_05650_),
    .S(_05635_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14700_ (.I0(\samples_real[6][6] ),
    .I1(_05309_),
    .S(_04040_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14701_ (.I0(_05308_),
    .I1(_05651_),
    .S(_05626_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14702_ (.I0(net76),
    .I1(_05652_),
    .S(_03595_),
    .Z(_05653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14703_ (.I0(\samples_real[6][6] ),
    .I1(_05653_),
    .S(_05635_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14704_ (.I0(\samples_real[6][7] ),
    .I1(_05316_),
    .S(_04040_),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14705_ (.I0(_05315_),
    .I1(_05654_),
    .S(_05626_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14706_ (.I0(net77),
    .I1(_05655_),
    .S(_03595_),
    .Z(_05656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14707_ (.I0(\samples_real[6][7] ),
    .I1(_05656_),
    .S(_05635_),
    .Z(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14708_ (.I0(\samples_real[6][8] ),
    .I1(_05322_),
    .S(_04040_),
    .Z(_05657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14709_ (.I0(_05321_),
    .I1(_05657_),
    .S(_04995_),
    .Z(_05658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14710_ (.I0(net78),
    .I1(_05658_),
    .S(_03595_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14711_ (.I0(\samples_real[6][8] ),
    .I1(_05659_),
    .S(_05635_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14712_ (.I0(\samples_real[6][9] ),
    .I1(_05329_),
    .S(_04040_),
    .Z(_05660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14713_ (.I0(_05328_),
    .I1(_05660_),
    .S(_04995_),
    .Z(_05661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14714_ (.I0(net79),
    .I1(_05661_),
    .S(_03595_),
    .Z(_05662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14715_ (.I0(\samples_real[6][9] ),
    .I1(_05662_),
    .S(_05635_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14716_ (.A1(\samples_real[7][0] ),
    .A2(_05051_),
    .B1(_05055_),
    .B2(_05178_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14717_ (.A1(_05059_),
    .A2(_05211_),
    .B1(_05663_),
    .B2(_03753_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14718_ (.A1(_05065_),
    .A2(_05664_),
    .Z(_05665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14719_ (.I0(_05214_),
    .I1(\samples_real[7][0] ),
    .S(_05054_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14720_ (.A1(_05665_),
    .A2(_05666_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14721_ (.I0(\samples_real[7][10] ),
    .I1(_05231_),
    .S(_05093_),
    .Z(_05667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14722_ (.I0(_05229_),
    .I1(_05667_),
    .S(_05095_),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14723_ (.I0(net65),
    .I1(_05668_),
    .S(_05107_),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14724_ (.I0(_05669_),
    .I1(\samples_real[7][10] ),
    .S(_05101_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14725_ (.I0(\samples_real[7][11] ),
    .I1(_05239_),
    .S(_05093_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14726_ (.I0(_05238_),
    .I1(_05670_),
    .S(_05095_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14727_ (.I0(net66),
    .I1(_05671_),
    .S(_05107_),
    .Z(_05672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14728_ (.I0(_05672_),
    .I1(\samples_real[7][11] ),
    .S(_05101_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14729_ (.I0(\samples_real[7][12] ),
    .I1(_05249_),
    .S(_05093_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14730_ (.I0(_05248_),
    .I1(_05673_),
    .S(_05095_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14731_ (.I0(net67),
    .I1(_05674_),
    .S(_05107_),
    .Z(_05675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14732_ (.I0(_05675_),
    .I1(\samples_real[7][12] ),
    .S(_05101_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14733_ (.I0(\samples_real[7][13] ),
    .I1(_05255_),
    .S(_05093_),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14734_ (.I0(_05254_),
    .I1(_05676_),
    .S(_05095_),
    .Z(_05677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14735_ (.I0(net68),
    .I1(_05677_),
    .S(_05107_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14736_ (.I0(_05678_),
    .I1(\samples_real[7][13] ),
    .S(_05101_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14737_ (.I(_04013_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14738_ (.I0(\samples_real[7][14] ),
    .I1(_05264_),
    .S(_05679_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14739_ (.I(_05057_),
    .Z(_05681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14740_ (.I0(_05263_),
    .I1(_05680_),
    .S(_05681_),
    .Z(_05682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14741_ (.I0(net69),
    .I1(_05682_),
    .S(_05107_),
    .Z(_05683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14742_ (.I0(_05683_),
    .I1(\samples_real[7][14] ),
    .S(_05101_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14743_ (.I0(\samples_real[7][15] ),
    .I1(_05269_),
    .S(_05679_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14744_ (.I0(_05208_),
    .I1(_05684_),
    .S(_05681_),
    .Z(_05685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14745_ (.I0(net70),
    .I1(_05685_),
    .S(_05107_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _14746_ (.I(_05054_),
    .Z(_05687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14747_ (.I0(_05686_),
    .I1(\samples_real[7][15] ),
    .S(_05687_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14748_ (.I0(\samples_real[7][1] ),
    .I1(_05277_),
    .S(_05679_),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14749_ (.I0(_05276_),
    .I1(_05688_),
    .S(_05681_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14750_ (.I0(net71),
    .I1(_05689_),
    .S(_05107_),
    .Z(_05690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14751_ (.I0(_05690_),
    .I1(\samples_real[7][1] ),
    .S(_05687_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14752_ (.I0(\samples_real[7][2] ),
    .I1(_05283_),
    .S(_05679_),
    .Z(_05691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14753_ (.I0(_05282_),
    .I1(_05691_),
    .S(_05681_),
    .Z(_05692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14754_ (.I0(net72),
    .I1(_05692_),
    .S(_04578_),
    .Z(_05693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14755_ (.I0(_05693_),
    .I1(\samples_real[7][2] ),
    .S(_05687_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14756_ (.I0(\samples_real[7][3] ),
    .I1(_05290_),
    .S(_05679_),
    .Z(_05694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14757_ (.I0(_05289_),
    .I1(_05694_),
    .S(_05681_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14758_ (.I0(net73),
    .I1(_05695_),
    .S(_04578_),
    .Z(_05696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14759_ (.I0(_05696_),
    .I1(\samples_real[7][3] ),
    .S(_05687_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14760_ (.I0(\samples_real[7][4] ),
    .I1(_05296_),
    .S(_05679_),
    .Z(_05697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14761_ (.I0(_05295_),
    .I1(_05697_),
    .S(_05681_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14762_ (.I0(net74),
    .I1(_05698_),
    .S(_04578_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14763_ (.I0(_05699_),
    .I1(\samples_real[7][4] ),
    .S(_05687_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14764_ (.I0(\samples_real[7][5] ),
    .I1(_05303_),
    .S(_05679_),
    .Z(_05700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14765_ (.I0(_05302_),
    .I1(_05700_),
    .S(_05681_),
    .Z(_05701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14766_ (.I0(net75),
    .I1(_05701_),
    .S(_04578_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14767_ (.I0(_05702_),
    .I1(\samples_real[7][5] ),
    .S(_05687_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14768_ (.I0(\samples_real[7][6] ),
    .I1(_05309_),
    .S(_05679_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14769_ (.I0(_05308_),
    .I1(_05703_),
    .S(_05681_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14770_ (.I0(net76),
    .I1(_05704_),
    .S(_04578_),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14771_ (.I0(_05705_),
    .I1(\samples_real[7][6] ),
    .S(_05687_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14772_ (.I0(\samples_real[7][7] ),
    .I1(_05316_),
    .S(_05679_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14773_ (.I0(_05315_),
    .I1(_05706_),
    .S(_05681_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14774_ (.I0(net77),
    .I1(_05707_),
    .S(_04578_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14775_ (.I0(_05708_),
    .I1(\samples_real[7][7] ),
    .S(_05687_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14776_ (.I0(\samples_real[7][8] ),
    .I1(_05322_),
    .S(_05679_),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14777_ (.I0(_05321_),
    .I1(_05709_),
    .S(_05681_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14778_ (.I0(net78),
    .I1(_05710_),
    .S(_04578_),
    .Z(_05711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14779_ (.I0(_05711_),
    .I1(\samples_real[7][8] ),
    .S(_05687_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14780_ (.I0(\samples_real[7][9] ),
    .I1(_05329_),
    .S(_04013_),
    .Z(_05712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14781_ (.I0(_05328_),
    .I1(_05712_),
    .S(_05057_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14782_ (.I0(net79),
    .I1(_05713_),
    .S(_04578_),
    .Z(_05714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14783_ (.I0(_05714_),
    .I1(\samples_real[7][9] ),
    .S(_05687_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14784_ (.A1(_05065_),
    .A2(_07773_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14785_ (.A1(_07789_),
    .A2(_03634_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14786_ (.A1(_05716_),
    .A2(_04257_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14787_ (.I0(\stage[0] ),
    .I1(_05715_),
    .S(_05717_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14788_ (.A1(_05065_),
    .A2(_07776_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14789_ (.I0(\stage[1] ),
    .I1(_05718_),
    .S(_05717_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14790_ (.A1(_05065_),
    .A2(_07790_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14791_ (.I0(_00567_),
    .I1(_05719_),
    .S(_05717_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14792_ (.I(_08207_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14793_ (.I(_07073_),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _14794_ (.A1(_05721_),
    .A2(_08297_),
    .A3(_08299_),
    .A4(_08301_),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14795_ (.A1(_08308_),
    .A2(_06803_),
    .B(_08307_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14796_ (.A1(_05722_),
    .A2(_05723_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14797_ (.A1(_08254_),
    .A2(_08290_),
    .A3(_08236_),
    .A4(_08266_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14798_ (.A1(_08296_),
    .A2(_05724_),
    .B(_05725_),
    .C(_08283_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14799_ (.I(_08253_),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14800_ (.A1(_08289_),
    .A2(_08283_),
    .Z(_05728_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14801_ (.A1(_08282_),
    .A2(_05728_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14802_ (.A1(_08266_),
    .A2(_05729_),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14803_ (.A1(_08265_),
    .A2(_05730_),
    .B(_08254_),
    .ZN(_05731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14804_ (.A1(_05727_),
    .A2(_05731_),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14805_ (.A1(_08236_),
    .A2(_05732_),
    .B(_08235_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14806_ (.A1(_05726_),
    .A2(_05733_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14807_ (.A1(_08222_),
    .A2(_05734_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14808_ (.A1(_08221_),
    .A2(_05735_),
    .B(_08208_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14809_ (.A1(_05720_),
    .A2(_05736_),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14810_ (.A1(_08193_),
    .A2(_05737_),
    .B(_08192_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14811_ (.A1(_03845_),
    .A2(_03875_),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14812_ (.A1(_03789_),
    .A2(_03817_),
    .A3(_05739_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14813_ (.A1(_00011_),
    .A2(_05740_),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14814_ (.I0(\samples_imag[2][15] ),
    .I1(\samples_imag[6][15] ),
    .S(_03679_),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14815_ (.A1(_03717_),
    .A2(\samples_imag[4][15] ),
    .Z(_05743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14816_ (.I0(\samples_imag[3][15] ),
    .I1(\samples_imag[7][15] ),
    .S(_03678_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14817_ (.A1(_03688_),
    .A2(\samples_imag[1][15] ),
    .Z(_05745_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _14818_ (.I0(_05742_),
    .I1(_05743_),
    .I2(_05744_),
    .I3(_05745_),
    .S0(_03693_),
    .S1(_03676_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14819_ (.A1(\samples_imag[5][15] ),
    .A2(_03820_),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _14820_ (.A1(\samples_imag[0][15] ),
    .A2(_03712_),
    .B1(_05746_),
    .B2(_05747_),
    .C(_00009_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14821_ (.A1(_06918_),
    .A2(_05748_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14822_ (.A1(_06567_),
    .A2(_06745_),
    .A3(_05749_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14823_ (.A1(_03724_),
    .A2(_03887_),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14824_ (.A1(_03700_),
    .A2(_04001_),
    .A3(_05751_),
    .ZN(_05752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14825_ (.A1(_03725_),
    .A2(_05752_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14826_ (.A1(_05741_),
    .A2(_05750_),
    .A3(_05753_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14827_ (.A1(_06609_),
    .A2(_06614_),
    .ZN(_05755_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14828_ (.A1(_06598_),
    .A2(_06661_),
    .A3(_05755_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14829_ (.A1(_08103_),
    .A2(_08106_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14830_ (.A1(_08113_),
    .A2(_08131_),
    .A3(_05757_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14831_ (.A1(_06519_),
    .A2(_06499_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14832_ (.A1(_06508_),
    .A2(_06531_),
    .A3(_05759_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14833_ (.A1(_06675_),
    .A2(_08138_),
    .Z(_05761_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14834_ (.A1(_06672_),
    .A2(_06603_),
    .A3(_05761_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14835_ (.A1(_05760_),
    .A2(_05762_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14836_ (.A1(_05756_),
    .A2(_05758_),
    .A3(_05763_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14837_ (.A1(_00016_),
    .A2(_00017_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14838_ (.A1(_06557_),
    .A2(_06589_),
    .A3(_05765_),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14839_ (.A1(_08167_),
    .A2(_06544_),
    .A3(_05766_),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14840_ (.A1(_03714_),
    .A2(_03979_),
    .Z(_05768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14841_ (.A1(_00010_),
    .A2(_05768_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14842_ (.A1(_05764_),
    .A2(_05767_),
    .A3(_05769_),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14843_ (.A1(_00012_),
    .A2(_03989_),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14844_ (.I(_03925_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14845_ (.A1(_00016_),
    .A2(_05772_),
    .Z(_05773_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14846_ (.A1(_06523_),
    .A2(_06513_),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14847_ (.A1(_06561_),
    .A2(_06526_),
    .A3(_05774_),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14848_ (.A1(_06553_),
    .A2(_06621_),
    .Z(_05776_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14849_ (.A1(_08129_),
    .A2(_06728_),
    .A3(_05776_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14850_ (.A1(_08117_),
    .A2(_06776_),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14851_ (.A1(_08109_),
    .A2(_08128_),
    .A3(_05778_),
    .ZN(_05779_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14852_ (.A1(_05775_),
    .A2(_05777_),
    .A3(_05779_),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14853_ (.I(_03969_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14854_ (.A1(_00017_),
    .A2(_05781_),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14855_ (.A1(_05780_),
    .A2(_05782_),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14856_ (.A1(_05771_),
    .A2(_05773_),
    .A3(_05783_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14857_ (.A1(_05770_),
    .A2(_05784_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14858_ (.A1(_05738_),
    .A2(_05754_),
    .A3(_05785_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14859_ (.I0(\temp_imag[0] ),
    .I1(_05786_),
    .S(_03636_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14860_ (.I(_07972_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _14861_ (.A1(_08017_),
    .A2(_08030_),
    .A3(_08041_),
    .A4(_08066_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14862_ (.A1(_08086_),
    .A2(_08093_),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14863_ (.A1(_08085_),
    .A2(_05789_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14864_ (.A1(_08094_),
    .A2(_08096_),
    .A3(_08100_),
    .A4(_08086_),
    .Z(_05791_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14865_ (.A1(_08099_),
    .A2(_06341_),
    .ZN(_05792_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14866_ (.A1(_08076_),
    .A2(_03981_),
    .A3(_05791_),
    .A4(_05792_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _14867_ (.A1(_08076_),
    .A2(_05790_),
    .B(_05793_),
    .C(_08075_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14868_ (.I(_08029_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14869_ (.A1(_08065_),
    .A2(_08041_),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14870_ (.A1(_08040_),
    .A2(_05796_),
    .B(_08030_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14871_ (.A1(_05795_),
    .A2(_05797_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14872_ (.A1(_08017_),
    .A2(_05798_),
    .B(_08016_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14873_ (.A1(_05788_),
    .A2(_05794_),
    .B(_05799_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14874_ (.A1(_07998_),
    .A2(_05800_),
    .Z(_05801_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14875_ (.A1(_07997_),
    .A2(_05801_),
    .Z(_05802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14876_ (.A1(_07983_),
    .A2(_05802_),
    .Z(_05803_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14877_ (.A1(_07982_),
    .A2(_05803_),
    .B(_07973_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14878_ (.A1(_05787_),
    .A2(_05804_),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14879_ (.A1(_07964_),
    .A2(_05805_),
    .B(_07963_),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14880_ (.A1(_00016_),
    .A2(_05781_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14881_ (.A1(_00011_),
    .A2(_03865_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14882_ (.A1(_05889_),
    .A2(_05902_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14883_ (.A1(_05929_),
    .A2(_05934_),
    .A3(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14884_ (.A1(_05884_),
    .A2(_07893_),
    .Z(_05811_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14885_ (.A1(_07902_),
    .A2(_06005_),
    .A3(_05811_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14886_ (.A1(_05810_),
    .A2(_05812_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14887_ (.A1(_06008_),
    .A2(_06027_),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14888_ (.A1(_06059_),
    .A2(_06079_),
    .A3(_05814_),
    .ZN(_05815_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14889_ (.A1(_06074_),
    .A2(_05937_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14890_ (.A1(_05941_),
    .A2(_05962_),
    .A3(_05816_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14891_ (.A1(_05815_),
    .A2(_05817_),
    .ZN(_05818_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14892_ (.A1(_07957_),
    .A2(_07894_),
    .Z(_05819_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14893_ (.A1(_05898_),
    .A2(_05920_),
    .A3(_05819_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14894_ (.A1(_07899_),
    .A2(_05977_),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14895_ (.A1(_05990_),
    .A2(_06023_),
    .A3(_05821_),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14896_ (.A1(_07912_),
    .A2(_07915_),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14897_ (.A1(_07910_),
    .A2(_05985_),
    .A3(_05823_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14898_ (.A1(_05820_),
    .A2(_05822_),
    .A3(_05824_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14899_ (.A1(_05813_),
    .A2(_05818_),
    .A3(_05825_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14900_ (.A1(_00012_),
    .A2(_04001_),
    .Z(_05827_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14901_ (.A1(_07909_),
    .A2(_05826_),
    .A3(_05827_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14902_ (.A1(_05807_),
    .A2(_05808_),
    .A3(_05828_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14903_ (.A1(_07908_),
    .A2(_05950_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14904_ (.A1(_06094_),
    .A2(_06256_),
    .A3(_05830_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14905_ (.A1(_03725_),
    .A2(_03989_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14906_ (.A1(_00017_),
    .A2(_05772_),
    .Z(_05833_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14907_ (.A1(_05832_),
    .A2(_05833_),
    .ZN(_05834_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14908_ (.A1(_05917_),
    .A2(_05969_),
    .A3(_05834_),
    .ZN(_05835_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14909_ (.A1(_03827_),
    .A2(_05751_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14910_ (.A1(_00010_),
    .A2(_05836_),
    .Z(_05837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14911_ (.I0(\samples_real[3][15] ),
    .I1(\samples_real[7][15] ),
    .S(_03680_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14912_ (.A1(\samples_real[5][15] ),
    .A2(_03703_),
    .B1(_05838_),
    .B2(_03672_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14913_ (.A1(_03689_),
    .A2(\samples_real[4][15] ),
    .Z(_05840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14914_ (.A1(_03689_),
    .A2(\samples_real[1][15] ),
    .B1(_05840_),
    .B2(_03684_),
    .ZN(_05841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14915_ (.I0(\samples_real[2][15] ),
    .I1(\samples_real[6][15] ),
    .S(_03680_),
    .Z(_05842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14916_ (.A1(_03745_),
    .A2(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _14917_ (.A1(_03685_),
    .A2(_05839_),
    .B1(_05841_),
    .B2(_03673_),
    .C(_05843_),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14918_ (.A1(\samples_real[0][15] ),
    .A2(_03712_),
    .B(_05844_),
    .C(_00009_),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14919_ (.A1(_06125_),
    .A2(_06182_),
    .A3(_05765_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14920_ (.A1(_07938_),
    .A2(_05995_),
    .A3(_05846_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14921_ (.A1(_05964_),
    .A2(_05845_),
    .A3(_05847_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14922_ (.A1(_05892_),
    .A2(_05837_),
    .A3(_05848_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14923_ (.A1(_05831_),
    .A2(_05835_),
    .A3(_05849_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _14924_ (.A1(_05806_),
    .A2(_05829_),
    .A3(_05850_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14925_ (.I0(\temp_real[0] ),
    .I1(_05851_),
    .S(_03636_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14926_ (.A1(_00000_),
    .A2(_00002_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14927_ (.A(_05852_),
    .B(_05853_),
    .CI(_05854_),
    .CO(_05855_),
    .S(_05856_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14928_ (.A(_05852_),
    .B(_05857_),
    .CI(_05858_),
    .CO(_05859_),
    .S(_05860_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14929_ (.A(_05862_),
    .B(_05863_),
    .CI(_05864_),
    .CO(_05865_),
    .S(_05866_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14930_ (.A(_05867_),
    .B(_05868_),
    .CI(_05869_),
    .CO(_05870_),
    .S(_05871_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14931_ (.A(_05867_),
    .B(_05872_),
    .CI(_05873_),
    .CO(_05874_),
    .S(_05875_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14932_ (.A(_05877_),
    .B(_00014_),
    .CI(_05878_),
    .CO(_05879_),
    .S(_05880_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14933_ (.A(_05881_),
    .B(_05882_),
    .CI(_05883_),
    .CO(_05884_),
    .S(_05885_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14934_ (.A(_05886_),
    .B(_05887_),
    .CI(_05888_),
    .CO(_05889_),
    .S(_05890_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14935_ (.A(_05891_),
    .B(_05892_),
    .CI(_05893_),
    .CO(_05887_),
    .S(_05894_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14936_ (.A(_05895_),
    .B(_05896_),
    .CI(_05897_),
    .CO(_05898_),
    .S(_05899_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14937_ (.A(_05890_),
    .B(_05900_),
    .CI(_05901_),
    .CO(_05902_),
    .S(_05903_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14938_ (.A(_05894_),
    .B(_05904_),
    .CI(_05905_),
    .CO(_05900_),
    .S(_05906_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14939_ (.A(_05907_),
    .B(_05908_),
    .CI(_05909_),
    .CO(_05910_),
    .S(_05911_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14940_ (.A(_05912_),
    .B(_05913_),
    .CI(_05914_),
    .CO(_05915_),
    .S(_05916_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14941_ (.A(_05917_),
    .B(_05918_),
    .CI(_05919_),
    .CO(_05920_),
    .S(_05921_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14942_ (.A(_05922_),
    .B(_05923_),
    .CI(_05924_),
    .CO(_05925_),
    .S(_05926_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14943_ (.A(_05893_),
    .B(_05927_),
    .CI(_05928_),
    .CO(_05929_),
    .S(_05930_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14944_ (.A(_05931_),
    .B(_05932_),
    .CI(_05933_),
    .CO(_05934_),
    .S(_05935_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14945_ (.A(_05930_),
    .B(_05936_),
    .CI(_05935_),
    .CO(_05937_),
    .S(_05938_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14946_ (.A(_05903_),
    .B(_05939_),
    .CI(_05940_),
    .CO(_05941_),
    .S(_05942_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14947_ (.A(_05906_),
    .B(_05943_),
    .CI(_05944_),
    .CO(_05939_),
    .S(_05945_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14948_ (.A(_05946_),
    .B(_05947_),
    .CI(_05948_),
    .CO(_05943_),
    .S(_05949_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14949_ (.A(_05908_),
    .B(_05950_),
    .CI(_05951_),
    .CO(_05952_),
    .S(_05953_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14950_ (.A(_05954_),
    .B(_05955_),
    .CI(_05956_),
    .CO(_05957_),
    .S(_05958_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14951_ (.A(_05959_),
    .B(_05960_),
    .CI(_05961_),
    .CO(_05962_),
    .S(_05963_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14952_ (.A(_05964_),
    .B(_05965_),
    .CI(_05966_),
    .CO(_05967_),
    .S(_05968_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14953_ (.A(_05909_),
    .B(_05951_),
    .CI(_05969_),
    .CO(_05970_),
    .S(_05971_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14954_ (.A(_05973_),
    .B(_05974_),
    .CI(_05975_),
    .CO(_05976_),
    .S(_05977_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14955_ (.A(_05971_),
    .B(_05978_),
    .CI(_05977_),
    .CO(_05979_),
    .S(_05980_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14956_ (.A(_05982_),
    .B(_05983_),
    .CI(_05984_),
    .CO(_05985_),
    .S(_05986_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14957_ (.A(_05987_),
    .B(_05988_),
    .CI(_05989_),
    .CO(_05990_),
    .S(_05991_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14958_ (.A(_05992_),
    .B(_05993_),
    .CI(_05994_),
    .CO(_05995_),
    .S(_05996_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14959_ (.A(_05989_),
    .B(_05997_),
    .CI(_05998_),
    .CO(_05999_),
    .S(_06000_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14960_ (.A(_06001_),
    .B(_06002_),
    .CI(_06003_),
    .CO(_06004_),
    .S(_06005_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14961_ (.A(_06006_),
    .B(_05996_),
    .CI(_06007_),
    .CO(_06008_),
    .S(_06009_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14962_ (.A(_05928_),
    .B(_05972_),
    .CI(_05932_),
    .CO(_05981_),
    .S(_06010_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14963_ (.A(_05933_),
    .B(_06011_),
    .CI(_06001_),
    .CO(_06012_),
    .S(_06013_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14964_ (.A(_06012_),
    .B(_06000_),
    .CI(_06014_),
    .CO(_06007_),
    .S(_06015_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14965_ (.A(_05998_),
    .B(_06016_),
    .CI(_06017_),
    .CO(_06018_),
    .S(_06019_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14966_ (.A(_06020_),
    .B(_06021_),
    .CI(_06022_),
    .CO(_06023_),
    .S(_06024_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14967_ (.A(_05942_),
    .B(_06025_),
    .CI(_06026_),
    .CO(_06027_),
    .S(_06028_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14968_ (.A(_05945_),
    .B(_06029_),
    .CI(_06030_),
    .CO(_06025_),
    .S(_06031_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14969_ (.A(_05949_),
    .B(_06032_),
    .CI(_06033_),
    .CO(_06029_),
    .S(_06034_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14970_ (.A(_06035_),
    .B(_06036_),
    .CI(_06037_),
    .CO(_06032_),
    .S(_06038_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14971_ (.A(_06039_),
    .B(_06040_),
    .CI(_05972_),
    .CO(_06036_),
    .S(_06041_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14972_ (.A(_06042_),
    .B(_06043_),
    .CI(_06044_),
    .CO(_06045_),
    .S(_06046_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14973_ (.A(_06047_),
    .B(_06048_),
    .CI(_05980_),
    .CO(_05984_),
    .S(_06049_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14974_ (.A(_05927_),
    .B(_06050_),
    .CI(_06051_),
    .CO(_06052_),
    .S(_06053_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14975_ (.A(_06010_),
    .B(_06054_),
    .CI(_06055_),
    .CO(_06056_),
    .S(_06057_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _14976_ (.A(_06009_),
    .B(_06058_),
    .CI(_06024_),
    .CO(_06059_),
    .S(_06060_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14977_ (.A(_06056_),
    .B(_06061_),
    .CI(_06062_),
    .CO(_06058_),
    .S(_06063_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14978_ (.A(_05972_),
    .B(_05932_),
    .CI(_06065_),
    .CO(_06054_),
    .S(_06066_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14979_ (.A(_05975_),
    .B(_05989_),
    .CI(_05997_),
    .CO(_06067_),
    .S(_06068_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14980_ (.A(_06069_),
    .B(_06067_),
    .CI(_06070_),
    .CO(_06064_),
    .S(_06071_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14981_ (.A(_06072_),
    .B(_06060_),
    .CI(_06073_),
    .CO(_06074_),
    .S(_06075_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14982_ (.A(_06028_),
    .B(_06077_),
    .CI(_06078_),
    .CO(_06079_),
    .S(_06080_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14983_ (.A(_06031_),
    .B(_06081_),
    .CI(_06082_),
    .CO(_06077_),
    .S(_06083_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14984_ (.A(_06034_),
    .B(_06085_),
    .CI(_06045_),
    .CO(_06081_),
    .S(_06086_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14985_ (.A(_06038_),
    .B(_06087_),
    .CI(_06088_),
    .CO(_06085_),
    .S(_06089_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14986_ (.A(_06041_),
    .B(_06090_),
    .CI(_06091_),
    .CO(_06087_),
    .S(_06092_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14987_ (.A(_06093_),
    .B(_06094_),
    .CI(_06095_),
    .CO(_06096_),
    .S(_06097_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14988_ (.A(_06098_),
    .B(_06099_),
    .CI(_06100_),
    .CO(_06101_),
    .S(_06102_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14989_ (.A(_05928_),
    .B(_06103_),
    .CI(_06104_),
    .CO(_06105_),
    .S(_06106_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14990_ (.A(_06066_),
    .B(_06107_),
    .CI(_06068_),
    .CO(_06108_),
    .S(_06109_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14991_ (.A(_06063_),
    .B(_06111_),
    .CI(_06112_),
    .CO(_06073_),
    .S(_06113_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14992_ (.A(_06108_),
    .B(_06114_),
    .CI(_06115_),
    .CO(_06111_),
    .S(_06116_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14993_ (.A(_06095_),
    .B(_05974_),
    .CI(_05987_),
    .CO(_06110_),
    .S(_06117_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14994_ (.A(_06118_),
    .B(_06113_),
    .CI(_06119_),
    .CO(_06120_),
    .S(_06121_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14995_ (.A(_06080_),
    .B(_06123_),
    .CI(_06124_),
    .CO(_06125_),
    .S(_06126_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14996_ (.A(_06083_),
    .B(_06127_),
    .CI(_06128_),
    .CO(_06123_),
    .S(_06129_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14997_ (.A(_06086_),
    .B(_06130_),
    .CI(_06131_),
    .CO(_06127_),
    .S(_06132_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14998_ (.A(_06089_),
    .B(_06134_),
    .CI(_06135_),
    .CO(_06130_),
    .S(_06136_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _14999_ (.A(_06092_),
    .B(_06138_),
    .CI(_06139_),
    .CO(_06134_),
    .S(_06140_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15000_ (.A(_06141_),
    .B(_06142_),
    .CI(_06143_),
    .CO(_06138_),
    .S(_06144_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15001_ (.A(_06145_),
    .B(_06094_),
    .CI(_05974_),
    .CO(_06146_),
    .S(_06147_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15002_ (.A(_06148_),
    .B(_06149_),
    .CI(_06150_),
    .CO(_06151_),
    .S(_06152_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15003_ (.A(_05969_),
    .B(_06153_),
    .CI(_06154_),
    .CO(_06155_),
    .S(_06156_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15004_ (.A(_06157_),
    .B(_06158_),
    .CI(_06005_),
    .CO(_06159_),
    .S(_06160_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15005_ (.A(_06116_),
    .B(_06162_),
    .CI(_06163_),
    .CO(_06119_),
    .S(_06164_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15006_ (.A(_06159_),
    .B(_06165_),
    .CI(_06166_),
    .CO(_06162_),
    .S(_06167_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15007_ (.A(_05974_),
    .B(_05987_),
    .CI(_05997_),
    .CO(_06161_),
    .S(_06168_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15008_ (.A(_06170_),
    .B(_06171_),
    .CI(_06172_),
    .CO(_06173_),
    .S(_06174_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15009_ (.A(_06175_),
    .B(_06176_),
    .CI(_06177_),
    .CO(_06178_),
    .S(_06179_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15010_ (.A(_06126_),
    .B(_06180_),
    .CI(_06181_),
    .CO(_06182_),
    .S(_06183_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15011_ (.A(_06129_),
    .B(_06184_),
    .CI(_06185_),
    .CO(_06180_),
    .S(_06186_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15012_ (.A(_06132_),
    .B(_06187_),
    .CI(_06188_),
    .CO(_06184_),
    .S(_06189_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15013_ (.A(_06136_),
    .B(_06190_),
    .CI(_06191_),
    .CO(_06187_),
    .S(_06192_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15014_ (.A(_06140_),
    .B(_06194_),
    .CI(_06195_),
    .CO(_06190_),
    .S(_06196_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15015_ (.A(_06144_),
    .B(_06198_),
    .CI(_06199_),
    .CO(_06194_),
    .S(_06200_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15016_ (.A(_06201_),
    .B(_06202_),
    .CI(_06203_),
    .CO(_06198_),
    .S(_06204_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15017_ (.A(_06145_),
    .B(_06205_),
    .CI(_05987_),
    .CO(_06206_),
    .S(_06207_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15018_ (.A(_06208_),
    .B(_06209_),
    .CI(_06210_),
    .CO(_06211_),
    .S(_06212_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15019_ (.A(_05932_),
    .B(_06213_),
    .CI(_06214_),
    .CO(_06215_),
    .S(_06216_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15020_ (.A(_06217_),
    .B(_06218_),
    .CI(_06174_),
    .CO(_06219_),
    .S(_06220_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15021_ (.A(_06221_),
    .B(_06222_),
    .CI(_06223_),
    .CO(_06177_),
    .S(_06224_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15022_ (.A(_06011_),
    .B(_06169_),
    .CI(_06003_),
    .CO(_06218_),
    .S(_06225_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15023_ (.A(_06226_),
    .B(_06224_),
    .CI(_06227_),
    .CO(_06228_),
    .S(_06229_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15024_ (.A(_06186_),
    .B(_06230_),
    .CI(_06231_),
    .CO(_06232_),
    .S(_06233_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15025_ (.A(_06189_),
    .B(_06234_),
    .CI(_06235_),
    .CO(_06230_),
    .S(_06236_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15026_ (.A(_06192_),
    .B(_06237_),
    .CI(_06238_),
    .CO(_06234_),
    .S(_06239_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15027_ (.A(_06196_),
    .B(_06240_),
    .CI(_06241_),
    .CO(_06237_),
    .S(_06242_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15028_ (.A(_06200_),
    .B(_06244_),
    .CI(_06245_),
    .CO(_06240_),
    .S(_06246_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15029_ (.A(_06204_),
    .B(_06248_),
    .CI(_06249_),
    .CO(_06244_),
    .S(_06250_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15030_ (.A(_06251_),
    .B(_06252_),
    .CI(_06253_),
    .CO(_06248_),
    .S(_06254_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15031_ (.A(_06255_),
    .B(_06256_),
    .CI(_06169_),
    .CO(_06252_),
    .S(_06257_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15032_ (.A(_06258_),
    .B(_06259_),
    .CI(_06260_),
    .CO(_06261_),
    .S(_06262_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15033_ (.A(_06065_),
    .B(_06263_),
    .CI(_06264_),
    .CO(_06265_),
    .S(_06266_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15034_ (.A(_06225_),
    .B(_06267_),
    .CI(_06268_),
    .CO(_06269_),
    .S(_06270_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15035_ (.A(_06271_),
    .B(_06272_),
    .CI(_06273_),
    .CO(_06227_),
    .S(_06274_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15036_ (.A(_06275_),
    .B(_06276_),
    .CI(_06277_),
    .CO(_06278_),
    .S(_06279_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15037_ (.A(_06236_),
    .B(_06281_),
    .CI(_06282_),
    .CO(_06283_),
    .S(_06284_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15038_ (.A(_06239_),
    .B(_06285_),
    .CI(_06286_),
    .CO(_06281_),
    .S(_06287_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15039_ (.A(_06242_),
    .B(_06288_),
    .CI(_06279_),
    .CO(_06285_),
    .S(_06289_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15040_ (.A(_06246_),
    .B(_06290_),
    .CI(_06291_),
    .CO(_06288_),
    .S(_06292_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15041_ (.A(_06254_),
    .B(_06295_),
    .CI(_06296_),
    .CO(_06297_),
    .S(_06298_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15042_ (.A(_06257_),
    .B(_06300_),
    .CI(_06301_),
    .CO(_06295_),
    .S(_06302_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15043_ (.A(_06256_),
    .B(_06303_),
    .CI(_06003_),
    .CO(_06300_),
    .S(_06304_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15044_ (.A(_06305_),
    .B(_06306_),
    .CI(_06307_),
    .CO(_06308_),
    .S(_06309_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15045_ (.A(_06011_),
    .B(_06310_),
    .CI(_06311_),
    .CO(_06312_),
    .S(_06313_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15046_ (.A(_06169_),
    .B(_06003_),
    .CI(_06172_),
    .CO(_06267_),
    .S(_06314_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15047_ (.A(_06171_),
    .B(_06314_),
    .CI(_06315_),
    .CO(_06316_),
    .S(_06317_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15048_ (.A(_06318_),
    .B(_06319_),
    .CI(_06320_),
    .CO(_06321_),
    .S(_06322_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15049_ (.A(_06287_),
    .B(_06323_),
    .CI(_06324_),
    .CO(_06325_),
    .S(_06326_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15050_ (.A(_06289_),
    .B(_06327_),
    .CI(_06328_),
    .CO(_06323_),
    .S(_06329_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15051_ (.A(_06292_),
    .B(_06330_),
    .CI(_06322_),
    .CO(_06327_),
    .S(_06331_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15052_ (.A(_06333_),
    .B(_06334_),
    .CI(_06335_),
    .CO(_06332_),
    .S(_06336_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15053_ (.A(_06337_),
    .B(_06304_),
    .CI(_06338_),
    .CO(_06339_),
    .S(_06340_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15054_ (.A(_06343_),
    .B(_06344_),
    .CI(_06345_),
    .CO(_06346_),
    .S(_06347_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15055_ (.A(_05997_),
    .B(_06348_),
    .CI(_06349_),
    .CO(_06350_),
    .S(_06351_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15056_ (.A(_06003_),
    .B(_06172_),
    .CI(_06352_),
    .CO(_06315_),
    .S(_06353_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15057_ (.A(_06354_),
    .B(_06355_),
    .CI(_06356_),
    .CO(_06357_),
    .S(_06358_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15058_ (.A(_06329_),
    .B(_06359_),
    .CI(_06360_),
    .CO(_06361_),
    .S(_06362_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15059_ (.A(_06331_),
    .B(_06363_),
    .CI(_06364_),
    .CO(_06359_),
    .S(_06365_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15060_ (.A(_06366_),
    .B(_06367_),
    .CI(_06358_),
    .CO(_06363_),
    .S(_06368_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15061_ (.A(_06370_),
    .B(_06371_),
    .CI(_06372_),
    .CO(_06369_),
    .S(_06373_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15062_ (.A(_06374_),
    .B(_06375_),
    .CI(_06376_),
    .CO(_06377_),
    .S(_06378_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15063_ (.A(_06381_),
    .B(_06382_),
    .CI(_06383_),
    .CO(_06384_),
    .S(_06385_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15064_ (.A(_06365_),
    .B(_06386_),
    .CI(_06387_),
    .CO(_06388_),
    .S(_06389_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15065_ (.A(_06368_),
    .B(_06390_),
    .CI(_06391_),
    .CO(_06386_),
    .S(_06392_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15066_ (.A(_06393_),
    .B(_06394_),
    .CI(_06385_),
    .CO(_06390_),
    .S(_06395_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15067_ (.A(_06397_),
    .B(_06398_),
    .CI(_06399_),
    .CO(_06400_),
    .S(_06401_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15068_ (.A(_06404_),
    .B(_06405_),
    .CI(_06406_),
    .CO(_06407_),
    .S(_06408_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15069_ (.A(_06392_),
    .B(_06409_),
    .CI(_06410_),
    .CO(_06411_),
    .S(_06412_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15070_ (.A(_06395_),
    .B(_06413_),
    .CI(_06414_),
    .CO(_06409_),
    .S(_06415_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15071_ (.A(_06416_),
    .B(_06417_),
    .CI(_06418_),
    .CO(_06413_),
    .S(_06419_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15072_ (.A(_06337_),
    .B(_06422_),
    .CI(_06423_),
    .CO(_06424_),
    .S(_06425_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15073_ (.A(_06428_),
    .B(_06429_),
    .CI(_06430_),
    .CO(_06431_),
    .S(_06432_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15074_ (.A(_06435_),
    .B(_06436_),
    .CI(_06437_),
    .CO(_06438_),
    .S(_06439_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15075_ (.A(_06415_),
    .B(_06440_),
    .CI(_06441_),
    .CO(_06442_),
    .S(_06443_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15076_ (.A(_06419_),
    .B(_06444_),
    .CI(_06445_),
    .CO(_06440_),
    .S(_06446_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15077_ (.A(_06447_),
    .B(_06448_),
    .CI(_06449_),
    .CO(_06444_),
    .S(_06450_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15078_ (.A(_06205_),
    .B(_06451_),
    .CI(_06452_),
    .CO(_06453_),
    .S(_06454_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15079_ (.A(_06446_),
    .B(_06455_),
    .CI(_06456_),
    .CO(_06457_),
    .S(_06458_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15080_ (.A(_06450_),
    .B(_06459_),
    .CI(_06453_),
    .CO(_06455_),
    .S(_06460_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15081_ (.A(_06462_),
    .B(_06463_),
    .CI(_06464_),
    .CO(_06461_),
    .S(_06465_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15082_ (.A(_06299_),
    .B(_06467_),
    .CI(_06468_),
    .CO(_06469_),
    .S(_06470_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15083_ (.A(_06471_),
    .B(_06472_),
    .CI(_06473_),
    .CO(_06474_),
    .S(_06475_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15084_ (.A(_06460_),
    .B(_06478_),
    .CI(_06479_),
    .CO(_06480_),
    .S(_06481_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15085_ (.A(_06482_),
    .B(_06483_),
    .CI(_06484_),
    .CO(_06478_),
    .S(_06485_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15086_ (.A(_06485_),
    .B(_06487_),
    .CI(_06488_),
    .CO(_06489_),
    .S(_06490_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15087_ (.A(_06491_),
    .B(_06492_),
    .CI(_06493_),
    .CO(_06494_),
    .S(_06495_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15088_ (.A(_06496_),
    .B(_06497_),
    .CI(_06498_),
    .CO(_06499_),
    .S(_06500_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15089_ (.A(_06501_),
    .B(_06497_),
    .CI(_06502_),
    .CO(_06503_),
    .S(_06504_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15090_ (.A(_06505_),
    .B(_06506_),
    .CI(_06507_),
    .CO(_06508_),
    .S(_06509_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15091_ (.A(_06510_),
    .B(_06511_),
    .CI(_06512_),
    .CO(_06513_),
    .S(_06514_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15092_ (.A(_06515_),
    .B(_06516_),
    .CI(_06517_),
    .CO(_06518_),
    .S(_06519_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15093_ (.A(_06520_),
    .B(_06521_),
    .CI(_06522_),
    .CO(_06523_),
    .S(_06524_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15094_ (.A(_06516_),
    .B(_06517_),
    .CI(_06525_),
    .CO(_06526_),
    .S(_06527_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15095_ (.A(_06528_),
    .B(_06529_),
    .CI(_06530_),
    .CO(_06531_),
    .S(_06532_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15096_ (.A(_06533_),
    .B(_06534_),
    .CI(_06535_),
    .CO(_06512_),
    .S(_06536_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15097_ (.A(_06537_),
    .B(_06538_),
    .CI(_06539_),
    .CO(_06540_),
    .S(_06541_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15098_ (.A(_06542_),
    .B(_06543_),
    .CI(_06527_),
    .CO(_06544_),
    .S(_06545_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15099_ (.A(_06546_),
    .B(_06547_),
    .CI(_06521_),
    .CO(_06548_),
    .S(_06549_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15100_ (.A(_06550_),
    .B(_06551_),
    .CI(_06552_),
    .CO(_06553_),
    .S(_06554_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15101_ (.A(_06518_),
    .B(_06555_),
    .CI(_06556_),
    .CO(_06557_),
    .S(_06558_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15102_ (.A(_06559_),
    .B(_06560_),
    .CI(_06554_),
    .CO(_06561_),
    .S(_06562_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15103_ (.A(_06563_),
    .B(_06564_),
    .CI(_06541_),
    .CO(_06565_),
    .S(_06566_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15104_ (.A(_06567_),
    .B(_06568_),
    .CI(_06569_),
    .CO(_06570_),
    .S(_06571_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15105_ (.A(_06572_),
    .B(_06573_),
    .CI(_06519_),
    .CO(_06574_),
    .S(_06575_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15106_ (.A(_06577_),
    .B(_06578_),
    .CI(_06547_),
    .CO(_06576_),
    .S(_06579_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15107_ (.A(_06521_),
    .B(_06522_),
    .CI(_06580_),
    .CO(_06581_),
    .S(_06582_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15108_ (.A(_06583_),
    .B(_06575_),
    .CI(_06584_),
    .CO(_06585_),
    .S(_06586_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15109_ (.A(_06558_),
    .B(_06587_),
    .CI(_06588_),
    .CO(_06589_),
    .S(_06590_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15110_ (.A(_06591_),
    .B(_06592_),
    .CI(_06593_),
    .CO(_06587_),
    .S(_06594_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15111_ (.A(_06595_),
    .B(_06596_),
    .CI(_06597_),
    .CO(_06598_),
    .S(_06599_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15112_ (.A(_06600_),
    .B(_06601_),
    .CI(_06602_),
    .CO(_06603_),
    .S(_06604_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15113_ (.A(_06606_),
    .B(_06607_),
    .CI(_06608_),
    .CO(_06609_),
    .S(_06610_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15114_ (.A(_06611_),
    .B(_06612_),
    .CI(_06613_),
    .CO(_06614_),
    .S(_06615_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15115_ (.A(_06601_),
    .B(_06618_),
    .CI(_06602_),
    .CO(_06617_),
    .S(_06619_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15116_ (.A(_06562_),
    .B(_06620_),
    .CI(_06599_),
    .CO(_06621_),
    .S(_06622_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15117_ (.A(_06623_),
    .B(_06624_),
    .CI(_06625_),
    .CO(_06620_),
    .S(_06626_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15118_ (.A(_06627_),
    .B(_06628_),
    .CI(_06629_),
    .CO(_06624_),
    .S(_06630_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15119_ (.A(_06631_),
    .B(_06632_),
    .CI(_06535_),
    .CO(_06633_),
    .S(_06634_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15120_ (.A(_06635_),
    .B(_06636_),
    .CI(_06582_),
    .CO(_06584_),
    .S(_06637_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15121_ (.A(_06533_),
    .B(_06534_),
    .CI(_06578_),
    .CO(_06638_),
    .S(_06639_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15122_ (.A(_06547_),
    .B(_06521_),
    .CI(_06522_),
    .CO(_06640_),
    .S(_06641_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15123_ (.A(_06642_),
    .B(_06637_),
    .CI(_06643_),
    .CO(_06644_),
    .S(_06645_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15124_ (.A(_06594_),
    .B(_06646_),
    .CI(_06647_),
    .CO(_06648_),
    .S(_06649_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15125_ (.A(_06650_),
    .B(_06651_),
    .CI(_06652_),
    .CO(_06646_),
    .S(_06653_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15126_ (.A(_06654_),
    .B(_06655_),
    .CI(_06656_),
    .CO(_06657_),
    .S(_06658_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15127_ (.A(_06610_),
    .B(_06659_),
    .CI(_06660_),
    .CO(_06661_),
    .S(_06662_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15128_ (.A(_06663_),
    .B(_06619_),
    .CI(_06664_),
    .CO(_06665_),
    .S(_06666_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15129_ (.A(_06667_),
    .B(_06668_),
    .CI(_06605_),
    .CO(_06669_),
    .S(_06670_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15130_ (.A(_06657_),
    .B(_06662_),
    .CI(_06671_),
    .CO(_06672_),
    .S(_06673_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15131_ (.A(_06622_),
    .B(_06674_),
    .CI(_06673_),
    .CO(_06675_),
    .S(_06676_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15132_ (.A(_06626_),
    .B(_06677_),
    .CI(_06658_),
    .CO(_06674_),
    .S(_06678_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15133_ (.A(_06679_),
    .B(_06680_),
    .CI(_06645_),
    .CO(_06681_),
    .S(_06682_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15134_ (.A(_06501_),
    .B(_06683_),
    .CI(_06502_),
    .CO(_06684_),
    .S(_06685_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15135_ (.A(_06686_),
    .B(_06687_),
    .CI(_06641_),
    .CO(_06643_),
    .S(_06688_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15136_ (.A(_06568_),
    .B(_06534_),
    .CI(_06569_),
    .CO(_06689_),
    .S(_06690_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15137_ (.A(_06507_),
    .B(_06691_),
    .CI(_06692_),
    .CO(_06693_),
    .S(_06694_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15138_ (.A(_06695_),
    .B(_06688_),
    .CI(_06696_),
    .CO(_06697_),
    .S(_06698_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15139_ (.A(_06699_),
    .B(_06653_),
    .CI(_06700_),
    .CO(_06701_),
    .S(_06702_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15140_ (.A(_06693_),
    .B(_06703_),
    .CI(_06704_),
    .CO(_06700_),
    .S(_06705_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15141_ (.A(_06706_),
    .B(_06707_),
    .CI(_06708_),
    .CO(_06709_),
    .S(_06710_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15142_ (.A(_06711_),
    .B(_06712_),
    .CI(_06713_),
    .CO(_06671_),
    .S(_06714_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15143_ (.A(_06601_),
    .B(_06715_),
    .CI(_06716_),
    .CO(_06717_),
    .S(_06718_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15144_ (.A(_06667_),
    .B(_06668_),
    .CI(_06719_),
    .CO(_06720_),
    .S(_06721_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15145_ (.A(_06709_),
    .B(_06714_),
    .CI(_06722_),
    .CO(_06723_),
    .S(_06724_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15146_ (.A(_06725_),
    .B(_06726_),
    .CI(_06727_),
    .CO(_06728_),
    .S(_06729_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15147_ (.A(_06678_),
    .B(_06731_),
    .CI(_06724_),
    .CO(_06730_),
    .S(_06732_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15148_ (.A(_06733_),
    .B(_06734_),
    .CI(_06710_),
    .CO(_06731_),
    .S(_06735_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15149_ (.A(_06736_),
    .B(_06737_),
    .CI(_06698_),
    .CO(_06738_),
    .S(_06739_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15150_ (.A(_06740_),
    .B(_06741_),
    .CI(_06694_),
    .CO(_06696_),
    .S(_06742_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15151_ (.A(_06632_),
    .B(_06569_),
    .CI(_06535_),
    .CO(_06743_),
    .S(_06744_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15152_ (.A(_06745_),
    .B(_06507_),
    .CI(_06691_),
    .CO(_06746_),
    .S(_06747_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15153_ (.A(_06748_),
    .B(_06705_),
    .CI(_06749_),
    .CO(_06750_),
    .S(_06751_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15154_ (.A(_06746_),
    .B(_06752_),
    .CI(_06753_),
    .CO(_06749_),
    .S(_06754_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15155_ (.A(_06755_),
    .B(_06751_),
    .CI(_06756_),
    .CO(_06757_),
    .S(_06758_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15156_ (.A(_06759_),
    .B(_06760_),
    .CI(_06761_),
    .CO(_06722_),
    .S(_06762_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15157_ (.A(_06602_),
    .B(_06763_),
    .CI(_06764_),
    .CO(_06765_),
    .S(_06766_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15158_ (.A(_06767_),
    .B(_06667_),
    .CI(_06719_),
    .CO(_06768_),
    .S(_06769_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15159_ (.A(_06770_),
    .B(_06762_),
    .CI(_06771_),
    .CO(_06772_),
    .S(_06773_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15160_ (.A(_06729_),
    .B(_06774_),
    .CI(_06775_),
    .CO(_06776_),
    .S(_06777_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15161_ (.A(_06778_),
    .B(_06779_),
    .CI(_06780_),
    .CO(_06774_),
    .S(_06781_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15162_ (.A(_06735_),
    .B(_06783_),
    .CI(_06773_),
    .CO(_06782_),
    .S(_06784_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15163_ (.A(_06785_),
    .B(_06786_),
    .CI(_06787_),
    .CO(_06783_),
    .S(_06788_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15164_ (.A(_06789_),
    .B(_06790_),
    .CI(_06791_),
    .CO(_06792_),
    .S(_06793_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15165_ (.A(_06794_),
    .B(_06795_),
    .CI(_06747_),
    .CO(_06796_),
    .S(_06797_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15166_ (.A(_06799_),
    .B(_06567_),
    .CI(_06535_),
    .CO(_06798_),
    .S(_06800_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15167_ (.A(_06534_),
    .B(_06569_),
    .CI(_06578_),
    .CO(_06801_),
    .S(_06802_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15168_ (.A(_06803_),
    .B(_06754_),
    .CI(_06804_),
    .CO(_06756_),
    .S(_06805_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15169_ (.A(_06806_),
    .B(_06807_),
    .CI(_06808_),
    .CO(_06804_),
    .S(_06809_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15170_ (.A(_06810_),
    .B(_06811_),
    .CI(_06812_),
    .CO(_06813_),
    .S(_06814_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15171_ (.A(_06815_),
    .B(_06816_),
    .CI(_06817_),
    .CO(_06771_),
    .S(_06818_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15172_ (.A(_06618_),
    .B(_06819_),
    .CI(_06820_),
    .CO(_06821_),
    .S(_06822_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15173_ (.A(_06823_),
    .B(_06767_),
    .CI(_06719_),
    .CO(_06824_),
    .S(_06825_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15174_ (.A(_06826_),
    .B(_06827_),
    .CI(_06828_),
    .CO(_06829_),
    .S(_06830_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15175_ (.A(_06781_),
    .B(_06831_),
    .CI(_06832_),
    .CO(_06833_),
    .S(_06834_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15176_ (.A(_06835_),
    .B(_06836_),
    .CI(_06837_),
    .CO(_06831_),
    .S(_06838_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15177_ (.A(_06788_),
    .B(_06840_),
    .CI(_06841_),
    .CO(_06839_),
    .S(_06842_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _15178_ (.A(_06843_),
    .B(_06844_),
    .CI(_06814_),
    .CO(_06840_),
    .S(_06845_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15179_ (.A(_06846_),
    .B(_06847_),
    .CI(_06848_),
    .CO(_06844_),
    .S(_06849_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15180_ (.A(_06850_),
    .B(_06851_),
    .CI(_06852_),
    .CO(_06853_),
    .S(_06854_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15181_ (.A(_06856_),
    .B(_06567_),
    .CI(_06631_),
    .CO(_06855_),
    .S(_06857_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15182_ (.A(_06534_),
    .B(_06569_),
    .CI(_06535_),
    .CO(_06858_),
    .S(_06859_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15183_ (.A(_06860_),
    .B(_06861_),
    .CI(_06862_),
    .CO(_06863_),
    .S(_06864_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15184_ (.A(_06865_),
    .B(_06866_),
    .CI(_06867_),
    .CO(_06868_),
    .S(_06869_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15185_ (.A(_06667_),
    .B(_06825_),
    .CI(_06870_),
    .CO(_06871_),
    .S(_06872_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15186_ (.A(_06823_),
    .B(_06873_),
    .CI(_06767_),
    .CO(_06870_),
    .S(_06874_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15187_ (.A(_06875_),
    .B(_06876_),
    .CI(_06877_),
    .CO(_06878_),
    .S(_06879_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15188_ (.A(_06838_),
    .B(_06880_),
    .CI(_06881_),
    .CO(_06882_),
    .S(_06883_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15189_ (.A(_06884_),
    .B(_06885_),
    .CI(_06886_),
    .CO(_06880_),
    .S(_06887_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15190_ (.A(_06845_),
    .B(_06889_),
    .CI(_06890_),
    .CO(_06888_),
    .S(_06891_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15191_ (.A(_06892_),
    .B(_06893_),
    .CI(_06894_),
    .CO(_06895_),
    .S(_06896_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15192_ (.A(_06857_),
    .B(_06897_),
    .CI(_06859_),
    .CO(_06898_),
    .S(_06899_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15193_ (.A(_06567_),
    .B(_06569_),
    .CI(_06535_),
    .CO(_06901_),
    .S(_06902_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15194_ (.A(_06903_),
    .B(_06904_),
    .CI(_06905_),
    .CO(_06906_),
    .S(_06907_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15195_ (.A(_06908_),
    .B(_06909_),
    .CI(_06910_),
    .CO(_06911_),
    .S(_06912_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15196_ (.A(_06913_),
    .B(_06914_),
    .CI(_06915_),
    .CO(_06916_),
    .S(_06917_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15197_ (.A(_06918_),
    .B(_06823_),
    .CI(_06873_),
    .CO(_06919_),
    .S(_06920_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15198_ (.A(_06921_),
    .B(_06922_),
    .CI(_06923_),
    .CO(_06924_),
    .S(_06925_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15199_ (.A(_06887_),
    .B(_06926_),
    .CI(_06927_),
    .CO(_06928_),
    .S(_06929_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15200_ (.A(_06930_),
    .B(_06931_),
    .CI(_06932_),
    .CO(_06926_),
    .S(_06933_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15201_ (.A(_06935_),
    .B(_06936_),
    .CI(_06937_),
    .CO(_06934_),
    .S(_06938_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15202_ (.A(_06939_),
    .B(_06940_),
    .CI(_06941_),
    .CO(_06942_),
    .S(_06943_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15203_ (.A(_06567_),
    .B(_06631_),
    .CI(_06535_),
    .CO(_06944_),
    .S(_06945_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15204_ (.A(_06946_),
    .B(_06947_),
    .CI(_06948_),
    .CO(_06949_),
    .S(_06950_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15205_ (.A(_06951_),
    .B(_06952_),
    .CI(_06953_),
    .CO(_06954_),
    .S(_06955_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15206_ (.A(_06956_),
    .B(_06957_),
    .CI(_06958_),
    .CO(_06959_),
    .S(_06960_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15207_ (.A(_06699_),
    .B(_06748_),
    .CI(_06961_),
    .CO(_06958_),
    .S(_06962_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15208_ (.A(_06963_),
    .B(_06964_),
    .CI(_06965_),
    .CO(_06966_),
    .S(_06967_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15209_ (.A(_06933_),
    .B(_06968_),
    .CI(_06969_),
    .CO(_06970_),
    .S(_06971_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15210_ (.A(_06972_),
    .B(_06973_),
    .CI(_06974_),
    .CO(_06968_),
    .S(_06975_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15211_ (.A(_06977_),
    .B(_06978_),
    .CI(_06979_),
    .CO(_06976_),
    .S(_06980_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15212_ (.A(_06981_),
    .B(_06982_),
    .CI(_06983_),
    .CO(_06984_),
    .S(_06985_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15213_ (.A(_06986_),
    .B(_06987_),
    .CI(_06988_),
    .CO(_06989_),
    .S(_06990_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15214_ (.A(_06823_),
    .B(_06991_),
    .CI(_06992_),
    .CO(_06993_),
    .S(_06994_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15215_ (.A(_06699_),
    .B(_06748_),
    .CI(_06803_),
    .CO(_06995_),
    .S(_06996_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15216_ (.A(_06997_),
    .B(_06998_),
    .CI(_06999_),
    .CO(_07000_),
    .S(_07001_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15217_ (.A(_06975_),
    .B(_07002_),
    .CI(_07003_),
    .CO(_07004_),
    .S(_07005_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15218_ (.A(_07006_),
    .B(_07007_),
    .CI(_07008_),
    .CO(_07002_),
    .S(_07009_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15219_ (.A(_06985_),
    .B(_07010_),
    .CI(_07011_),
    .CO(_07007_),
    .S(_07012_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15220_ (.A(_07013_),
    .B(_07014_),
    .CI(_07015_),
    .CO(_07010_),
    .S(_07016_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15221_ (.A(_06683_),
    .B(_06496_),
    .CI(_06502_),
    .CO(_06986_),
    .S(_07017_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15222_ (.A(_06897_),
    .B(_07018_),
    .CI(_07019_),
    .CO(_07020_),
    .S(_07021_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15223_ (.A(_07009_),
    .B(_07022_),
    .CI(_07023_),
    .CO(_07024_),
    .S(_07025_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15224_ (.A(_07012_),
    .B(_07026_),
    .CI(_07027_),
    .CO(_07022_),
    .S(_07028_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15225_ (.A(_07016_),
    .B(_07029_),
    .CI(_07030_),
    .CO(_07026_),
    .S(_07031_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15226_ (.A(_07032_),
    .B(_07033_),
    .CI(_07034_),
    .CO(_07029_),
    .S(_07035_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15227_ (.A(_06961_),
    .B(_07036_),
    .CI(_06996_),
    .CO(_07037_),
    .S(_07038_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15228_ (.A(_07039_),
    .B(_07040_),
    .CI(_07041_),
    .CO(_07042_),
    .S(_07043_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15229_ (.A(_07028_),
    .B(_07044_),
    .CI(_07045_),
    .CO(_07046_),
    .S(_07047_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15230_ (.A(_07031_),
    .B(_07048_),
    .CI(_07049_),
    .CO(_07044_),
    .S(_07050_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15231_ (.A(_07035_),
    .B(_07051_),
    .CI(_07052_),
    .CO(_07048_),
    .S(_07053_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15232_ (.A(_07054_),
    .B(_07055_),
    .CI(_07056_),
    .CO(_07051_),
    .S(_07057_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15233_ (.A(_07058_),
    .B(_07053_),
    .CI(_07059_),
    .CO(_07060_),
    .S(_07061_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15234_ (.A(_07057_),
    .B(_07062_),
    .CI(_07063_),
    .CO(_07059_),
    .S(_07064_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15235_ (.A(_07066_),
    .B(_07067_),
    .CI(_07068_),
    .CO(_07065_),
    .S(_07069_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _15236_ (.A(_07069_),
    .B(_07070_),
    .CI(_07071_),
    .CO(_07072_),
    .S(_07073_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15237_ (.A(_07076_),
    .B(net369),
    .CO(_07077_),
    .S(_07078_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15238_ (.A(_05862_),
    .B(_07079_),
    .CO(_07080_),
    .S(_07081_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15239_ (.A(_07082_),
    .B(_07083_),
    .CO(_07084_),
    .S(_07085_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15240_ (.A(_05862_),
    .B(_07086_),
    .CO(_07087_),
    .S(_07088_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15241_ (.A(_07076_),
    .B(net342),
    .CO(_07089_),
    .S(_07090_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15242_ (.A(_07092_),
    .B(_07091_),
    .CO(_07093_),
    .S(_07094_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15243_ (.A(_07095_),
    .B(_07082_),
    .CO(_07096_),
    .S(_07097_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15244_ (.A(_05862_),
    .B(_07098_),
    .CO(_07099_),
    .S(_07100_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15245_ (.A(_07076_),
    .B(net343),
    .CO(_07101_),
    .S(_07102_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15246_ (.A(_07104_),
    .B(_07103_),
    .CO(_07105_),
    .S(_07106_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15247_ (.A(_07091_),
    .B(_07107_),
    .CO(_07108_),
    .S(_07109_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15248_ (.A(_07082_),
    .B(_07110_),
    .CO(_07111_),
    .S(_07112_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15249_ (.A(_05862_),
    .B(_07113_),
    .CO(_07114_),
    .S(_07115_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15250_ (.A(_07076_),
    .B(net344),
    .CO(_07116_),
    .S(_07117_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15251_ (.A(_05862_),
    .B(_07118_),
    .CO(_07119_),
    .S(_07120_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15252_ (.A(_07076_),
    .B(net345),
    .CO(_07121_),
    .S(_07122_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15253_ (.A(_07123_),
    .B(_07124_),
    .CO(_07125_),
    .S(_07126_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15254_ (.A(_07127_),
    .B(_07103_),
    .CO(_07128_),
    .S(_07129_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15255_ (.A(_07091_),
    .B(_07130_),
    .CO(_07131_),
    .S(_07132_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15256_ (.A(_07082_),
    .B(_07133_),
    .CO(_07134_),
    .S(_07135_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15257_ (.A(_07136_),
    .B(_07137_),
    .CO(_07138_),
    .S(_07139_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15258_ (.A(_07123_),
    .B(_07140_),
    .CO(_07141_),
    .S(_07142_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15259_ (.A(_07143_),
    .B(_07103_),
    .CO(_07144_),
    .S(_07145_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15260_ (.A(_07091_),
    .B(_07146_),
    .CO(_07147_),
    .S(_07148_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15261_ (.A(_07082_),
    .B(_07149_),
    .CO(_07150_),
    .S(_07151_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15262_ (.A(_05862_),
    .B(_07152_),
    .CO(_07153_),
    .S(_07154_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15263_ (.A(_07076_),
    .B(net346),
    .CO(_07155_),
    .S(_07156_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15264_ (.A(_07157_),
    .B(_07136_),
    .CO(_07158_),
    .S(_07159_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15265_ (.A(_07160_),
    .B(_07123_),
    .CO(_07161_),
    .S(_07162_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15266_ (.A(_07103_),
    .B(_07163_),
    .CO(_07164_),
    .S(_07165_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15267_ (.A(_07091_),
    .B(_07166_),
    .CO(_07167_),
    .S(_07168_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15268_ (.A(_07082_),
    .B(_07169_),
    .CO(_07170_),
    .S(_07171_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15269_ (.A(_05862_),
    .B(_07172_),
    .CO(_07173_),
    .S(_07174_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15270_ (.A(_07076_),
    .B(net347),
    .CO(_07175_),
    .S(_07176_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15271_ (.A(_07177_),
    .B(_07178_),
    .CO(_07179_),
    .S(_07180_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15272_ (.A(_07136_),
    .B(_07181_),
    .CO(_07182_),
    .S(_07183_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15273_ (.A(_07123_),
    .B(_07184_),
    .CO(_07185_),
    .S(_07186_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15274_ (.A(net19),
    .B(_07187_),
    .CO(_07188_),
    .S(_07189_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15275_ (.A(_07091_),
    .B(_07190_),
    .CO(_07191_),
    .S(_07192_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15276_ (.A(_07082_),
    .B(_07193_),
    .CO(_07194_),
    .S(_07195_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15277_ (.A(_05862_),
    .B(_07196_),
    .CO(_07197_),
    .S(_07198_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15278_ (.A(_07076_),
    .B(net348),
    .CO(_07199_),
    .S(_07200_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15279_ (.A(_07136_),
    .B(_07201_),
    .CO(_07202_),
    .S(_07203_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15280_ (.A(_07123_),
    .B(_07204_),
    .CO(_07205_),
    .S(_07206_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15281_ (.A(_07207_),
    .B(net19),
    .CO(_07208_),
    .S(_07209_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15282_ (.A(_07091_),
    .B(_07210_),
    .CO(_07211_),
    .S(_07212_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15283_ (.A(_07082_),
    .B(_07213_),
    .CO(_07214_),
    .S(_07215_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15284_ (.A(_05862_),
    .B(_07216_),
    .CO(_07217_),
    .S(_07218_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15285_ (.A(net8),
    .B(net349),
    .CO(_07219_),
    .S(_07220_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15286_ (.A(_07136_),
    .B(_07221_),
    .CO(_07222_),
    .S(_07223_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15287_ (.A(_07123_),
    .B(_07224_),
    .CO(_07225_),
    .S(_07226_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15288_ (.A(net19),
    .B(_07227_),
    .CO(_07228_),
    .S(_07229_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15289_ (.A(_07230_),
    .B(_07082_),
    .CO(_07231_),
    .S(_07232_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15290_ (.A(_07233_),
    .B(_05862_),
    .CO(_07234_),
    .S(_07235_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15291_ (.A(net8),
    .B(net350),
    .CO(_07236_),
    .S(_07237_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15292_ (.A(_07091_),
    .B(_07238_),
    .CO(_07239_),
    .S(_07240_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15293_ (.A(_07136_),
    .B(_07241_),
    .CO(_07242_),
    .S(_07243_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15294_ (.A(_07123_),
    .B(_07244_),
    .CO(_07245_),
    .S(_07246_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15295_ (.A(net19),
    .B(_07247_),
    .CO(_07248_),
    .S(_07249_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15296_ (.A(_07091_),
    .B(_07250_),
    .CO(_07251_),
    .S(_07252_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15297_ (.A(_07082_),
    .B(_07253_),
    .CO(_07254_),
    .S(_07255_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15298_ (.A(_05862_),
    .B(_07256_),
    .CO(_07257_),
    .S(_07258_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15299_ (.A(net8),
    .B(net351),
    .CO(_07259_),
    .S(_07260_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15300_ (.A(_07082_),
    .B(_07261_),
    .CO(_07262_),
    .S(_07263_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15301_ (.A(_05862_),
    .B(_07264_),
    .CO(_07265_),
    .S(_07266_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15302_ (.A(net19),
    .B(_07267_),
    .CO(_07268_),
    .S(_07269_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15303_ (.A(_07091_),
    .B(_07270_),
    .CO(_07271_),
    .S(_07272_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15304_ (.A(net8),
    .B(net352),
    .CO(_07273_),
    .S(_07274_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15305_ (.A(_07136_),
    .B(_07275_),
    .CO(_07276_),
    .S(_07277_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15306_ (.A(_07123_),
    .B(_07278_),
    .CO(_07279_),
    .S(_07280_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15307_ (.A(_07136_),
    .B(_07281_),
    .CO(_07282_),
    .S(_07283_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15308_ (.A(_07123_),
    .B(_07284_),
    .CO(_07285_),
    .S(_07286_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15309_ (.A(net19),
    .B(_07287_),
    .CO(_07288_),
    .S(_07289_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15310_ (.A(_07091_),
    .B(_07290_),
    .CO(_07291_),
    .S(_07292_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15311_ (.A(_07082_),
    .B(_07293_),
    .CO(_07294_),
    .S(_07295_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15312_ (.A(_05862_),
    .B(_07296_),
    .CO(_07297_),
    .S(_07298_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15313_ (.A(net8),
    .B(net353),
    .CO(_07299_),
    .S(_07300_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15314_ (.A(_07136_),
    .B(_07301_),
    .CO(_07302_),
    .S(_07303_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15315_ (.A(_07123_),
    .B(_07304_),
    .CO(_07305_),
    .S(_07306_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15316_ (.A(net19),
    .B(_07307_),
    .CO(_07308_),
    .S(_07309_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15317_ (.A(_07091_),
    .B(_07310_),
    .CO(_07311_),
    .S(_07312_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15318_ (.A(_07082_),
    .B(_07313_),
    .CO(_07314_),
    .S(_07315_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15319_ (.A(_05862_),
    .B(_07316_),
    .CO(_07317_),
    .S(_07318_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15320_ (.A(net8),
    .B(net354),
    .CO(_07319_),
    .S(_07320_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15321_ (.A(_07136_),
    .B(_07321_),
    .CO(_07322_),
    .S(_07323_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15322_ (.A(_07123_),
    .B(_07324_),
    .CO(_07325_),
    .S(_07326_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15323_ (.A(net19),
    .B(_07327_),
    .CO(_07328_),
    .S(_07329_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15324_ (.A(_07091_),
    .B(_07330_),
    .CO(_07331_),
    .S(_07332_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15325_ (.A(_07082_),
    .B(_07333_),
    .CO(_07334_),
    .S(_07335_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15326_ (.A(_05862_),
    .B(_07336_),
    .CO(_07337_),
    .S(_07338_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15327_ (.A(net8),
    .B(net355),
    .CO(_07339_),
    .S(_07340_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15328_ (.A(net8),
    .B(net356),
    .CO(_07341_),
    .S(_07342_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15329_ (.A(_07136_),
    .B(_07343_),
    .CO(_07344_),
    .S(_07345_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15330_ (.A(_07123_),
    .B(_07346_),
    .CO(_07347_),
    .S(_07348_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15331_ (.A(net2),
    .B(_07349_),
    .CO(_07350_),
    .S(_07351_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15332_ (.A(_07091_),
    .B(_07352_),
    .CO(_07353_),
    .S(_07354_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15333_ (.A(_07082_),
    .B(_07355_),
    .CO(_07356_),
    .S(_07357_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15334_ (.A(_05862_),
    .B(_07358_),
    .CO(_07359_),
    .S(_07360_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15335_ (.A(_05862_),
    .B(_07361_),
    .CO(_07362_),
    .S(_07363_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15336_ (.A(net1),
    .B(net357),
    .CO(_07364_),
    .S(_07365_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15337_ (.A(_07136_),
    .B(_07366_),
    .CO(_07367_),
    .S(_07368_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15338_ (.A(_07123_),
    .B(_07369_),
    .CO(_07370_),
    .S(_07371_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15339_ (.A(net2),
    .B(_07372_),
    .CO(_07373_),
    .S(_07374_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15340_ (.A(_07091_),
    .B(_07375_),
    .CO(_07376_),
    .S(_07377_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15341_ (.A(_07082_),
    .B(_07378_),
    .CO(_07379_),
    .S(_07380_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15342_ (.A(_07082_),
    .B(_07381_),
    .CO(_07382_),
    .S(_07383_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15343_ (.A(_05862_),
    .B(_07384_),
    .CO(_07385_),
    .S(_07386_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15344_ (.A(net1),
    .B(net358),
    .CO(_07387_),
    .S(_07388_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15345_ (.A(_07136_),
    .B(_07389_),
    .CO(_07390_),
    .S(_07391_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15346_ (.A(_07123_),
    .B(_07392_),
    .CO(_07393_),
    .S(_07394_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15347_ (.A(net2),
    .B(_07395_),
    .CO(_07396_),
    .S(_07397_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15348_ (.A(_07091_),
    .B(_07398_),
    .CO(_07399_),
    .S(_07400_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15349_ (.A(_07091_),
    .B(_07401_),
    .CO(_07402_),
    .S(_07403_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15350_ (.A(_07082_),
    .B(_07404_),
    .CO(_07405_),
    .S(_07406_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15351_ (.A(_05862_),
    .B(_07407_),
    .CO(_07408_),
    .S(_07409_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15352_ (.A(net1),
    .B(net359),
    .CO(_07410_),
    .S(_07411_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15353_ (.A(_07136_),
    .B(_07412_),
    .CO(_07413_),
    .S(_07414_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15354_ (.A(_07123_),
    .B(_07415_),
    .CO(_07416_),
    .S(_07417_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15355_ (.A(net2),
    .B(_07418_),
    .CO(_07419_),
    .S(_07420_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15356_ (.A(net2),
    .B(_07421_),
    .CO(_07422_),
    .S(_07423_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15357_ (.A(_07091_),
    .B(_07424_),
    .CO(_07425_),
    .S(_07426_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15358_ (.A(_07082_),
    .B(_07427_),
    .CO(_07428_),
    .S(_07429_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15359_ (.A(_05862_),
    .B(_07430_),
    .CO(_07431_),
    .S(_07432_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15360_ (.A(net1),
    .B(net360),
    .CO(_07433_),
    .S(_07434_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15361_ (.A(_07136_),
    .B(_07435_),
    .CO(_07436_),
    .S(_07437_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15362_ (.A(_07123_),
    .B(_07438_),
    .CO(_07439_),
    .S(_07440_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15363_ (.A(_07123_),
    .B(_07441_),
    .CO(_07442_),
    .S(_07443_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15364_ (.A(net2),
    .B(_07444_),
    .CO(_07445_),
    .S(_07446_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15365_ (.A(_07091_),
    .B(_07447_),
    .CO(_07448_),
    .S(_07449_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15366_ (.A(_07082_),
    .B(_07450_),
    .CO(_07451_),
    .S(_07452_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15367_ (.A(_05862_),
    .B(_07453_),
    .CO(_07454_),
    .S(_07455_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15368_ (.A(net1),
    .B(net361),
    .CO(_07456_),
    .S(_07457_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15369_ (.A(_07136_),
    .B(_07458_),
    .CO(_07459_),
    .S(_07460_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15370_ (.A(_07136_),
    .B(_07461_),
    .CO(_07462_),
    .S(_07463_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15371_ (.A(_07123_),
    .B(_07464_),
    .CO(_07465_),
    .S(_07466_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15372_ (.A(net2),
    .B(_07467_),
    .CO(_07468_),
    .S(_07469_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15373_ (.A(_07091_),
    .B(_07470_),
    .CO(_07471_),
    .S(_07472_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15374_ (.A(_07082_),
    .B(_07473_),
    .CO(_07474_),
    .S(_07475_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15375_ (.A(_05862_),
    .B(_07476_),
    .CO(_07477_),
    .S(_07478_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15376_ (.A(net1),
    .B(net362),
    .CO(_07479_),
    .S(_07480_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15377_ (.A(_07136_),
    .B(_07481_),
    .CO(_07482_),
    .S(_07483_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15378_ (.A(_07123_),
    .B(_07484_),
    .CO(_07485_),
    .S(_07486_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15379_ (.A(net2),
    .B(_07487_),
    .CO(_07488_),
    .S(_07489_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15380_ (.A(_07091_),
    .B(_07490_),
    .CO(_07491_),
    .S(_07492_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15381_ (.A(_07082_),
    .B(_07493_),
    .CO(_07494_),
    .S(_07495_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15382_ (.A(_05862_),
    .B(_07496_),
    .CO(_07497_),
    .S(_07498_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15383_ (.A(net1),
    .B(net363),
    .CO(_07499_),
    .S(_07500_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15384_ (.A(net1),
    .B(net364),
    .CO(_07501_),
    .S(_07502_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15385_ (.A(_07136_),
    .B(_07503_),
    .CO(_07504_),
    .S(_07505_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15386_ (.A(_07123_),
    .B(_07506_),
    .CO(_07507_),
    .S(_07508_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15387_ (.A(net2),
    .B(_07509_),
    .CO(_07510_),
    .S(_07511_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15388_ (.A(_07091_),
    .B(_07512_),
    .CO(_07513_),
    .S(_07514_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15389_ (.A(_07082_),
    .B(_07515_),
    .CO(_07516_),
    .S(_07517_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15390_ (.A(_05862_),
    .B(_07518_),
    .CO(_07519_),
    .S(_07520_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15391_ (.A(_05862_),
    .B(_07521_),
    .CO(_07522_),
    .S(_07523_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15392_ (.A(net1),
    .B(net365),
    .CO(_07524_),
    .S(_07525_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15393_ (.A(_07177_),
    .B(_07526_),
    .CO(_07527_),
    .S(_07528_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15394_ (.A(_07136_),
    .B(_07529_),
    .CO(_07530_),
    .S(_07531_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15395_ (.A(_07123_),
    .B(_07532_),
    .CO(_07533_),
    .S(_07534_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15396_ (.A(net2),
    .B(_07535_),
    .CO(_07536_),
    .S(_07537_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15397_ (.A(_07091_),
    .B(_07538_),
    .CO(_07539_),
    .S(_07540_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15398_ (.A(_07082_),
    .B(_07541_),
    .CO(_07542_),
    .S(_07543_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15399_ (.A(net1),
    .B(net366),
    .CO(_07544_),
    .S(_07545_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15400_ (.A(_07082_),
    .B(_07546_),
    .CO(_07547_),
    .S(_07548_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15401_ (.A(_05862_),
    .B(_07549_),
    .CO(_07550_),
    .S(_07551_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15402_ (.A(_07177_),
    .B(_07552_),
    .CO(_07553_),
    .S(_07554_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15403_ (.A(_07136_),
    .B(_07555_),
    .CO(_07556_),
    .S(_07557_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15404_ (.A(_07123_),
    .B(_07558_),
    .CO(_07559_),
    .S(_07560_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15405_ (.A(net2),
    .B(_07561_),
    .CO(_07562_),
    .S(_07563_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15406_ (.A(_07091_),
    .B(_07564_),
    .CO(_07565_),
    .S(_07566_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15407_ (.A(_07091_),
    .B(_07567_),
    .CO(_07568_),
    .S(_07569_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15408_ (.A(_07082_),
    .B(_07570_),
    .CO(_07571_),
    .S(_07572_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15409_ (.A(_05862_),
    .B(_07573_),
    .CO(_07574_),
    .S(_07575_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15410_ (.A(net1),
    .B(net367),
    .CO(_07576_),
    .S(_07577_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15411_ (.A(_07177_),
    .B(_07578_),
    .CO(_07579_),
    .S(_07580_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15412_ (.A(_07136_),
    .B(_07581_),
    .CO(_07582_),
    .S(_07583_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15413_ (.A(_07123_),
    .B(_07584_),
    .CO(_07585_),
    .S(_07586_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15414_ (.A(net2),
    .B(_07587_),
    .CO(_07588_),
    .S(_07589_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15415_ (.A(net1),
    .B(net368),
    .CO(_07590_),
    .S(_07591_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15416_ (.A(_07082_),
    .B(_07592_),
    .CO(_07593_),
    .S(_07594_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15417_ (.A(_05862_),
    .B(_07595_),
    .CO(_07596_),
    .S(_07597_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15418_ (.A(net2),
    .B(_07598_),
    .CO(_07599_),
    .S(_07600_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15419_ (.A(_07091_),
    .B(_07601_),
    .CO(_07602_),
    .S(_07603_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15420_ (.A(_07136_),
    .B(_07604_),
    .CO(_07605_),
    .S(_07606_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15421_ (.A(_07123_),
    .B(_07607_),
    .CO(_07608_),
    .S(_07609_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15422_ (.A(_07177_),
    .B(_07610_),
    .CO(_07611_),
    .S(_07612_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15423_ (.A(_05862_),
    .B(_07613_),
    .CO(_07614_),
    .S(_07615_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15424_ (.A(\butterfly_count[2] ),
    .B(net1),
    .CO(_07616_),
    .S(_07617_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15425_ (.A(_07123_),
    .B(_07618_),
    .CO(_07619_),
    .S(_07620_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15426_ (.A(net2),
    .B(_07621_),
    .CO(_07622_),
    .S(_07623_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15427_ (.A(_07091_),
    .B(_07624_),
    .CO(_07625_),
    .S(_07626_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15428_ (.A(_07082_),
    .B(_07627_),
    .CO(_07628_),
    .S(_07629_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15429_ (.A(_07177_),
    .B(_07630_),
    .CO(_07631_),
    .S(_07632_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15430_ (.A(_07136_),
    .B(_07633_),
    .CO(_07634_),
    .S(_07635_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15431_ (.A(_07636_),
    .B(_07637_),
    .CO(_07638_),
    .S(_07639_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15432_ (.A(\butterfly_count[1] ),
    .B(net1),
    .CO(_07640_),
    .S(_07641_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15433_ (.A(_07082_),
    .B(_07642_),
    .CO(_07643_),
    .S(_07644_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15434_ (.A(_05862_),
    .B(_07645_),
    .CO(_07646_),
    .S(_07647_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15435_ (.A(_07136_),
    .B(_07648_),
    .CO(_07649_),
    .S(_07650_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15436_ (.A(_07123_),
    .B(_07651_),
    .CO(_07652_),
    .S(_07653_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15437_ (.A(net2),
    .B(_07654_),
    .CO(_07655_),
    .S(_07656_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15438_ (.A(_07091_),
    .B(_07657_),
    .CO(_07658_),
    .S(_07659_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15439_ (.A(_07660_),
    .B(_07661_),
    .CO(_07662_),
    .S(_07663_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15440_ (.A(_07664_),
    .B(_07665_),
    .CO(_07666_),
    .S(_07667_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15441_ (.A(_07669_),
    .B(_07668_),
    .CO(_07670_),
    .S(_07671_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15442_ (.A(_07672_),
    .B(_07673_),
    .CO(_07674_),
    .S(_07675_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15443_ (.A(_07676_),
    .B(_07677_),
    .CO(_07678_),
    .S(_07679_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15444_ (.A(_07680_),
    .B(_07681_),
    .CO(_07682_),
    .S(_07683_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15445_ (.A(_05862_),
    .B(_05863_),
    .CO(_07684_),
    .S(_07685_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15446_ (.A(_07686_),
    .B(_07637_),
    .CO(_07687_),
    .S(_07688_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15447_ (.A(\butterfly_count[0] ),
    .B(net1),
    .CO(_07689_),
    .S(_07690_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15448_ (.A(_05852_),
    .B(_07691_),
    .CO(_07692_),
    .S(_07693_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15449_ (.A(\temp_real[0] ),
    .B(_07691_),
    .CO(_07694_),
    .S(_07695_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15450_ (.A(_05852_),
    .B(_07696_),
    .CO(_07697_),
    .S(_07698_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15451_ (.A(\temp_real[0] ),
    .B(_07696_),
    .CO(_07699_),
    .S(_07700_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15452_ (.A(\temp_real[0] ),
    .B(_07702_),
    .CO(_07701_),
    .S(_07703_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15453_ (.A(\temp_real[0] ),
    .B(_07704_),
    .CO(_05861_),
    .S(_07705_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15454_ (.A(_07706_),
    .B(_07707_),
    .CO(_07708_),
    .S(_07709_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15455_ (.A(_05852_),
    .B(_07710_),
    .CO(_07711_),
    .S(_07712_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15456_ (.A(\temp_real[0] ),
    .B(_07710_),
    .CO(_07713_),
    .S(_07714_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15457_ (.A(_05852_),
    .B(_07715_),
    .CO(_07716_),
    .S(_07717_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15458_ (.A(\temp_real[0] ),
    .B(_07715_),
    .CO(_07718_),
    .S(_07719_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15459_ (.A(_05852_),
    .B(_07720_),
    .CO(_07721_),
    .S(_07722_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15460_ (.A(\temp_real[0] ),
    .B(_07720_),
    .CO(_07723_),
    .S(_07724_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15461_ (.A(_05852_),
    .B(_07725_),
    .CO(_07726_),
    .S(_07727_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15462_ (.A(\temp_real[0] ),
    .B(_07725_),
    .CO(_07728_),
    .S(_07729_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15463_ (.A(_05852_),
    .B(_07730_),
    .CO(_07731_),
    .S(_07732_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15464_ (.A(\temp_real[0] ),
    .B(_07730_),
    .CO(_07733_),
    .S(_07734_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15465_ (.A(_05852_),
    .B(_07735_),
    .CO(_07736_),
    .S(_07737_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15466_ (.A(\temp_real[0] ),
    .B(_07735_),
    .CO(_07738_),
    .S(_07739_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15467_ (.A(_05852_),
    .B(_07740_),
    .CO(_07741_),
    .S(_07742_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15468_ (.A(\temp_real[0] ),
    .B(_07740_),
    .CO(_07743_),
    .S(_07744_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15469_ (.A(_05852_),
    .B(_07745_),
    .CO(_07746_),
    .S(_07747_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15470_ (.A(\temp_real[0] ),
    .B(_07745_),
    .CO(_07748_),
    .S(_07749_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15471_ (.A(_05852_),
    .B(_07750_),
    .CO(_07751_),
    .S(_07752_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15472_ (.A(\temp_real[0] ),
    .B(_07750_),
    .CO(_07753_),
    .S(_07754_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15473_ (.A(_05852_),
    .B(_07755_),
    .CO(_07756_),
    .S(_07757_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15474_ (.A(\temp_real[0] ),
    .B(_07755_),
    .CO(_07758_),
    .S(_07759_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15475_ (.A(_05852_),
    .B(_07760_),
    .CO(_07761_),
    .S(_07762_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15476_ (.A(\temp_real[0] ),
    .B(_07760_),
    .CO(_07763_),
    .S(_07764_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15477_ (.A(_05852_),
    .B(_05857_),
    .CO(_07765_),
    .S(_07766_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15478_ (.A(\temp_real[0] ),
    .B(_05857_),
    .CO(_07767_),
    .S(_07768_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15479_ (.A(_07686_),
    .B(_07636_),
    .CO(_07769_),
    .S(_07770_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15480_ (.A(\butterfly_count[0] ),
    .B(\butterfly_count[1] ),
    .CO(_07771_),
    .S(_07772_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15481_ (.A(_07773_),
    .B(_07774_),
    .CO(_07775_),
    .S(_07776_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15482_ (.A(_07773_),
    .B(_07774_),
    .CO(_07777_),
    .S(_07778_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15483_ (.A(_07773_),
    .B(\stage[1] ),
    .CO(_07779_),
    .S(_07780_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15484_ (.A(\stage[0] ),
    .B(_07774_),
    .CO(_07781_),
    .S(_07782_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15485_ (.A(\stage[0] ),
    .B(_07774_),
    .CO(_07783_),
    .S(_07784_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15486_ (.A(\stage[0] ),
    .B(\stage[1] ),
    .CO(_07785_),
    .S(_07786_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15487_ (.A(_07787_),
    .B(_07788_),
    .CO(_07789_),
    .S(_07790_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15488_ (.A(_07787_),
    .B(_07785_),
    .CO(_07791_),
    .S(_07792_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15489_ (.A(_07787_),
    .B(_07785_),
    .CO(_07676_),
    .S(_07793_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15490_ (.A(\stage[2] ),
    .B(_07785_),
    .CO(_07794_),
    .S(_07795_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15491_ (.A(\stage[2] ),
    .B(_07785_),
    .CO(_07660_),
    .S(_07796_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15492_ (.A(_07797_),
    .B(_07798_),
    .CO(_07799_),
    .S(_07800_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15493_ (.A(\sample_count[0] ),
    .B(\sample_count[1] ),
    .CO(_07801_),
    .S(_07802_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15494_ (.A(\sample_count[2] ),
    .B(_07801_),
    .CO(_07803_),
    .S(_07804_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15495_ (.A(_05867_),
    .B(_07805_),
    .CO(_07806_),
    .S(_07807_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15496_ (.A(\temp_imag[0] ),
    .B(_07805_),
    .CO(_07808_),
    .S(_07809_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15497_ (.A(_05867_),
    .B(_07810_),
    .CO(_07811_),
    .S(_07812_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15498_ (.A(\temp_imag[0] ),
    .B(_07810_),
    .CO(_07813_),
    .S(_07814_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _15499_ (.A(\temp_imag[0] ),
    .B(_07816_),
    .CO(_07815_),
    .S(_07817_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15500_ (.A(\temp_imag[0] ),
    .B(_07818_),
    .CO(_05876_),
    .S(_07819_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15501_ (.A(_07820_),
    .B(_07821_),
    .CO(_07822_),
    .S(_07823_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15502_ (.A(_05867_),
    .B(_07824_),
    .CO(_07825_),
    .S(_07826_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15503_ (.A(\temp_imag[0] ),
    .B(_07824_),
    .CO(_07827_),
    .S(_07828_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15504_ (.A(_05867_),
    .B(_07829_),
    .CO(_07830_),
    .S(_07831_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15505_ (.A(\temp_imag[0] ),
    .B(_07829_),
    .CO(_07832_),
    .S(_07833_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15506_ (.A(_05867_),
    .B(_07834_),
    .CO(_07835_),
    .S(_07836_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15507_ (.A(\temp_imag[0] ),
    .B(_07834_),
    .CO(_07837_),
    .S(_07838_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15508_ (.A(_05867_),
    .B(_07839_),
    .CO(_07840_),
    .S(_07841_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15509_ (.A(\temp_imag[0] ),
    .B(_07839_),
    .CO(_07842_),
    .S(_07843_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15510_ (.A(_05867_),
    .B(_07844_),
    .CO(_07845_),
    .S(_07846_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15511_ (.A(\temp_imag[0] ),
    .B(_07844_),
    .CO(_07847_),
    .S(_07848_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15512_ (.A(_05867_),
    .B(_07849_),
    .CO(_07850_),
    .S(_07851_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15513_ (.A(\temp_imag[0] ),
    .B(_07849_),
    .CO(_07852_),
    .S(_07853_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15514_ (.A(_05867_),
    .B(_07854_),
    .CO(_07855_),
    .S(_07856_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15515_ (.A(\temp_imag[0] ),
    .B(_07854_),
    .CO(_07857_),
    .S(_07858_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15516_ (.A(_05867_),
    .B(_07859_),
    .CO(_07860_),
    .S(_07861_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15517_ (.A(\temp_imag[0] ),
    .B(_07859_),
    .CO(_07862_),
    .S(_07863_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15518_ (.A(_05867_),
    .B(_07864_),
    .CO(_07865_),
    .S(_07866_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15519_ (.A(\temp_imag[0] ),
    .B(_07864_),
    .CO(_07867_),
    .S(_07868_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15520_ (.A(_05867_),
    .B(_07869_),
    .CO(_07870_),
    .S(_07871_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15521_ (.A(\temp_imag[0] ),
    .B(_07869_),
    .CO(_07872_),
    .S(_07873_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15522_ (.A(_05867_),
    .B(_07874_),
    .CO(_07875_),
    .S(_07876_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15523_ (.A(\temp_imag[0] ),
    .B(_07874_),
    .CO(_07877_),
    .S(_07878_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15524_ (.A(_05867_),
    .B(_05872_),
    .CO(_07879_),
    .S(_07880_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15525_ (.A(\temp_imag[0] ),
    .B(_05872_),
    .CO(_07881_),
    .S(_07882_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15526_ (.A(\butterfly_in_group[0] ),
    .B(_07883_),
    .CO(_07884_),
    .S(_00013_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15527_ (.A(\butterfly_in_group[1] ),
    .B(_07885_),
    .CO(_07886_),
    .S(_07887_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15528_ (.A(_07887_),
    .B(_07888_),
    .CO(_07889_),
    .S(_07890_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15529_ (.A(_07890_),
    .B(_07884_),
    .CO(_07891_),
    .S(_00014_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15530_ (.A(_07637_),
    .B(_00013_),
    .CO(_05878_),
    .S(_00015_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15531_ (.A(_05882_),
    .B(_05883_),
    .CO(_07892_),
    .S(_07893_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15532_ (.A(_06093_),
    .B(_06145_),
    .CO(_07894_),
    .S(_07895_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15533_ (.A(_06094_),
    .B(_06205_),
    .CO(_07896_),
    .S(_05913_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15534_ (.A(_05915_),
    .B(_07898_),
    .CO(_07899_),
    .S(_07900_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15535_ (.A(_05921_),
    .B(_07901_),
    .CO(_07902_),
    .S(_07903_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15536_ (.A(_06145_),
    .B(_06471_),
    .CO(_05914_),
    .S(_05955_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15537_ (.A(_05957_),
    .B(_06341_),
    .CO(_05982_),
    .S(_07905_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15538_ (.A(_07906_),
    .B(_05967_),
    .CO(_07907_),
    .S(_06047_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15539_ (.A(_07908_),
    .B(_07909_),
    .CO(_07910_),
    .S(_07911_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15540_ (.A(_06171_),
    .B(_06172_),
    .CO(_07912_),
    .S(_07913_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15541_ (.A(_07914_),
    .B(_07913_),
    .CO(_07915_),
    .S(_07916_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15542_ (.A(_07908_),
    .B(_05882_),
    .CO(_06022_),
    .S(_07917_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15543_ (.A(_06205_),
    .B(_07898_),
    .CO(_05956_),
    .S(_07919_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15544_ (.A(_05968_),
    .B(_07920_),
    .CO(_06048_),
    .S(_06098_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15545_ (.A(_06049_),
    .B(_06101_),
    .CO(_06076_),
    .S(_06084_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15546_ (.A(_07921_),
    .B(_06352_),
    .CO(_07918_),
    .S(_07922_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15547_ (.A(_07922_),
    .B(_07923_),
    .CO(_07924_),
    .S(_06112_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15548_ (.A(_07925_),
    .B(_06255_),
    .CO(_07926_),
    .S(_07927_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15549_ (.A(_06145_),
    .B(_06205_),
    .CO(_07928_),
    .S(_07929_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15550_ (.A(_06471_),
    .B(_06341_),
    .CO(_07930_),
    .S(_07931_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15551_ (.A(_07928_),
    .B(_07931_),
    .CO(_06137_),
    .S(_07932_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15552_ (.A(_07933_),
    .B(_07934_),
    .CO(_06099_),
    .S(_06148_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15553_ (.A(_06102_),
    .B(_06151_),
    .CO(_06122_),
    .S(_06133_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15554_ (.A(_07913_),
    .B(_06004_),
    .CO(_06115_),
    .S(_06165_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15555_ (.A(_07935_),
    .B(_07936_),
    .CO(_07937_),
    .S(_06163_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15556_ (.A(_06120_),
    .B(_07924_),
    .CO(_07938_),
    .S(_06124_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15557_ (.A(_06205_),
    .B(_06471_),
    .CO(_07939_),
    .S(_07940_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15558_ (.A(_07898_),
    .B(_07939_),
    .CO(_06197_),
    .S(_07941_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15559_ (.A(_07942_),
    .B(_06155_),
    .CO(_06149_),
    .S(_06208_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15560_ (.A(_06152_),
    .B(_06211_),
    .CO(_06175_),
    .S(_06193_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15561_ (.A(_06352_),
    .B(_06173_),
    .CO(_06166_),
    .S(_07943_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15562_ (.A(_05883_),
    .B(_05907_),
    .CO(_07944_),
    .S(_07945_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15563_ (.A(_07946_),
    .B(_07947_),
    .CO(_07948_),
    .S(_07949_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15564_ (.A(_07951_),
    .B(_07937_),
    .CO(_06181_),
    .S(_06185_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15565_ (.A(_06341_),
    .B(_07952_),
    .CO(_06247_),
    .S(_07953_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15566_ (.A(_06156_),
    .B(_07954_),
    .CO(_06209_),
    .S(_06258_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15567_ (.A(_06212_),
    .B(_06261_),
    .CO(_06226_),
    .S(_06243_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15568_ (.A(_06219_),
    .B(_07943_),
    .CO(_07950_),
    .S(_07955_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15569_ (.A(_06002_),
    .B(_06352_),
    .CO(_07956_),
    .S(_06268_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15570_ (.A(_05907_),
    .B(_05908_),
    .CO(_07957_),
    .S(_07958_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15571_ (.A(_05895_),
    .B(_05888_),
    .CO(_07959_),
    .S(_07960_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15572_ (.A(_07962_),
    .B(_07948_),
    .CO(_06231_),
    .S(_06235_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15573_ (.A(_06183_),
    .B(_06232_),
    .CO(_07963_),
    .S(_07964_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15574_ (.A(_07965_),
    .B(_07966_),
    .CO(_06259_),
    .S(_06305_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15575_ (.A(_06262_),
    .B(_06308_),
    .CO(_06280_),
    .S(_06294_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15576_ (.A(_05908_),
    .B(_05950_),
    .CO(_07967_),
    .S(_07968_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15577_ (.A(_07897_),
    .B(_05905_),
    .CO(_07969_),
    .S(_07970_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15578_ (.A(_06269_),
    .B(_07956_),
    .CO(_07961_),
    .S(_07971_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15579_ (.A(_06278_),
    .B(_07959_),
    .CO(_06282_),
    .S(_06286_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15580_ (.A(_06233_),
    .B(_06283_),
    .CO(_07972_),
    .S(_07973_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15581_ (.A(_07974_),
    .B(_07975_),
    .CO(_06293_),
    .S(_06333_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15582_ (.A(_07976_),
    .B(_07977_),
    .CO(_06306_),
    .S(_06343_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15583_ (.A(_06309_),
    .B(_06346_),
    .CO(_07978_),
    .S(_06335_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15584_ (.A(_07970_),
    .B(_07971_),
    .CO(_06277_),
    .S(_06319_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15585_ (.A(_05950_),
    .B(_06093_),
    .CO(_05912_),
    .S(_07979_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15586_ (.A(_07904_),
    .B(_05948_),
    .CO(_07980_),
    .S(_07981_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15587_ (.A(_06321_),
    .B(_07969_),
    .CO(_06324_),
    .S(_06328_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15588_ (.A(_06284_),
    .B(_06325_),
    .CO(_07982_),
    .S(_07983_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15589_ (.A(_07984_),
    .B(_07985_),
    .CO(_06334_),
    .S(_06370_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15590_ (.A(_07986_),
    .B(_07987_),
    .CO(_07985_),
    .S(_07988_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15591_ (.A(_07898_),
    .B(_06404_),
    .CO(_06342_),
    .S(_06426_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15592_ (.A(_07989_),
    .B(_06350_),
    .CO(_06344_),
    .S(_06379_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15593_ (.A(_06353_),
    .B(_07990_),
    .CO(_07991_),
    .S(_06376_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15594_ (.A(_06347_),
    .B(_07992_),
    .CO(_07993_),
    .S(_06372_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15595_ (.A(_07981_),
    .B(_06316_),
    .CO(_06320_),
    .S(_06355_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15596_ (.A(_06093_),
    .B(_06094_),
    .CO(_05954_),
    .S(_07994_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15597_ (.A(_06042_),
    .B(_06037_),
    .CO(_07995_),
    .S(_07996_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15598_ (.A(_06357_),
    .B(_07980_),
    .CO(_06360_),
    .S(_06364_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15599_ (.A(_06326_),
    .B(_06361_),
    .CO(_07997_),
    .S(_07998_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15600_ (.A(_07988_),
    .B(_07999_),
    .CO(_06371_),
    .S(_08000_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15601_ (.A(_06351_),
    .B(_08001_),
    .CO(_06380_),
    .S(_06402_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15602_ (.A(_06016_),
    .B(_08002_),
    .CO(_08001_),
    .S(_08003_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15603_ (.A(_06172_),
    .B(_06352_),
    .CO(_07990_),
    .S(_08004_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15604_ (.A(_08004_),
    .B(_08005_),
    .CO(_08006_),
    .S(_06399_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15605_ (.A(_08007_),
    .B(_08008_),
    .CO(_08009_),
    .S(_08010_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15606_ (.A(_07996_),
    .B(_07991_),
    .CO(_06356_),
    .S(_06382_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15607_ (.A(_06145_),
    .B(_06094_),
    .CO(_08011_),
    .S(_08012_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15608_ (.A(_08013_),
    .B(_06091_),
    .CO(_08014_),
    .S(_08015_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15609_ (.A(_06384_),
    .B(_07995_),
    .CO(_06387_),
    .S(_06391_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15610_ (.A(_06362_),
    .B(_06388_),
    .CO(_08016_),
    .S(_08017_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15611_ (.A(_08000_),
    .B(_08010_),
    .CO(_06396_),
    .S(_06420_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15612_ (.A(_08018_),
    .B(_08019_),
    .CO(_07999_),
    .S(_08020_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15613_ (.A(_08003_),
    .B(_06407_),
    .CO(_06403_),
    .S(_06433_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15614_ (.A(_06352_),
    .B(_08021_),
    .CO(_08005_),
    .S(_06430_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15615_ (.A(_08022_),
    .B(_08023_),
    .CO(_08024_),
    .S(_08025_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15616_ (.A(_08015_),
    .B(_08006_),
    .CO(_06383_),
    .S(_08026_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15617_ (.A(_08027_),
    .B(_08026_),
    .CO(_08028_),
    .S(_06416_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15618_ (.A(_08028_),
    .B(_08014_),
    .CO(_06410_),
    .S(_06414_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15619_ (.A(_06389_),
    .B(_06411_),
    .CO(_08029_),
    .S(_08030_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15620_ (.A(_08020_),
    .B(_08025_),
    .CO(_06421_),
    .S(_08031_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15621_ (.A(_06408_),
    .B(_06438_),
    .CO(_06434_),
    .S(_08032_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15622_ (.A(_08033_),
    .B(_08034_),
    .CO(_08035_),
    .S(_08036_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15623_ (.A(_08037_),
    .B(_08038_),
    .CO(_08039_),
    .S(_06449_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15624_ (.A(_06412_),
    .B(_06442_),
    .CO(_08040_),
    .S(_08041_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15625_ (.A(_08042_),
    .B(_08036_),
    .CO(_08043_),
    .S(_06462_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15626_ (.A(_06341_),
    .B(_06435_),
    .CO(_06427_),
    .S(_08044_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15627_ (.A(_08045_),
    .B(_08046_),
    .CO(_08047_),
    .S(_08048_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15628_ (.A(_06439_),
    .B(_08049_),
    .CO(_08050_),
    .S(_08051_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15629_ (.A(_08052_),
    .B(_08053_),
    .CO(_08054_),
    .S(_08055_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15630_ (.A(_08056_),
    .B(_08057_),
    .CO(_08058_),
    .S(_08059_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15631_ (.A(_06205_),
    .B(_06451_),
    .CO(_08060_),
    .S(_08061_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15632_ (.A(_06452_),
    .B(_08061_),
    .CO(_08062_),
    .S(_08063_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15633_ (.A(_08062_),
    .B(_08060_),
    .CO(_06456_),
    .S(_08064_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15634_ (.A(_06443_),
    .B(_06457_),
    .CO(_08065_),
    .S(_08066_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15635_ (.A(_08067_),
    .B(_08068_),
    .CO(_06466_),
    .S(_08069_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15636_ (.A(_08070_),
    .B(_08055_),
    .CO(_08071_),
    .S(_08072_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15637_ (.A(_06471_),
    .B(_07898_),
    .CO(_07952_),
    .S(_06468_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15638_ (.A(_06296_),
    .B(_06253_),
    .CO(_06477_),
    .S(_08073_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15639_ (.A(_08072_),
    .B(_08073_),
    .CO(_06476_),
    .S(_08074_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15640_ (.A(_06458_),
    .B(_06480_),
    .CO(_08075_),
    .S(_08076_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15641_ (.A(_08077_),
    .B(_06470_),
    .CO(_06486_),
    .S(_06491_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15642_ (.A(_07898_),
    .B(_06341_),
    .CO(_06299_),
    .S(_08078_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15643_ (.A(_08079_),
    .B(_08078_),
    .CO(_06493_),
    .S(_08080_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15644_ (.A(_08081_),
    .B(_08078_),
    .CO(_08082_),
    .S(_08083_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15645_ (.A(_06481_),
    .B(_06489_),
    .CO(_08085_),
    .S(_08086_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15646_ (.A(_06467_),
    .B(_08087_),
    .CO(_08084_),
    .S(_08088_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15647_ (.A(_08089_),
    .B(_08090_),
    .CO(_08081_),
    .S(_08091_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15648_ (.A(_06490_),
    .B(_08092_),
    .CO(_08093_),
    .S(_08094_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15649_ (.A(_06495_),
    .B(_08095_),
    .CO(_08092_),
    .S(_08096_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15650_ (.A(_08088_),
    .B(_08097_),
    .CO(_08098_),
    .S(_08099_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15651_ (.A(_06341_),
    .B(_08091_),
    .CO(_08097_),
    .S(_08100_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15652_ (.A(_08101_),
    .B(_08102_),
    .CO(_08103_),
    .S(_08104_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15653_ (.A(_08105_),
    .B(_08104_),
    .CO(_08106_),
    .S(_06528_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15654_ (.A(_08107_),
    .B(_06691_),
    .CO(_08108_),
    .S(_08109_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15655_ (.A(_06504_),
    .B(_06616_),
    .CO(_06529_),
    .S(_06563_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15656_ (.A(_08101_),
    .B(_06501_),
    .CO(_06537_),
    .S(_08110_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15657_ (.A(_08111_),
    .B(_08112_),
    .CO(_08113_),
    .S(_06555_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15658_ (.A(_08114_),
    .B(_08115_),
    .CO(_06556_),
    .S(_06592_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15659_ (.A(_06748_),
    .B(_08116_),
    .CO(_08117_),
    .S(_06588_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15660_ (.A(_08110_),
    .B(_06663_),
    .CO(_06564_),
    .S(_08118_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15661_ (.A(_08119_),
    .B(_08120_),
    .CO(_06583_),
    .S(_08121_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15662_ (.A(_08123_),
    .B(_08124_),
    .CO(_06593_),
    .S(_06651_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15663_ (.A(_06803_),
    .B(_06961_),
    .CO(_08125_),
    .S(_06647_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15664_ (.A(_06956_),
    .B(_08126_),
    .CO(_08127_),
    .S(_08128_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15665_ (.A(_06618_),
    .B(_06913_),
    .CO(_08129_),
    .S(_08130_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15666_ (.A(_08127_),
    .B(_08130_),
    .CO(_08131_),
    .S(_08132_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15667_ (.A(_08116_),
    .B(_06913_),
    .CO(_08134_),
    .S(_08135_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15668_ (.A(_08128_),
    .B(_08134_),
    .CO(_08133_),
    .S(_08136_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15669_ (.A(_08137_),
    .B(_06665_),
    .CO(_08138_),
    .S(_08139_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15670_ (.A(_08141_),
    .B(_06684_),
    .CO(_06642_),
    .S(_08142_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15671_ (.A(_08101_),
    .B(_06601_),
    .CO(_08122_),
    .S(_08143_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15672_ (.A(_08144_),
    .B(_08145_),
    .CO(_06652_),
    .S(_06703_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15673_ (.A(_08146_),
    .B(_08136_),
    .CO(_08140_),
    .S(_08147_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15674_ (.A(_06961_),
    .B(_06956_),
    .CO(_08148_),
    .S(_08149_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15675_ (.A(_08148_),
    .B(_08135_),
    .CO(_08146_),
    .S(_08150_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15676_ (.A(_06666_),
    .B(_06717_),
    .CO(_08151_),
    .S(_08152_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15677_ (.A(_08142_),
    .B(_08143_),
    .CO(_06680_),
    .S(_06736_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15678_ (.A(_06685_),
    .B(_08154_),
    .CO(_06695_),
    .S(_08155_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15679_ (.A(_08156_),
    .B(_08157_),
    .CO(_06704_),
    .S(_06752_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15680_ (.A(_08158_),
    .B(_08150_),
    .CO(_08153_),
    .S(_08159_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15681_ (.A(_06699_),
    .B(_08116_),
    .CO(_08160_),
    .S(_08161_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15682_ (.A(_08160_),
    .B(_08149_),
    .CO(_08158_),
    .S(_08162_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15683_ (.A(_06718_),
    .B(_06765_),
    .CO(_08163_),
    .S(_08164_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15684_ (.A(_08166_),
    .B(_08151_),
    .CO(_08167_),
    .S(_06727_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15685_ (.A(_06602_),
    .B(_08155_),
    .CO(_06737_),
    .S(_06789_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15686_ (.A(_08101_),
    .B(_06496_),
    .CO(_08154_),
    .S(_08168_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15687_ (.A(_06742_),
    .B(_06796_),
    .CO(_06755_),
    .S(_06791_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15688_ (.A(_08169_),
    .B(_08170_),
    .CO(_06753_),
    .S(_06807_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15689_ (.A(_08171_),
    .B(_08162_),
    .CO(_08165_),
    .S(_08172_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15690_ (.A(_06748_),
    .B(_06961_),
    .CO(_08173_),
    .S(_08174_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15691_ (.A(_08173_),
    .B(_08161_),
    .CO(_08171_),
    .S(_08175_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15692_ (.A(_06766_),
    .B(_06821_),
    .CO(_08176_),
    .S(_08177_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15693_ (.A(_08179_),
    .B(_08163_),
    .CO(_06775_),
    .S(_06780_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15694_ (.A(_06618_),
    .B(_08168_),
    .CO(_06790_),
    .S(_08180_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15695_ (.A(_06797_),
    .B(_06853_),
    .CO(_08181_),
    .S(_08182_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15696_ (.A(_08184_),
    .B(_08185_),
    .CO(_06808_),
    .S(_06861_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15697_ (.A(_06822_),
    .B(_08187_),
    .CO(_08188_),
    .S(_08189_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15698_ (.A(_08190_),
    .B(_08175_),
    .CO(_08178_),
    .S(_08191_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15699_ (.A(_06829_),
    .B(_08176_),
    .CO(_06832_),
    .S(_06837_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15700_ (.A(_06777_),
    .B(_06833_),
    .CO(_08192_),
    .S(_08193_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15701_ (.A(_06854_),
    .B(_08194_),
    .CO(_08195_),
    .S(_08196_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15702_ (.A(_06502_),
    .B(_08126_),
    .CO(_08183_),
    .S(_08197_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15703_ (.A(_06809_),
    .B(_06863_),
    .CO(_08186_),
    .S(_08198_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15704_ (.A(_08199_),
    .B(_08200_),
    .CO(_06862_),
    .S(_06904_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15705_ (.A(_08189_),
    .B(_08191_),
    .CO(_06828_),
    .S(_06876_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15706_ (.A(_08202_),
    .B(_06916_),
    .CO(_08203_),
    .S(_08204_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15707_ (.A(_08205_),
    .B(_08174_),
    .CO(_08190_),
    .S(_08206_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15708_ (.A(_06878_),
    .B(_08188_),
    .CO(_06881_),
    .S(_06886_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15709_ (.A(_06834_),
    .B(_06882_),
    .CO(_08207_),
    .S(_08208_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15710_ (.A(_08196_),
    .B(_08197_),
    .CO(_06893_),
    .S(_06939_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15711_ (.A(_06496_),
    .B(_06502_),
    .CO(_06900_),
    .S(_08209_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15712_ (.A(_08210_),
    .B(_08211_),
    .CO(_08212_),
    .S(_08213_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15713_ (.A(_06864_),
    .B(_06906_),
    .CO(_08201_),
    .S(_08214_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15714_ (.A(_08215_),
    .B(_08216_),
    .CO(_06905_),
    .S(_06947_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15715_ (.A(_08204_),
    .B(_08206_),
    .CO(_06877_),
    .S(_06922_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15716_ (.A(_06917_),
    .B(_06959_),
    .CO(_08218_),
    .S(_08219_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15717_ (.A(_06699_),
    .B(_06803_),
    .CO(_08205_),
    .S(_08220_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15718_ (.A(_06924_),
    .B(_08203_),
    .CO(_06927_),
    .S(_06932_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15719_ (.A(_06883_),
    .B(_06928_),
    .CO(_08221_),
    .S(_08222_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15720_ (.A(_06913_),
    .B(_08213_),
    .CO(_06940_),
    .S(_06981_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15721_ (.A(_08223_),
    .B(_08209_),
    .CO(_08211_),
    .S(_08224_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15722_ (.A(_08224_),
    .B(_08225_),
    .CO(_08226_),
    .S(_08227_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15723_ (.A(_06907_),
    .B(_06949_),
    .CO(_08217_),
    .S(_08228_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15724_ (.A(_08229_),
    .B(_08230_),
    .CO(_06948_),
    .S(_06987_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15725_ (.A(_08219_),
    .B(_08220_),
    .CO(_06923_),
    .S(_06964_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15726_ (.A(_06748_),
    .B(_06803_),
    .CO(_07036_),
    .S(_07074_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15727_ (.A(_06960_),
    .B(_08232_),
    .CO(_08233_),
    .S(_08234_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15728_ (.A(_06966_),
    .B(_08218_),
    .CO(_06969_),
    .S(_06974_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15729_ (.A(_06929_),
    .B(_06970_),
    .CO(_08235_),
    .S(_08236_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15730_ (.A(_06956_),
    .B(_08227_),
    .CO(_06982_),
    .S(_07013_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15731_ (.A(_06502_),
    .B(_08237_),
    .CO(_08225_),
    .S(_08238_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15732_ (.A(_06950_),
    .B(_06989_),
    .CO(_08231_),
    .S(_08239_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15733_ (.A(_08240_),
    .B(_08241_),
    .CO(_06988_),
    .S(_08242_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15734_ (.A(_08239_),
    .B(_08243_),
    .CO(_08244_),
    .S(_07015_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15735_ (.A(_06748_),
    .B(_08234_),
    .CO(_06965_),
    .S(_08245_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15736_ (.A(_06699_),
    .B(_07074_),
    .CO(_08246_),
    .S(_08247_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15737_ (.A(_07036_),
    .B(_06996_),
    .CO(_07058_),
    .S(_07063_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15738_ (.A(_08248_),
    .B(_07037_),
    .CO(_08249_),
    .S(_08250_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15739_ (.A(_08252_),
    .B(_08233_),
    .CO(_07003_),
    .S(_07008_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15740_ (.A(_06971_),
    .B(_07004_),
    .CO(_08253_),
    .S(_08254_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15741_ (.A(_08116_),
    .B(_08238_),
    .CO(_07014_),
    .S(_07032_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15742_ (.A(_06990_),
    .B(_08255_),
    .CO(_08243_),
    .S(_08256_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15743_ (.A(_08258_),
    .B(_08259_),
    .CO(_08257_),
    .S(_08260_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15744_ (.A(_08256_),
    .B(_08261_),
    .CO(_08262_),
    .S(_07034_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15745_ (.A(_06803_),
    .B(_08250_),
    .CO(_08251_),
    .S(_08263_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15746_ (.A(_08262_),
    .B(_08263_),
    .CO(_08264_),
    .S(_07030_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15747_ (.A(_08264_),
    .B(_08249_),
    .CO(_07023_),
    .S(_07027_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15748_ (.A(_07005_),
    .B(_07024_),
    .CO(_08265_),
    .S(_08266_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15749_ (.A(_06961_),
    .B(_07017_),
    .CO(_07033_),
    .S(_07054_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15750_ (.A(_08267_),
    .B(_08268_),
    .CO(_08261_),
    .S(_08269_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15751_ (.A(_08270_),
    .B(_08260_),
    .CO(_08268_),
    .S(_08271_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15752_ (.A(_08272_),
    .B(_08273_),
    .CO(_08270_),
    .S(_08274_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _15753_ (.A(_08269_),
    .B(_08275_),
    .CO(_08276_),
    .S(_07056_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15754_ (.A(_08246_),
    .B(_07038_),
    .CO(_08277_),
    .S(_08278_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15755_ (.A(_08276_),
    .B(_08278_),
    .CO(_08279_),
    .S(_08280_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15756_ (.A(_08279_),
    .B(_08277_),
    .CO(_07045_),
    .S(_08281_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15757_ (.A(_07025_),
    .B(_07046_),
    .CO(_08282_),
    .S(_08283_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15758_ (.A(_06699_),
    .B(_08209_),
    .CO(_07055_),
    .S(_08284_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15759_ (.A(_08271_),
    .B(_08285_),
    .CO(_08275_),
    .S(_08286_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15760_ (.A(_07047_),
    .B(_08288_),
    .CO(_08289_),
    .S(_08290_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15761_ (.A(_07050_),
    .B(_07060_),
    .CO(_08288_),
    .S(_08291_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15762_ (.A(_08292_),
    .B(_08274_),
    .CO(_08285_),
    .S(_08293_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15763_ (.A(_06502_),
    .B(_06748_),
    .CO(_08287_),
    .S(_08294_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15764_ (.A(_08291_),
    .B(_08295_),
    .CO(_08296_),
    .S(_08297_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15765_ (.A(_07061_),
    .B(_08298_),
    .CO(_08295_),
    .S(_08299_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15766_ (.A(_07064_),
    .B(_08300_),
    .CO(_08298_),
    .S(_08301_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15767_ (.A(_08293_),
    .B(_08294_),
    .CO(_07075_),
    .S(_08302_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15768_ (.A(_08303_),
    .B(_08304_),
    .CO(_08292_),
    .S(_08305_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _15769_ (.A(_08302_),
    .B(_08306_),
    .CO(_08307_),
    .S(_08308_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 _15770_ (.D(_00002_),
    .CLK(clknet_leaf_0_clk),
    .Q(_00011_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 _15771_ (.D(_00001_),
    .CLK(clknet_leaf_0_clk),
    .Q(_00010_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _15772_ (.D(_00000_),
    .CLK(clknet_leaf_21_clk),
    .Q(_00008_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 _15773_ (.D(_00018_),
    .CLK(clknet_leaf_0_clk),
    .Q(_00009_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _15774_ (.D(_00019_),
    .CLK(clknet_leaf_0_clk),
    .Q(_00012_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _15775_ (.D(_00020_),
    .CLK(clknet_leaf_0_clk),
    .Q(_00016_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _15776_ (.D(_00021_),
    .CLK(clknet_leaf_0_clk),
    .Q(_00017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__tieh _15237__322 (.Z(net369));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_rev_idx[0]$_DFFE_PN0P_  (.D(_00022_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\bit_rev_idx[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_rev_idx[1]$_DFFE_PN0P_  (.D(_00023_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\bit_rev_idx[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_rev_idx[2]$_DFFE_PN0P_  (.D(_00024_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\bit_rev_idx[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \busy$_DFFE_PN0P_  (.D(_00025_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(net83));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \butterfly_count[0]$_DFFE_PN0P_  (.D(_00026_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\butterfly_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \butterfly_count[1]$_DFFE_PN0P_  (.D(_00027_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\butterfly_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \butterfly_count[2]$_DFFE_PN0P_  (.D(_00028_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\butterfly_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \butterfly_in_group[0]$_DFFE_PP_  (.D(_00029_),
    .CLK(clknet_leaf_20_clk),
    .Q(\butterfly_in_group[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \butterfly_in_group[1]$_DFFE_PP_  (.D(_00030_),
    .CLK(clknet_leaf_20_clk),
    .Q(\butterfly_in_group[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \butterfly_in_group[2]$_DFFE_PP_  (.D(_00031_),
    .CLK(clknet_leaf_20_clk),
    .Q(\butterfly_in_group[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[0]$_DFFE_PN0P_  (.D(_00032_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(net84));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[100]$_DFFE_PN0P_  (.D(_00033_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net85));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[101]$_DFFE_PN0P_  (.D(_00034_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net86));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[102]$_DFFE_PN0P_  (.D(_00035_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net87));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[103]$_DFFE_PN0P_  (.D(_00036_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net88));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[104]$_DFFE_PN0P_  (.D(_00037_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net89));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[105]$_DFFE_PN0P_  (.D(_00038_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net90));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[106]$_DFFE_PN0P_  (.D(_00039_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net91));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[107]$_DFFE_PN0P_  (.D(_00040_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(net92));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[108]$_DFFE_PN0P_  (.D(_00041_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net93));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[109]$_DFFE_PN0P_  (.D(_00042_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net94));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[10]$_DFFE_PN0P_  (.D(_00043_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net95));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[110]$_DFFE_PN0P_  (.D(_00044_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net96));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[111]$_DFFE_PN0P_  (.D(_00045_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net97));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[112]$_DFFE_PN0P_  (.D(_00046_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net98));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[113]$_DFFE_PN0P_  (.D(_00047_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net99));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[114]$_DFFE_PN0P_  (.D(_00048_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[115]$_DFFE_PN0P_  (.D(_00049_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[116]$_DFFE_PN0P_  (.D(_00050_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[117]$_DFFE_PN0P_  (.D(_00051_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[118]$_DFFE_PN0P_  (.D(_00052_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[119]$_DFFE_PN0P_  (.D(_00053_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[11]$_DFFE_PN0P_  (.D(_00054_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[120]$_DFFE_PN0P_  (.D(_00055_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[121]$_DFFE_PN0P_  (.D(_00056_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[122]$_DFFE_PN0P_  (.D(_00057_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[123]$_DFFE_PN0P_  (.D(_00058_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[124]$_DFFE_PN0P_  (.D(_00059_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[125]$_DFFE_PN0P_  (.D(_00060_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[126]$_DFFE_PN0P_  (.D(_00061_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[127]$_DFFE_PN0P_  (.D(_00062_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[12]$_DFFE_PN0P_  (.D(_00063_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[13]$_DFFE_PN0P_  (.D(_00064_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[14]$_DFFE_PN0P_  (.D(_00065_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[15]$_DFFE_PN0P_  (.D(_00066_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[16]$_DFFE_PN0P_  (.D(_00067_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[17]$_DFFE_PN0P_  (.D(_00068_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[18]$_DFFE_PN0P_  (.D(_00069_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[19]$_DFFE_PN0P_  (.D(_00070_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[1]$_DFFE_PN0P_  (.D(_00071_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[20]$_DFFE_PN0P_  (.D(_00072_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[21]$_DFFE_PN0P_  (.D(_00073_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[22]$_DFFE_PN0P_  (.D(_00074_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[23]$_DFFE_PN0P_  (.D(_00075_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(net127));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[24]$_DFFE_PN0P_  (.D(_00076_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(net128));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[25]$_DFFE_PN0P_  (.D(_00077_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(net129));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[26]$_DFFE_PN0P_  (.D(_00078_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net130));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[27]$_DFFE_PN0P_  (.D(_00079_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net131));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[28]$_DFFE_PN0P_  (.D(_00080_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net132));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[29]$_DFFE_PN0P_  (.D(_00081_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net133));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[2]$_DFFE_PN0P_  (.D(_00082_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net134));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[30]$_DFFE_PN0P_  (.D(_00083_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net135));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[31]$_DFFE_PN0P_  (.D(_00084_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net136));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[32]$_DFFE_PN0P_  (.D(_00085_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net137));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[33]$_DFFE_PN0P_  (.D(_00086_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net138));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[34]$_DFFE_PN0P_  (.D(_00087_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net139));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[35]$_DFFE_PN0P_  (.D(_00088_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net140));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[36]$_DFFE_PN0P_  (.D(_00089_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net141));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[37]$_DFFE_PN0P_  (.D(_00090_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net142));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[38]$_DFFE_PN0P_  (.D(_00091_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net143));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[39]$_DFFE_PN0P_  (.D(_00092_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net144));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[3]$_DFFE_PN0P_  (.D(_00093_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net145));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[40]$_DFFE_PN0P_  (.D(_00094_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net146));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[41]$_DFFE_PN0P_  (.D(_00095_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net147));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[42]$_DFFE_PN0P_  (.D(_00096_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net148));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[43]$_DFFE_PN0P_  (.D(_00097_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net149));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[44]$_DFFE_PN0P_  (.D(_00098_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net150));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[45]$_DFFE_PN0P_  (.D(_00099_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net151));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[46]$_DFFE_PN0P_  (.D(_00100_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net152));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[47]$_DFFE_PN0P_  (.D(_00101_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net153));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[48]$_DFFE_PN0P_  (.D(_00102_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net154));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[49]$_DFFE_PN0P_  (.D(_00103_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net155));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[4]$_DFFE_PN0P_  (.D(_00104_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net156));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[50]$_DFFE_PN0P_  (.D(_00105_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net157));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[51]$_DFFE_PN0P_  (.D(_00106_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net158));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[52]$_DFFE_PN0P_  (.D(_00107_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net159));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[53]$_DFFE_PN0P_  (.D(_00108_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net160));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[54]$_DFFE_PN0P_  (.D(_00109_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net161));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[55]$_DFFE_PN0P_  (.D(_00110_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net162));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[56]$_DFFE_PN0P_  (.D(_00111_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net163));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[57]$_DFFE_PN0P_  (.D(_00112_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net164));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[58]$_DFFE_PN0P_  (.D(_00113_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net165));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[59]$_DFFE_PN0P_  (.D(_00114_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net166));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[5]$_DFFE_PN0P_  (.D(_00115_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net167));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[60]$_DFFE_PN0P_  (.D(_00116_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(net168));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[61]$_DFFE_PN0P_  (.D(_00117_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(net169));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[62]$_DFFE_PN0P_  (.D(_00118_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net170));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[63]$_DFFE_PN0P_  (.D(_00119_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net171));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[64]$_DFFE_PN0P_  (.D(_00120_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(net172));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[65]$_DFFE_PN0P_  (.D(_00121_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net173));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[66]$_DFFE_PN0P_  (.D(_00122_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net174));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[67]$_DFFE_PN0P_  (.D(_00123_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net175));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[68]$_DFFE_PN0P_  (.D(_00124_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net176));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[69]$_DFFE_PN0P_  (.D(_00125_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(net177));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[6]$_DFFE_PN0P_  (.D(_00126_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net178));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[70]$_DFFE_PN0P_  (.D(_00127_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(net179));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[71]$_DFFE_PN0P_  (.D(_00128_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(net180));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[72]$_DFFE_PN0P_  (.D(_00129_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net181));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[73]$_DFFE_PN0P_  (.D(_00130_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net182));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[74]$_DFFE_PN0P_  (.D(_00131_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net183));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[75]$_DFFE_PN0P_  (.D(_00132_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net184));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[76]$_DFFE_PN0P_  (.D(_00133_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net185));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[77]$_DFFE_PN0P_  (.D(_00134_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net186));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[78]$_DFFE_PN0P_  (.D(_00135_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net187));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[79]$_DFFE_PN0P_  (.D(_00136_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net188));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[7]$_DFFE_PN0P_  (.D(_00137_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net189));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[80]$_DFFE_PN0P_  (.D(_00138_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net190));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[81]$_DFFE_PN0P_  (.D(_00139_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net191));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[82]$_DFFE_PN0P_  (.D(_00140_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net192));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[83]$_DFFE_PN0P_  (.D(_00141_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net193));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[84]$_DFFE_PN0P_  (.D(_00142_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(net194));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[85]$_DFFE_PN0P_  (.D(_00143_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net195));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[86]$_DFFE_PN0P_  (.D(_00144_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net196));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[87]$_DFFE_PN0P_  (.D(_00145_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net197));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[88]$_DFFE_PN0P_  (.D(_00146_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net198));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[89]$_DFFE_PN0P_  (.D(_00147_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net199));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[8]$_DFFE_PN0P_  (.D(_00148_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net200));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[90]$_DFFE_PN0P_  (.D(_00149_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(net201));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[91]$_DFFE_PN0P_  (.D(_00150_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(net202));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[92]$_DFFE_PN0P_  (.D(_00151_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(net203));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[93]$_DFFE_PN0P_  (.D(_00152_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(net204));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[94]$_DFFE_PN0P_  (.D(_00153_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net205));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[95]$_DFFE_PN0P_  (.D(_00154_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(net206));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[96]$_DFFE_PN0P_  (.D(_00155_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(net207));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[97]$_DFFE_PN0P_  (.D(_00156_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net208));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[98]$_DFFE_PN0P_  (.D(_00157_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net209));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[99]$_DFFE_PN0P_  (.D(_00158_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(net210));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_imag[9]$_DFFE_PN0P_  (.D(_00159_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(net211));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[0]$_DFFE_PN0P_  (.D(_00160_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(net212));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[100]$_DFFE_PN0P_  (.D(_00161_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net213));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[101]$_DFFE_PN0P_  (.D(_00162_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net214));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[102]$_DFFE_PN0P_  (.D(_00163_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net215));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[103]$_DFFE_PN0P_  (.D(_00164_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net216));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[104]$_DFFE_PN0P_  (.D(_00165_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net217));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[105]$_DFFE_PN0P_  (.D(_00166_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net218));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[106]$_DFFE_PN0P_  (.D(_00167_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net219));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[107]$_DFFE_PN0P_  (.D(_00168_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(net220));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[108]$_DFFE_PN0P_  (.D(_00169_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net221));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[109]$_DFFE_PN0P_  (.D(_00170_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net222));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[10]$_DFFE_PN0P_  (.D(_00171_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net223));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[110]$_DFFE_PN0P_  (.D(_00172_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net224));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[111]$_DFFE_PN0P_  (.D(_00173_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net225));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[112]$_DFFE_PN0P_  (.D(_00174_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net226));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[113]$_DFFE_PN0P_  (.D(_00175_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net227));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[114]$_DFFE_PN0P_  (.D(_00176_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net228));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[115]$_DFFE_PN0P_  (.D(_00177_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net229));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[116]$_DFFE_PN0P_  (.D(_00178_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net230));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[117]$_DFFE_PN0P_  (.D(_00179_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net231));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[118]$_DFFE_PN0P_  (.D(_00180_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net232));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[119]$_DFFE_PN0P_  (.D(_00181_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net233));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[11]$_DFFE_PN0P_  (.D(_00182_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net234));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[120]$_DFFE_PN0P_  (.D(_00183_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net235));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[121]$_DFFE_PN0P_  (.D(_00184_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net236));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[122]$_DFFE_PN0P_  (.D(_00185_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net237));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[123]$_DFFE_PN0P_  (.D(_00186_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(net238));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[124]$_DFFE_PN0P_  (.D(_00187_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net239));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[125]$_DFFE_PN0P_  (.D(_00188_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net240));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[126]$_DFFE_PN0P_  (.D(_00189_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net241));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[127]$_DFFE_PN0P_  (.D(_00190_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net242));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[12]$_DFFE_PN0P_  (.D(_00191_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net243));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[13]$_DFFE_PN0P_  (.D(_00192_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net244));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[14]$_DFFE_PN0P_  (.D(_00193_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net245));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[15]$_DFFE_PN0P_  (.D(_00194_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net246));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[16]$_DFFE_PN0P_  (.D(_00195_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net247));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[17]$_DFFE_PN0P_  (.D(_00196_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net248));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[18]$_DFFE_PN0P_  (.D(_00197_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net249));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[19]$_DFFE_PN0P_  (.D(_00198_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net250));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[1]$_DFFE_PN0P_  (.D(_00199_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net251));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[20]$_DFFE_PN0P_  (.D(_00200_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net252));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[21]$_DFFE_PN0P_  (.D(_00201_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net253));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[22]$_DFFE_PN0P_  (.D(_00202_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net254));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[23]$_DFFE_PN0P_  (.D(_00203_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net255));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[24]$_DFFE_PN0P_  (.D(_00204_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net256));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[25]$_DFFE_PN0P_  (.D(_00205_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net257));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[26]$_DFFE_PN0P_  (.D(_00206_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net258));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[27]$_DFFE_PN0P_  (.D(_00207_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net259));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[28]$_DFFE_PN0P_  (.D(_00208_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net260));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[29]$_DFFE_PN0P_  (.D(_00209_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net261));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[2]$_DFFE_PN0P_  (.D(_00210_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net262));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[30]$_DFFE_PN0P_  (.D(_00211_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net263));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[31]$_DFFE_PN0P_  (.D(_00212_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net264));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[32]$_DFFE_PN0P_  (.D(_00213_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net265));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[33]$_DFFE_PN0P_  (.D(_00214_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net266));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[34]$_DFFE_PN0P_  (.D(_00215_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net267));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[35]$_DFFE_PN0P_  (.D(_00216_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net268));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[36]$_DFFE_PN0P_  (.D(_00217_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net269));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[37]$_DFFE_PN0P_  (.D(_00218_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net270));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[38]$_DFFE_PN0P_  (.D(_00219_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net271));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[39]$_DFFE_PN0P_  (.D(_00220_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net272));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[3]$_DFFE_PN0P_  (.D(_00221_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net273));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[40]$_DFFE_PN0P_  (.D(_00222_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net274));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[41]$_DFFE_PN0P_  (.D(_00223_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net275));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[42]$_DFFE_PN0P_  (.D(_00224_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net276));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[43]$_DFFE_PN0P_  (.D(_00225_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net277));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[44]$_DFFE_PN0P_  (.D(_00226_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net278));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[45]$_DFFE_PN0P_  (.D(_00227_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net279));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[46]$_DFFE_PN0P_  (.D(_00228_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net280));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[47]$_DFFE_PN0P_  (.D(_00229_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(net281));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[48]$_DFFE_PN0P_  (.D(_00230_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(net282));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[49]$_DFFE_PN0P_  (.D(_00231_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net283));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[4]$_DFFE_PN0P_  (.D(_00232_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net284));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[50]$_DFFE_PN0P_  (.D(_00233_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net285));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[51]$_DFFE_PN0P_  (.D(_00234_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net286));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[52]$_DFFE_PN0P_  (.D(_00235_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net287));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[53]$_DFFE_PN0P_  (.D(_00236_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net288));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[54]$_DFFE_PN0P_  (.D(_00237_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net289));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[55]$_DFFE_PN0P_  (.D(_00238_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net290));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[56]$_DFFE_PN0P_  (.D(_00239_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net291));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[57]$_DFFE_PN0P_  (.D(_00240_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net292));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[58]$_DFFE_PN0P_  (.D(_00241_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net293));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[59]$_DFFE_PN0P_  (.D(_00242_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net294));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[5]$_DFFE_PN0P_  (.D(_00243_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net295));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[60]$_DFFE_PN0P_  (.D(_00244_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net296));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[61]$_DFFE_PN0P_  (.D(_00245_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net297));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[62]$_DFFE_PN0P_  (.D(_00246_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net298));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[63]$_DFFE_PN0P_  (.D(_00247_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net299));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[64]$_DFFE_PN0P_  (.D(_00248_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(net300));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[65]$_DFFE_PN0P_  (.D(_00249_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net301));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[66]$_DFFE_PN0P_  (.D(_00250_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net302));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[67]$_DFFE_PN0P_  (.D(_00251_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net303));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[68]$_DFFE_PN0P_  (.D(_00252_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net304));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[69]$_DFFE_PN0P_  (.D(_00253_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net305));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[6]$_DFFE_PN0P_  (.D(_00254_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net306));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[70]$_DFFE_PN0P_  (.D(_00255_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(net307));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[71]$_DFFE_PN0P_  (.D(_00256_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net308));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[72]$_DFFE_PN0P_  (.D(_00257_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net309));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[73]$_DFFE_PN0P_  (.D(_00258_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net310));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[74]$_DFFE_PN0P_  (.D(_00259_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net311));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[75]$_DFFE_PN0P_  (.D(_00260_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net312));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[76]$_DFFE_PN0P_  (.D(_00261_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net313));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[77]$_DFFE_PN0P_  (.D(_00262_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(net314));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[78]$_DFFE_PN0P_  (.D(_00263_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net315));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[79]$_DFFE_PN0P_  (.D(_00264_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net316));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[7]$_DFFE_PN0P_  (.D(_00265_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net317));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[80]$_DFFE_PN0P_  (.D(_00266_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(net318));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[81]$_DFFE_PN0P_  (.D(_00267_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net319));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[82]$_DFFE_PN0P_  (.D(_00268_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net320));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[83]$_DFFE_PN0P_  (.D(_00269_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net321));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[84]$_DFFE_PN0P_  (.D(_00270_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(net322));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[85]$_DFFE_PN0P_  (.D(_00271_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net323));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[86]$_DFFE_PN0P_  (.D(_00272_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net324));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[87]$_DFFE_PN0P_  (.D(_00273_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net325));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[88]$_DFFE_PN0P_  (.D(_00274_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(net326));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[89]$_DFFE_PN0P_  (.D(_00275_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net327));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[8]$_DFFE_PN0P_  (.D(_00276_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(net328));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[90]$_DFFE_PN0P_  (.D(_00277_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net329));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[91]$_DFFE_PN0P_  (.D(_00278_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(net330));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[92]$_DFFE_PN0P_  (.D(_00279_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net331));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[93]$_DFFE_PN0P_  (.D(_00280_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net332));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[94]$_DFFE_PN0P_  (.D(_00281_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net333));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[95]$_DFFE_PN0P_  (.D(_00282_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(net334));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[96]$_DFFE_PN0P_  (.D(_00283_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(net335));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[97]$_DFFE_PN0P_  (.D(_00284_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net336));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[98]$_DFFE_PN0P_  (.D(_00285_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(net337));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[99]$_DFFE_PN0P_  (.D(_00286_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net338));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out_real[9]$_DFFE_PN0P_  (.D(_00287_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(net339));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \data_ready$_DFFE_PN1P_  (.D(_00288_),
    .SETN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(net340));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_valid_out$_DFFE_PN0P_  (.D(_00289_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(net341));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \group[0]$_DFFE_PP_  (.D(_00290_),
    .CLK(clknet_leaf_20_clk),
    .Q(\group[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \group[1]$_DFFE_PP_  (.D(_00291_),
    .CLK(clknet_leaf_20_clk),
    .Q(\group[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \group[2]$_DFFE_PP_  (.D(_00292_),
    .CLK(clknet_leaf_20_clk),
    .Q(\group[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \idx1[0]$_DFFE_PP_  (.D(_00293_),
    .CLK(clknet_leaf_17_clk),
    .Q(\idx1[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \idx1[1]$_DFFE_PP_  (.D(_00294_),
    .CLK(clknet_leaf_17_clk),
    .Q(\idx1[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \idx1[2]$_DFFE_PP_  (.D(_00295_),
    .CLK(clknet_leaf_9_clk),
    .Q(\idx1[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \idx2[0]$_DFFE_PP_  (.D(_00296_),
    .CLK(clknet_leaf_9_clk),
    .Q(\idx2[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \idx2[1]$_DFFE_PP_  (.D(_00297_),
    .CLK(clknet_leaf_9_clk),
    .Q(\idx2[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \idx2[2]$_DFFE_PP_  (.D(_00298_),
    .CLK(clknet_leaf_17_clk),
    .Q(\idx2[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \sample_count[0]$_DFFE_PN0P_  (.D(_00299_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\sample_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \sample_count[1]$_DFFE_PN0P_  (.D(_00300_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\sample_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \sample_count[2]$_DFFE_PN0P_  (.D(_00301_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\sample_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][0]$_DFFE_PN0P_  (.D(_00302_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][10]$_DFFE_PN0P_  (.D(_00303_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_imag[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][11]$_DFFE_PN0P_  (.D(_00304_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_imag[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][12]$_DFFE_PN0P_  (.D(_00305_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][13]$_DFFE_PN0P_  (.D(_00306_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][14]$_DFFE_PN0P_  (.D(_00307_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][15]$_DFFE_PN0P_  (.D(_00308_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][1]$_DFFE_PN0P_  (.D(_00309_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][2]$_DFFE_PN0P_  (.D(_00310_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][3]$_DFFE_PN0P_  (.D(_00311_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][4]$_DFFE_PN0P_  (.D(_00312_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][5]$_DFFE_PN0P_  (.D(_00313_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][6]$_DFFE_PN0P_  (.D(_00314_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][7]$_DFFE_PN0P_  (.D(_00315_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][8]$_DFFE_PN0P_  (.D(_00316_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[0][9]$_DFFE_PN0P_  (.D(_00317_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][0]$_DFFE_PN0P_  (.D(_00318_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][10]$_DFFE_PN0P_  (.D(_00319_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][11]$_DFFE_PN0P_  (.D(_00320_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][12]$_DFFE_PN0P_  (.D(_00321_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][13]$_DFFE_PN0P_  (.D(_00322_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][14]$_DFFE_PN0P_  (.D(_00323_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][15]$_DFFE_PN0P_  (.D(_00324_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][1]$_DFFE_PN0P_  (.D(_00325_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][2]$_DFFE_PN0P_  (.D(_00326_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][3]$_DFFE_PN0P_  (.D(_00327_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][4]$_DFFE_PN0P_  (.D(_00328_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][5]$_DFFE_PN0P_  (.D(_00329_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][6]$_DFFE_PN0P_  (.D(_00330_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][7]$_DFFE_PN0P_  (.D(_00331_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][8]$_DFFE_PN0P_  (.D(_00332_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[1][9]$_DFFE_PN0P_  (.D(_00333_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][0]$_DFFE_PN0P_  (.D(_00334_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][10]$_DFFE_PN0P_  (.D(_00335_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][11]$_DFFE_PN0P_  (.D(_00336_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][12]$_DFFE_PN0P_  (.D(_00337_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][13]$_DFFE_PN0P_  (.D(_00338_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][14]$_DFFE_PN0P_  (.D(_00339_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][15]$_DFFE_PN0P_  (.D(_00340_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][1]$_DFFE_PN0P_  (.D(_00341_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][2]$_DFFE_PN0P_  (.D(_00342_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][3]$_DFFE_PN0P_  (.D(_00343_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][4]$_DFFE_PN0P_  (.D(_00344_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][5]$_DFFE_PN0P_  (.D(_00345_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][6]$_DFFE_PN0P_  (.D(_00346_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][7]$_DFFE_PN0P_  (.D(_00347_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][8]$_DFFE_PN0P_  (.D(_00348_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[2][9]$_DFFE_PN0P_  (.D(_00349_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][0]$_DFFE_PN0P_  (.D(_00350_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][10]$_DFFE_PN0P_  (.D(_00351_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][11]$_DFFE_PN0P_  (.D(_00352_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][12]$_DFFE_PN0P_  (.D(_00353_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][13]$_DFFE_PN0P_  (.D(_00354_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][14]$_DFFE_PN0P_  (.D(_00355_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][15]$_DFFE_PN0P_  (.D(_00356_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][1]$_DFFE_PN0P_  (.D(_00357_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][2]$_DFFE_PN0P_  (.D(_00358_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][3]$_DFFE_PN0P_  (.D(_00359_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][4]$_DFFE_PN0P_  (.D(_00360_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][5]$_DFFE_PN0P_  (.D(_00361_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][6]$_DFFE_PN0P_  (.D(_00362_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][7]$_DFFE_PN0P_  (.D(_00363_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][8]$_DFFE_PN0P_  (.D(_00364_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_imag[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[3][9]$_DFFE_PN0P_  (.D(_00365_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_imag[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][0]$_DFFE_PN0P_  (.D(_00366_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][10]$_DFFE_PN0P_  (.D(_00367_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][11]$_DFFE_PN0P_  (.D(_00368_),
    .RN(net81),
    .CLK(clknet_leaf_15_clk),
    .Q(\samples_imag[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][12]$_DFFE_PN0P_  (.D(_00369_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][13]$_DFFE_PN0P_  (.D(_00370_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][14]$_DFFE_PN0P_  (.D(_00371_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][15]$_DFFE_PN0P_  (.D(_00372_),
    .RN(net81),
    .CLK(clknet_leaf_19_clk),
    .Q(\samples_imag[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][1]$_DFFE_PN0P_  (.D(_00373_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][2]$_DFFE_PN0P_  (.D(_00374_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][3]$_DFFE_PN0P_  (.D(_00375_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][4]$_DFFE_PN0P_  (.D(_00376_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][5]$_DFFE_PN0P_  (.D(_00377_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][6]$_DFFE_PN0P_  (.D(_00378_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][7]$_DFFE_PN0P_  (.D(_00379_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][8]$_DFFE_PN0P_  (.D(_00380_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[4][9]$_DFFE_PN0P_  (.D(_00381_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][0]$_DFFE_PN0P_  (.D(_00382_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][10]$_DFFE_PN0P_  (.D(_00383_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][11]$_DFFE_PN0P_  (.D(_00384_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][12]$_DFFE_PN0P_  (.D(_00385_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][13]$_DFFE_PN0P_  (.D(_00386_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][14]$_DFFE_PN0P_  (.D(_00387_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][15]$_DFFE_PN0P_  (.D(_00388_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][1]$_DFFE_PN0P_  (.D(_00389_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][2]$_DFFE_PN0P_  (.D(_00390_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][3]$_DFFE_PN0P_  (.D(_00391_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][4]$_DFFE_PN0P_  (.D(_00392_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][5]$_DFFE_PN0P_  (.D(_00393_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][6]$_DFFE_PN0P_  (.D(_00394_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][7]$_DFFE_PN0P_  (.D(_00395_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][8]$_DFFE_PN0P_  (.D(_00396_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[5][9]$_DFFE_PN0P_  (.D(_00397_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][0]$_DFFE_PN0P_  (.D(_00398_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][10]$_DFFE_PN0P_  (.D(_00399_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][11]$_DFFE_PN0P_  (.D(_00400_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][12]$_DFFE_PN0P_  (.D(_00401_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][13]$_DFFE_PN0P_  (.D(_00402_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][14]$_DFFE_PN0P_  (.D(_00403_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][15]$_DFFE_PN0P_  (.D(_00404_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][1]$_DFFE_PN0P_  (.D(_00405_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][2]$_DFFE_PN0P_  (.D(_00406_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][3]$_DFFE_PN0P_  (.D(_00407_),
    .RN(net81),
    .CLK(clknet_leaf_13_clk),
    .Q(\samples_imag[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][4]$_DFFE_PN0P_  (.D(_00408_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][5]$_DFFE_PN0P_  (.D(_00409_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][6]$_DFFE_PN0P_  (.D(_00410_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][7]$_DFFE_PN0P_  (.D(_00411_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][8]$_DFFE_PN0P_  (.D(_00412_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_imag[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[6][9]$_DFFE_PN0P_  (.D(_00413_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_imag[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][0]$_DFFE_PN0P_  (.D(_00414_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][10]$_DFFE_PN0P_  (.D(_00415_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_imag[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][11]$_DFFE_PN0P_  (.D(_00416_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][12]$_DFFE_PN0P_  (.D(_00417_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][13]$_DFFE_PN0P_  (.D(_00418_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][14]$_DFFE_PN0P_  (.D(_00419_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_imag[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][15]$_DFFE_PN0P_  (.D(_00420_),
    .RN(net81),
    .CLK(clknet_leaf_18_clk),
    .Q(\samples_imag[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][1]$_DFFE_PN0P_  (.D(_00421_),
    .RN(net81),
    .CLK(clknet_leaf_16_clk),
    .Q(\samples_imag[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][2]$_DFFE_PN0P_  (.D(_00422_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][3]$_DFFE_PN0P_  (.D(_00423_),
    .RN(net81),
    .CLK(clknet_leaf_14_clk),
    .Q(\samples_imag[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][4]$_DFFE_PN0P_  (.D(_00424_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][5]$_DFFE_PN0P_  (.D(_00425_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][6]$_DFFE_PN0P_  (.D(_00426_),
    .RN(net81),
    .CLK(clknet_leaf_12_clk),
    .Q(\samples_imag[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][7]$_DFFE_PN0P_  (.D(_00427_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][8]$_DFFE_PN0P_  (.D(_00428_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_imag[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_imag[7][9]$_DFFE_PN0P_  (.D(_00429_),
    .RN(net81),
    .CLK(clknet_leaf_11_clk),
    .Q(\samples_imag[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \samples_real[0][0]$_DFFE_PN0P_  (.D(_00430_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_real[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][10]$_DFFE_PN0P_  (.D(_00431_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_real[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][11]$_DFFE_PN0P_  (.D(_00432_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_real[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][12]$_DFFE_PN0P_  (.D(_00433_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][13]$_DFFE_PN0P_  (.D(_00434_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][14]$_DFFE_PN0P_  (.D(_00435_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][15]$_DFFE_PN0P_  (.D(_00436_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][1]$_DFFE_PN0P_  (.D(_00437_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][2]$_DFFE_PN0P_  (.D(_00438_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][3]$_DFFE_PN0P_  (.D(_00439_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][4]$_DFFE_PN0P_  (.D(_00440_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][5]$_DFFE_PN0P_  (.D(_00441_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][6]$_DFFE_PN0P_  (.D(_00442_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][7]$_DFFE_PN0P_  (.D(_00443_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][8]$_DFFE_PN0P_  (.D(_00444_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[0][9]$_DFFE_PN0P_  (.D(_00445_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][0]$_DFFE_PN0P_  (.D(_00446_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][10]$_DFFE_PN0P_  (.D(_00447_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][11]$_DFFE_PN0P_  (.D(_00448_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][12]$_DFFE_PN0P_  (.D(_00449_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][13]$_DFFE_PN0P_  (.D(_00450_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][14]$_DFFE_PN0P_  (.D(_00451_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][15]$_DFFE_PN0P_  (.D(_00452_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][1]$_DFFE_PN0P_  (.D(_00453_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][2]$_DFFE_PN0P_  (.D(_00454_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][3]$_DFFE_PN0P_  (.D(_00455_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][4]$_DFFE_PN0P_  (.D(_00456_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][5]$_DFFE_PN0P_  (.D(_00457_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][6]$_DFFE_PN0P_  (.D(_00458_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][7]$_DFFE_PN0P_  (.D(_00459_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][8]$_DFFE_PN0P_  (.D(_00460_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[1][9]$_DFFE_PN0P_  (.D(_00461_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \samples_real[2][0]$_DFFE_PN0P_  (.D(_00462_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_real[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][10]$_DFFE_PN0P_  (.D(_00463_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][11]$_DFFE_PN0P_  (.D(_00464_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][12]$_DFFE_PN0P_  (.D(_00465_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][13]$_DFFE_PN0P_  (.D(_00466_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][14]$_DFFE_PN0P_  (.D(_00467_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][15]$_DFFE_PN0P_  (.D(_00468_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][1]$_DFFE_PN0P_  (.D(_00469_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][2]$_DFFE_PN0P_  (.D(_00470_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][3]$_DFFE_PN0P_  (.D(_00471_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][4]$_DFFE_PN0P_  (.D(_00472_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][5]$_DFFE_PN0P_  (.D(_00473_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][6]$_DFFE_PN0P_  (.D(_00474_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][7]$_DFFE_PN0P_  (.D(_00475_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(\samples_real[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][8]$_DFFE_PN0P_  (.D(_00476_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[2][9]$_DFFE_PN0P_  (.D(_00477_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][0]$_DFFE_PN0P_  (.D(_00478_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][10]$_DFFE_PN0P_  (.D(_00479_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_real[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][11]$_DFFE_PN0P_  (.D(_00480_),
    .RN(net81),
    .CLK(clknet_leaf_9_clk),
    .Q(\samples_real[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][12]$_DFFE_PN0P_  (.D(_00481_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][13]$_DFFE_PN0P_  (.D(_00482_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][14]$_DFFE_PN0P_  (.D(_00483_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][15]$_DFFE_PN0P_  (.D(_00484_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][1]$_DFFE_PN0P_  (.D(_00485_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][2]$_DFFE_PN0P_  (.D(_00486_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][3]$_DFFE_PN0P_  (.D(_00487_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][4]$_DFFE_PN0P_  (.D(_00488_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][5]$_DFFE_PN0P_  (.D(_00489_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][6]$_DFFE_PN0P_  (.D(_00490_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][7]$_DFFE_PN0P_  (.D(_00491_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][8]$_DFFE_PN0P_  (.D(_00492_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[3][9]$_DFFE_PN0P_  (.D(_00493_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][0]$_DFFE_PN0P_  (.D(_00494_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \samples_real[4][10]$_DFFE_PN0P_  (.D(_00495_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][11]$_DFFE_PN0P_  (.D(_00496_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][12]$_DFFE_PN0P_  (.D(_00497_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][13]$_DFFE_PN0P_  (.D(_00498_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][14]$_DFFE_PN0P_  (.D(_00499_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][15]$_DFFE_PN0P_  (.D(_00500_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][1]$_DFFE_PN0P_  (.D(_00501_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][2]$_DFFE_PN0P_  (.D(_00502_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][3]$_DFFE_PN0P_  (.D(_00503_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][4]$_DFFE_PN0P_  (.D(_00504_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][5]$_DFFE_PN0P_  (.D(_00505_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][6]$_DFFE_PN0P_  (.D(_00506_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][7]$_DFFE_PN0P_  (.D(_00507_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][8]$_DFFE_PN0P_  (.D(_00508_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[4][9]$_DFFE_PN0P_  (.D(_00509_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][0]$_DFFE_PN0P_  (.D(_00510_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][10]$_DFFE_PN0P_  (.D(_00511_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][11]$_DFFE_PN0P_  (.D(_00512_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][12]$_DFFE_PN0P_  (.D(_00513_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][13]$_DFFE_PN0P_  (.D(_00514_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][14]$_DFFE_PN0P_  (.D(_00515_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][15]$_DFFE_PN0P_  (.D(_00516_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][1]$_DFFE_PN0P_  (.D(_00517_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][2]$_DFFE_PN0P_  (.D(_00518_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][3]$_DFFE_PN0P_  (.D(_00519_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][4]$_DFFE_PN0P_  (.D(_00520_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][5]$_DFFE_PN0P_  (.D(_00521_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][6]$_DFFE_PN0P_  (.D(_00522_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][7]$_DFFE_PN0P_  (.D(_00523_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][8]$_DFFE_PN0P_  (.D(_00524_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[5][9]$_DFFE_PN0P_  (.D(_00525_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][0]$_DFFE_PN0P_  (.D(_00526_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][10]$_DFFE_PN0P_  (.D(_00527_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][11]$_DFFE_PN0P_  (.D(_00528_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][12]$_DFFE_PN0P_  (.D(_00529_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][13]$_DFFE_PN0P_  (.D(_00530_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][14]$_DFFE_PN0P_  (.D(_00531_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][15]$_DFFE_PN0P_  (.D(_00532_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][1]$_DFFE_PN0P_  (.D(_00533_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][2]$_DFFE_PN0P_  (.D(_00534_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][3]$_DFFE_PN0P_  (.D(_00535_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][4]$_DFFE_PN0P_  (.D(_00536_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][5]$_DFFE_PN0P_  (.D(_00537_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][6]$_DFFE_PN0P_  (.D(_00538_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][7]$_DFFE_PN0P_  (.D(_00539_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][8]$_DFFE_PN0P_  (.D(_00540_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[6][9]$_DFFE_PN0P_  (.D(_00541_),
    .RN(net81),
    .CLK(clknet_leaf_4_clk),
    .Q(\samples_real[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][0]$_DFFE_PN0P_  (.D(_00542_),
    .RN(net81),
    .CLK(clknet_leaf_17_clk),
    .Q(\samples_real[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][10]$_DFFE_PN0P_  (.D(_00543_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][11]$_DFFE_PN0P_  (.D(_00544_),
    .RN(net81),
    .CLK(clknet_leaf_10_clk),
    .Q(\samples_real[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][12]$_DFFE_PN0P_  (.D(_00545_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][13]$_DFFE_PN0P_  (.D(_00546_),
    .RN(net81),
    .CLK(clknet_leaf_7_clk),
    .Q(\samples_real[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][14]$_DFFE_PN0P_  (.D(_00547_),
    .RN(net81),
    .CLK(clknet_leaf_6_clk),
    .Q(\samples_real[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][15]$_DFFE_PN0P_  (.D(_00548_),
    .RN(net81),
    .CLK(clknet_leaf_8_clk),
    .Q(\samples_real[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][1]$_DFFE_PN0P_  (.D(_00549_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][2]$_DFFE_PN0P_  (.D(_00550_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][3]$_DFFE_PN0P_  (.D(_00551_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][4]$_DFFE_PN0P_  (.D(_00552_),
    .RN(net81),
    .CLK(clknet_leaf_0_clk),
    .Q(\samples_real[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][5]$_DFFE_PN0P_  (.D(_00553_),
    .RN(net81),
    .CLK(clknet_leaf_1_clk),
    .Q(\samples_real[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][6]$_DFFE_PN0P_  (.D(_00554_),
    .RN(net81),
    .CLK(clknet_leaf_2_clk),
    .Q(\samples_real[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][7]$_DFFE_PN0P_  (.D(_00555_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(\samples_real[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][8]$_DFFE_PN0P_  (.D(_00556_),
    .RN(net81),
    .CLK(clknet_leaf_3_clk),
    .Q(\samples_real[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \samples_real[7][9]$_DFFE_PN0P_  (.D(_00557_),
    .RN(net81),
    .CLK(clknet_leaf_5_clk),
    .Q(\samples_real[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \stage[0]$_DFFE_PN0P_  (.D(_00558_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\stage[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \stage[1]$_DFFE_PN0P_  (.D(_00559_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\stage[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \stage[2]$_DFFE_PN0P_  (.D(_00560_),
    .RN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\stage[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \state[0]$_DFF_PN1_  (.D(_00004_),
    .SETN(net81),
    .CLK(clknet_leaf_20_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFF_PN0_  (.D(_00005_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[2]$_DFF_PN0_  (.D(_00006_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[3]$_DFF_PN0_  (.D(_00003_),
    .RN(net81),
    .CLK(clknet_leaf_21_clk),
    .Q(\state[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \temp_imag[0]$_DFFE_PP_  (.D(_00561_),
    .CLK(clknet_leaf_17_clk),
    .Q(\temp_imag[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \temp_real[0]$_DFFE_PP_  (.D(_00562_),
    .CLK(clknet_leaf_0_clk),
    .Q(\temp_real[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \twiddle_idx[0]$_DFFE_PP_  (.D(_00000_),
    .CLK(clknet_leaf_20_clk),
    .Q(\twiddle_idx[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \twiddle_idx[1]$_DFFE_PP_  (.D(_00007_),
    .CLK(clknet_leaf_20_clk),
    .Q(\twiddle_idx[1] ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone1 (.A1(net26),
    .A2(_07787_),
    .ZN(net1));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone2 (.A1(net26),
    .A2(_00567_),
    .ZN(net2));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 clone3 (.A1(net15),
    .A2(_02443_),
    .A3(_02478_),
    .A4(_02501_),
    .ZN(net3));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 clone4 (.A1(_02349_),
    .A2(_02310_),
    .ZN(net4));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 clone5 (.A1(_00608_),
    .A2(_00606_),
    .B1(_00613_),
    .B2(_00614_),
    .C(_00615_),
    .ZN(net5));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 clone6 (.A1(net21),
    .A2(_01039_),
    .A3(_00913_),
    .ZN(net6));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone7 (.A1(_02632_),
    .A2(_02630_),
    .B(_02633_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone8 (.A1(net26),
    .A2(_07787_),
    .ZN(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 clone9 (.I(_01982_),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 clone10 (.A1(_03416_),
    .A2(_03364_),
    .A3(_03345_),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clone11 (.I(_02636_),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clone12 (.I(_03005_),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 clone13 (.I(_01488_),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 clone14 (.I(_02548_),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone15 (.A1(_02458_),
    .A2(_02455_),
    .ZN(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 clone16 (.I(_03556_),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone17 (.I(_01928_),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clone18 (.I(_00582_),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone19 (.A1(net26),
    .A2(_00567_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 clone20 (.A1(_01972_),
    .A2(_01980_),
    .A3(_01977_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 split21 (.I(_07223_),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone22 (.I(_01486_),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone23 (.A1(_02637_),
    .A2(_02590_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone24 (.I(_02403_),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone25 (.A1(_02402_),
    .A2(_02350_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 split26 (.I(_07775_),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone27 (.I(_01747_),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone28 (.I(_01186_),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone29 (.I(_02700_),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone30 (.I(_01634_),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 clone32 (.I(_01294_),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 clone33 (.A1(_00772_),
    .A2(_00762_),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 clone34 (.A1(_07104_),
    .A2(_00737_),
    .B(_00771_),
    .C(_00770_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone35 (.I(_02843_),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone36 (.I(_07794_),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone37 (.I(net390),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone38 (.I(_01343_),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone39 (.I(_03107_),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone41 (.I(_02841_),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone42 (.I(_01276_),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone43 (.I(_02201_),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone44 (.I(_02275_),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone45 (.I(_02549_),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone46 (.I(net375),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone47 (.I(_03108_),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input1 (.I(data_in_imag[0]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input2 (.I(data_in_imag[10]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input3 (.I(data_in_imag[11]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input4 (.I(data_in_imag[12]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input5 (.I(data_in_imag[13]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input6 (.I(data_in_imag[14]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input7 (.I(data_in_imag[15]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input8 (.I(data_in_imag[1]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input9 (.I(data_in_imag[2]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input10 (.I(data_in_imag[3]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input11 (.I(data_in_imag[4]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input12 (.I(data_in_imag[5]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input13 (.I(data_in_imag[6]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input14 (.I(data_in_imag[7]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input15 (.I(data_in_imag[8]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input16 (.I(data_in_imag[9]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input17 (.I(data_in_real[0]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input18 (.I(data_in_real[10]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input19 (.I(data_in_real[11]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input20 (.I(data_in_real[12]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input21 (.I(data_in_real[13]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input22 (.I(data_in_real[14]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input23 (.I(data_in_real[15]),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input24 (.I(data_in_real[1]),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input25 (.I(data_in_real[2]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input26 (.I(data_in_real[3]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input27 (.I(data_in_real[4]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input28 (.I(data_in_real[5]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input29 (.I(data_in_real[6]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input30 (.I(data_in_real[7]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input31 (.I(data_in_real[8]),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input32 (.I(data_in_real[9]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input33 (.I(data_valid_in),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input34 (.I(rst_n),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input35 (.I(start),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output36 (.I(net83),
    .Z(busy));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net84),
    .Z(data_out_imag[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net85),
    .Z(data_out_imag[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net86),
    .Z(data_out_imag[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net87),
    .Z(data_out_imag[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net88),
    .Z(data_out_imag[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net89),
    .Z(data_out_imag[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net90),
    .Z(data_out_imag[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net91),
    .Z(data_out_imag[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net92),
    .Z(data_out_imag[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net93),
    .Z(data_out_imag[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net94),
    .Z(data_out_imag[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net95),
    .Z(data_out_imag[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net96),
    .Z(data_out_imag[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net97),
    .Z(data_out_imag[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net98),
    .Z(data_out_imag[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net99),
    .Z(data_out_imag[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net100),
    .Z(data_out_imag[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net101),
    .Z(data_out_imag[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net102),
    .Z(data_out_imag[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net103),
    .Z(data_out_imag[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net104),
    .Z(data_out_imag[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net105),
    .Z(data_out_imag[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net106),
    .Z(data_out_imag[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net107),
    .Z(data_out_imag[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net108),
    .Z(data_out_imag[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net109),
    .Z(data_out_imag[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net110),
    .Z(data_out_imag[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net111),
    .Z(data_out_imag[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net112),
    .Z(data_out_imag[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net113),
    .Z(data_out_imag[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net114),
    .Z(data_out_imag[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net115),
    .Z(data_out_imag[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net116),
    .Z(data_out_imag[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net117),
    .Z(data_out_imag[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net118),
    .Z(data_out_imag[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net119),
    .Z(data_out_imag[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net120),
    .Z(data_out_imag[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net121),
    .Z(data_out_imag[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net122),
    .Z(data_out_imag[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net123),
    .Z(data_out_imag[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net124),
    .Z(data_out_imag[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net125),
    .Z(data_out_imag[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net126),
    .Z(data_out_imag[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net127),
    .Z(data_out_imag[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net128),
    .Z(data_out_imag[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net129),
    .Z(data_out_imag[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net130),
    .Z(data_out_imag[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net131),
    .Z(data_out_imag[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net132),
    .Z(data_out_imag[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net133),
    .Z(data_out_imag[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net134),
    .Z(data_out_imag[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net135),
    .Z(data_out_imag[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net136),
    .Z(data_out_imag[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net137),
    .Z(data_out_imag[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net138),
    .Z(data_out_imag[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net139),
    .Z(data_out_imag[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net140),
    .Z(data_out_imag[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net141),
    .Z(data_out_imag[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net142),
    .Z(data_out_imag[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net143),
    .Z(data_out_imag[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net144),
    .Z(data_out_imag[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net145),
    .Z(data_out_imag[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net146),
    .Z(data_out_imag[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net147),
    .Z(data_out_imag[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net148),
    .Z(data_out_imag[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net149),
    .Z(data_out_imag[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net150),
    .Z(data_out_imag[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net151),
    .Z(data_out_imag[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net152),
    .Z(data_out_imag[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net153),
    .Z(data_out_imag[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net154),
    .Z(data_out_imag[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net155),
    .Z(data_out_imag[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net156),
    .Z(data_out_imag[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net157),
    .Z(data_out_imag[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net158),
    .Z(data_out_imag[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output112 (.I(net159),
    .Z(data_out_imag[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output113 (.I(net160),
    .Z(data_out_imag[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output114 (.I(net161),
    .Z(data_out_imag[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output115 (.I(net162),
    .Z(data_out_imag[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output116 (.I(net163),
    .Z(data_out_imag[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output117 (.I(net164),
    .Z(data_out_imag[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output118 (.I(net165),
    .Z(data_out_imag[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output119 (.I(net166),
    .Z(data_out_imag[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output120 (.I(net167),
    .Z(data_out_imag[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output121 (.I(net168),
    .Z(data_out_imag[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output122 (.I(net169),
    .Z(data_out_imag[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output123 (.I(net170),
    .Z(data_out_imag[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output124 (.I(net171),
    .Z(data_out_imag[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output125 (.I(net172),
    .Z(data_out_imag[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output126 (.I(net173),
    .Z(data_out_imag[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output127 (.I(net174),
    .Z(data_out_imag[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output128 (.I(net175),
    .Z(data_out_imag[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output129 (.I(net176),
    .Z(data_out_imag[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output130 (.I(net177),
    .Z(data_out_imag[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output131 (.I(net178),
    .Z(data_out_imag[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output132 (.I(net179),
    .Z(data_out_imag[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output133 (.I(net180),
    .Z(data_out_imag[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output134 (.I(net181),
    .Z(data_out_imag[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output135 (.I(net182),
    .Z(data_out_imag[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output136 (.I(net183),
    .Z(data_out_imag[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output137 (.I(net184),
    .Z(data_out_imag[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output138 (.I(net185),
    .Z(data_out_imag[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output139 (.I(net186),
    .Z(data_out_imag[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output140 (.I(net187),
    .Z(data_out_imag[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output141 (.I(net188),
    .Z(data_out_imag[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output142 (.I(net189),
    .Z(data_out_imag[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output143 (.I(net190),
    .Z(data_out_imag[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output144 (.I(net191),
    .Z(data_out_imag[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net192),
    .Z(data_out_imag[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output146 (.I(net193),
    .Z(data_out_imag[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output147 (.I(net194),
    .Z(data_out_imag[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output148 (.I(net195),
    .Z(data_out_imag[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output149 (.I(net196),
    .Z(data_out_imag[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output150 (.I(net197),
    .Z(data_out_imag[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output151 (.I(net198),
    .Z(data_out_imag[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output152 (.I(net199),
    .Z(data_out_imag[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output153 (.I(net200),
    .Z(data_out_imag[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output154 (.I(net201),
    .Z(data_out_imag[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output155 (.I(net202),
    .Z(data_out_imag[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net203),
    .Z(data_out_imag[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net204),
    .Z(data_out_imag[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net205),
    .Z(data_out_imag[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net206),
    .Z(data_out_imag[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output160 (.I(net207),
    .Z(data_out_imag[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net208),
    .Z(data_out_imag[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net209),
    .Z(data_out_imag[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net210),
    .Z(data_out_imag[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net211),
    .Z(data_out_imag[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net212),
    .Z(data_out_real[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net213),
    .Z(data_out_real[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net214),
    .Z(data_out_real[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net215),
    .Z(data_out_real[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net216),
    .Z(data_out_real[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net217),
    .Z(data_out_real[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net218),
    .Z(data_out_real[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net219),
    .Z(data_out_real[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net220),
    .Z(data_out_real[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output174 (.I(net221),
    .Z(data_out_real[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output175 (.I(net222),
    .Z(data_out_real[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output176 (.I(net223),
    .Z(data_out_real[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output177 (.I(net224),
    .Z(data_out_real[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output178 (.I(net225),
    .Z(data_out_real[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output179 (.I(net226),
    .Z(data_out_real[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output180 (.I(net227),
    .Z(data_out_real[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output181 (.I(net228),
    .Z(data_out_real[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output182 (.I(net229),
    .Z(data_out_real[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output183 (.I(net230),
    .Z(data_out_real[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output184 (.I(net231),
    .Z(data_out_real[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output185 (.I(net232),
    .Z(data_out_real[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output186 (.I(net233),
    .Z(data_out_real[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output187 (.I(net234),
    .Z(data_out_real[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output188 (.I(net235),
    .Z(data_out_real[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output189 (.I(net236),
    .Z(data_out_real[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output190 (.I(net237),
    .Z(data_out_real[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output191 (.I(net238),
    .Z(data_out_real[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output192 (.I(net239),
    .Z(data_out_real[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output193 (.I(net240),
    .Z(data_out_real[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output194 (.I(net241),
    .Z(data_out_real[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output195 (.I(net242),
    .Z(data_out_real[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output196 (.I(net243),
    .Z(data_out_real[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output197 (.I(net244),
    .Z(data_out_real[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output198 (.I(net245),
    .Z(data_out_real[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output199 (.I(net246),
    .Z(data_out_real[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output200 (.I(net247),
    .Z(data_out_real[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output201 (.I(net248),
    .Z(data_out_real[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output202 (.I(net249),
    .Z(data_out_real[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output203 (.I(net250),
    .Z(data_out_real[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output204 (.I(net251),
    .Z(data_out_real[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output205 (.I(net252),
    .Z(data_out_real[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output206 (.I(net253),
    .Z(data_out_real[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output207 (.I(net254),
    .Z(data_out_real[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output208 (.I(net255),
    .Z(data_out_real[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output209 (.I(net256),
    .Z(data_out_real[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output210 (.I(net257),
    .Z(data_out_real[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output211 (.I(net258),
    .Z(data_out_real[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output212 (.I(net259),
    .Z(data_out_real[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output213 (.I(net260),
    .Z(data_out_real[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output214 (.I(net261),
    .Z(data_out_real[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output215 (.I(net262),
    .Z(data_out_real[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output216 (.I(net263),
    .Z(data_out_real[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output217 (.I(net264),
    .Z(data_out_real[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output218 (.I(net265),
    .Z(data_out_real[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output219 (.I(net266),
    .Z(data_out_real[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output220 (.I(net267),
    .Z(data_out_real[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output221 (.I(net268),
    .Z(data_out_real[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output222 (.I(net269),
    .Z(data_out_real[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output223 (.I(net270),
    .Z(data_out_real[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output224 (.I(net271),
    .Z(data_out_real[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output225 (.I(net272),
    .Z(data_out_real[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output226 (.I(net273),
    .Z(data_out_real[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output227 (.I(net274),
    .Z(data_out_real[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output228 (.I(net275),
    .Z(data_out_real[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output229 (.I(net276),
    .Z(data_out_real[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output230 (.I(net277),
    .Z(data_out_real[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output231 (.I(net278),
    .Z(data_out_real[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output232 (.I(net279),
    .Z(data_out_real[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output233 (.I(net280),
    .Z(data_out_real[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output234 (.I(net281),
    .Z(data_out_real[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output235 (.I(net282),
    .Z(data_out_real[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output236 (.I(net283),
    .Z(data_out_real[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output237 (.I(net284),
    .Z(data_out_real[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output238 (.I(net285),
    .Z(data_out_real[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output239 (.I(net286),
    .Z(data_out_real[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output240 (.I(net287),
    .Z(data_out_real[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output241 (.I(net288),
    .Z(data_out_real[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output242 (.I(net289),
    .Z(data_out_real[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output243 (.I(net290),
    .Z(data_out_real[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output244 (.I(net291),
    .Z(data_out_real[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output245 (.I(net292),
    .Z(data_out_real[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output246 (.I(net293),
    .Z(data_out_real[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output247 (.I(net294),
    .Z(data_out_real[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output248 (.I(net295),
    .Z(data_out_real[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output249 (.I(net296),
    .Z(data_out_real[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output250 (.I(net297),
    .Z(data_out_real[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output251 (.I(net298),
    .Z(data_out_real[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output252 (.I(net299),
    .Z(data_out_real[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output253 (.I(net300),
    .Z(data_out_real[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output254 (.I(net301),
    .Z(data_out_real[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output255 (.I(net302),
    .Z(data_out_real[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output256 (.I(net303),
    .Z(data_out_real[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output257 (.I(net304),
    .Z(data_out_real[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output258 (.I(net305),
    .Z(data_out_real[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output259 (.I(net306),
    .Z(data_out_real[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output260 (.I(net307),
    .Z(data_out_real[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output261 (.I(net308),
    .Z(data_out_real[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output262 (.I(net309),
    .Z(data_out_real[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output263 (.I(net310),
    .Z(data_out_real[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output264 (.I(net311),
    .Z(data_out_real[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output265 (.I(net312),
    .Z(data_out_real[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output266 (.I(net313),
    .Z(data_out_real[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output267 (.I(net314),
    .Z(data_out_real[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output268 (.I(net315),
    .Z(data_out_real[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output269 (.I(net316),
    .Z(data_out_real[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output270 (.I(net317),
    .Z(data_out_real[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output271 (.I(net318),
    .Z(data_out_real[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output272 (.I(net319),
    .Z(data_out_real[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output273 (.I(net320),
    .Z(data_out_real[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output274 (.I(net321),
    .Z(data_out_real[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output275 (.I(net322),
    .Z(data_out_real[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output276 (.I(net323),
    .Z(data_out_real[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output277 (.I(net324),
    .Z(data_out_real[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output278 (.I(net325),
    .Z(data_out_real[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output279 (.I(net326),
    .Z(data_out_real[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output280 (.I(net327),
    .Z(data_out_real[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output281 (.I(net328),
    .Z(data_out_real[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output282 (.I(net329),
    .Z(data_out_real[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output283 (.I(net330),
    .Z(data_out_real[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output284 (.I(net331),
    .Z(data_out_real[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output285 (.I(net332),
    .Z(data_out_real[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output286 (.I(net333),
    .Z(data_out_real[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output287 (.I(net334),
    .Z(data_out_real[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output288 (.I(net335),
    .Z(data_out_real[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output289 (.I(net336),
    .Z(data_out_real[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output290 (.I(net337),
    .Z(data_out_real[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output291 (.I(net338),
    .Z(data_out_real[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output292 (.I(net339),
    .Z(data_out_real[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output293 (.I(net340),
    .Z(data_ready));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output294 (.I(net341),
    .Z(data_valid_out));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15241__295 (.ZN(net342));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15245__296 (.ZN(net343));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15250__297 (.ZN(net344));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15252__298 (.ZN(net345));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15263__299 (.ZN(net346));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15270__300 (.ZN(net347));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15278__301 (.ZN(net348));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15285__302 (.ZN(net349));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15291__303 (.ZN(net350));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15299__304 (.ZN(net351));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15304__305 (.ZN(net352));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15313__306 (.ZN(net353));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15320__307 (.ZN(net354));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15327__308 (.ZN(net355));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15328__309 (.ZN(net356));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15336__310 (.ZN(net357));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15344__311 (.ZN(net358));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15352__312 (.ZN(net359));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15360__313 (.ZN(net360));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15368__314 (.ZN(net361));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15376__315 (.ZN(net362));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15383__316 (.ZN(net363));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15384__317 (.ZN(net364));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15392__318 (.ZN(net365));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15399__319 (.ZN(net366));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15410__320 (.ZN(net367));
 gf180mcu_fd_sc_mcu9t5v0__tiel _15415__321 (.ZN(net368));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload1 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload2 (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload3 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload4 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload5 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload6 (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload7 (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload8 (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload9 (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload10 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload11 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload12 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload13 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload14 (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload15 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload16 (.I(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload17 (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload18 (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload19 (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload20 (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer1 (.I(_03430_),
    .Z(net370));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer2 (.I(_03430_),
    .Z(net371));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer3 (.I(net371),
    .Z(net372));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer4 (.I(_03106_),
    .Z(net373));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer5 (.I(_03294_),
    .Z(net374));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer6 (.I(_03294_),
    .Z(net375));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer7 (.I(_03294_),
    .Z(net376));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer8 (.I(_03230_),
    .Z(net377));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer9 (.I(_03108_),
    .Z(net378));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer10 (.I(_07627_),
    .Z(net379));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer11 (.I(_03004_),
    .Z(net380));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer12 (.I(_03229_),
    .Z(net381));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer13 (.I(_07629_),
    .Z(net382));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer14 (.I(net394),
    .Z(net383));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 clone21 (.A1(_02752_),
    .A2(_02842_),
    .Z(net384));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer23 (.I(_03212_),
    .Z(net386));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer24 (.I(_03126_),
    .Z(net387));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer25 (.I(_03305_),
    .Z(net388));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer26 (.I(_03124_),
    .Z(net389));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer27 (.I(net392),
    .Z(net390));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer31 (.I(net395),
    .Z(net394));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer32 (.I(net396),
    .Z(net395));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer33 (.I(_03231_),
    .Z(net396));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer15 (.I(_03004_),
    .Z(net385));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer16 (.I(_07629_),
    .Z(net391));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer17 (.I(net393),
    .Z(net392));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer18 (.I(net397),
    .Z(net393));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer19 (.I(net398),
    .Z(net397));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer20 (.I(net399),
    .Z(net398));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer21 (.I(net400),
    .Z(net399));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 rebuffer22 (.I(_03293_),
    .Z(net400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer28 (.I(_03295_),
    .Z(net401));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net100));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net208));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1732 ();
endmodule
