module async_fifo (almost_empty,
    almost_full,
    empty,
    full,
    pointer_wraparound_flag,
    rd_clk,
    rd_en,
    rd_rst_n,
    sync_error_flag,
    wr_clk,
    wr_en,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output almost_empty;
 output almost_full;
 output empty;
 output full;
 output pointer_wraparound_flag;
 input rd_clk;
 input rd_en;
 input rd_rst_n;
 output sync_error_flag;
 input wr_clk;
 input wr_en;
 input wr_rst_n;
 output [4:0] rd_count;
 output [7:0] rd_data;
 output [4:0] wr_count;
 input [7:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \rd_ptr_sync[0] ;
 wire \rd_ptr_sync[1] ;
 wire \rd_ptr_sync[2] ;
 wire \rd_ptr_sync[3] ;
 wire \rd_ptr_sync[4] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire \wr_ptr_sync[0] ;
 wire \wr_ptr_sync[1] ;
 wire \wr_ptr_sync[2] ;
 wire \wr_ptr_sync[3] ;
 wire \wr_ptr_sync[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;

 INV_X1 _0648_ (.A(_0616_),
    .ZN(net12));
 INV_X1 _0649_ (.A(_0609_),
    .ZN(_0169_));
 BUF_X1 _0650_ (.A(_0613_),
    .Z(_0170_));
 NAND4_X1 _0651_ (.A1(_0603_),
    .A2(_0170_),
    .A3(_0616_),
    .A4(_0607_),
    .ZN(_0171_));
 NOR2_X1 _0652_ (.A1(_0169_),
    .A2(_0171_),
    .ZN(_0000_));
 AOI21_X1 _0653_ (.A(_0612_),
    .B1(_0597_),
    .B2(_0170_),
    .ZN(_0172_));
 INV_X1 _0654_ (.A(_0172_),
    .ZN(_0173_));
 AOI21_X1 _0655_ (.A(_0602_),
    .B1(_0173_),
    .B2(_0603_),
    .ZN(_0174_));
 XNOR2_X1 _0656_ (.A(_0607_),
    .B(_0174_),
    .ZN(net16));
 XOR2_X1 _0657_ (.A(_0170_),
    .B(_0597_),
    .Z(net14));
 INV_X1 _0658_ (.A(_0608_),
    .ZN(_0175_));
 OAI21_X1 _0659_ (.A(_0175_),
    .B1(_0169_),
    .B2(_0618_),
    .ZN(_0176_));
 AOI21_X1 _0660_ (.A(_0612_),
    .B1(_0176_),
    .B2(_0170_),
    .ZN(_0177_));
 XNOR2_X1 _0661_ (.A(_0603_),
    .B(_0177_),
    .ZN(net15));
 INV_X1 _0662_ (.A(_0623_),
    .ZN(net26));
 INV_X1 _0663_ (.A(_0634_),
    .ZN(_0178_));
 INV_X1 _0664_ (.A(_0626_),
    .ZN(_0179_));
 INV_X1 _0665_ (.A(_0620_),
    .ZN(_0180_));
 OAI21_X1 _0666_ (.A(_0179_),
    .B1(_0624_),
    .B2(_0180_),
    .ZN(_0181_));
 BUF_X1 _0667_ (.A(_0630_),
    .Z(_0182_));
 AOI21_X1 _0668_ (.A(_0629_),
    .B1(_0181_),
    .B2(_0182_),
    .ZN(_0183_));
 XNOR2_X1 _0669_ (.A(_0178_),
    .B(_0183_),
    .ZN(_0184_));
 INV_X1 _0670_ (.A(_0184_),
    .ZN(net29));
 INV_X1 _0671_ (.A(_0633_),
    .ZN(_0185_));
 AOI21_X1 _0672_ (.A(_0629_),
    .B1(_0600_),
    .B2(_0182_),
    .ZN(_0186_));
 OAI21_X1 _0673_ (.A(_0185_),
    .B1(_0186_),
    .B2(_0178_),
    .ZN(_0187_));
 XNOR2_X1 _0674_ (.A(_0638_),
    .B(_0187_),
    .ZN(_0188_));
 INV_X1 _0675_ (.A(_0188_),
    .ZN(net30));
 NOR4_X1 _0676_ (.A1(\rd_ptr_sync[1] ),
    .A2(\rd_ptr_sync[0] ),
    .A3(\rd_ptr_sync[3] ),
    .A4(\rd_ptr_sync[2] ),
    .ZN(_0189_));
 CLKBUF_X3 _0677_ (.A(_0640_),
    .Z(_0190_));
 CLKBUF_X3 _0678_ (.A(\wr_ptr_bin[3] ),
    .Z(_0191_));
 BUF_X4 _0679_ (.A(\wr_ptr_bin[2] ),
    .Z(_0192_));
 NOR2_X4 _0680_ (.A1(_0191_),
    .A2(_0192_),
    .ZN(_0193_));
 NAND3_X1 _0681_ (.A1(\wr_ptr_bin[4] ),
    .A2(_0190_),
    .A3(_0193_),
    .ZN(_0194_));
 NOR2_X1 _0682_ (.A1(_0189_),
    .A2(_0194_),
    .ZN(_0010_));
 NAND3_X1 _0683_ (.A1(_0620_),
    .A2(_0634_),
    .A3(_0182_),
    .ZN(_0195_));
 NOR3_X1 _0684_ (.A1(net26),
    .A2(_0638_),
    .A3(_0195_),
    .ZN(_0001_));
 XOR2_X2 _0685_ (.A(\wr_ptr_gray_sync2[4] ),
    .B(\wr_ptr_gray_sync2[3] ),
    .Z(_0005_));
 XOR2_X2 _0686_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(_0005_),
    .Z(_0004_));
 XOR2_X2 _0687_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(_0004_),
    .Z(_0003_));
 XOR2_X1 _0688_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(_0003_),
    .Z(_0002_));
 XOR2_X2 _0689_ (.A(\rd_ptr_gray_sync2[4] ),
    .B(\rd_ptr_gray_sync2[3] ),
    .Z(_0009_));
 XOR2_X2 _0690_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(_0009_),
    .Z(_0008_));
 XOR2_X2 _0691_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(_0008_),
    .Z(_0007_));
 XOR2_X1 _0692_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(_0007_),
    .Z(_0006_));
 INV_X1 _0693_ (.A(_0618_),
    .ZN(_0596_));
 INV_X1 _0694_ (.A(_0624_),
    .ZN(_0599_));
 BUF_X1 _0695_ (.A(wr_data[0]),
    .Z(_0196_));
 BUF_X2 _0696_ (.A(_0196_),
    .Z(_0197_));
 INV_X1 _0697_ (.A(net5),
    .ZN(_0198_));
 NOR2_X1 _0698_ (.A1(_0198_),
    .A2(net10),
    .ZN(_0199_));
 BUF_X8 _0699_ (.A(_0199_),
    .Z(_0200_));
 NAND3_X4 _0700_ (.A1(_0190_),
    .A2(_0193_),
    .A3(_0200_),
    .ZN(_0201_));
 MUX2_X1 _0701_ (.A(_0197_),
    .B(\mem[0][0] ),
    .S(_0201_),
    .Z(_0015_));
 CLKBUF_X2 _0702_ (.A(wr_data[1]),
    .Z(_0202_));
 BUF_X2 _0703_ (.A(_0202_),
    .Z(_0203_));
 MUX2_X1 _0704_ (.A(_0203_),
    .B(\mem[0][1] ),
    .S(_0201_),
    .Z(_0016_));
 CLKBUF_X2 _0705_ (.A(wr_data[2]),
    .Z(_0204_));
 BUF_X2 _0706_ (.A(_0204_),
    .Z(_0205_));
 MUX2_X1 _0707_ (.A(_0205_),
    .B(\mem[0][2] ),
    .S(_0201_),
    .Z(_0017_));
 CLKBUF_X2 _0708_ (.A(wr_data[3]),
    .Z(_0206_));
 BUF_X2 _0709_ (.A(_0206_),
    .Z(_0207_));
 MUX2_X1 _0710_ (.A(_0207_),
    .B(\mem[0][3] ),
    .S(_0201_),
    .Z(_0018_));
 BUF_X1 _0711_ (.A(wr_data[4]),
    .Z(_0208_));
 BUF_X2 _0712_ (.A(_0208_),
    .Z(_0209_));
 MUX2_X1 _0713_ (.A(_0209_),
    .B(\mem[0][4] ),
    .S(_0201_),
    .Z(_0019_));
 CLKBUF_X2 _0714_ (.A(wr_data[5]),
    .Z(_0210_));
 BUF_X2 _0715_ (.A(_0210_),
    .Z(_0211_));
 MUX2_X1 _0716_ (.A(_0211_),
    .B(\mem[0][5] ),
    .S(_0201_),
    .Z(_0020_));
 CLKBUF_X2 _0717_ (.A(wr_data[6]),
    .Z(_0212_));
 BUF_X2 _0718_ (.A(_0212_),
    .Z(_0213_));
 MUX2_X1 _0719_ (.A(_0213_),
    .B(\mem[0][6] ),
    .S(_0201_),
    .Z(_0021_));
 CLKBUF_X2 _0720_ (.A(wr_data[7]),
    .Z(_0214_));
 BUF_X2 _0721_ (.A(_0214_),
    .Z(_0215_));
 MUX2_X1 _0722_ (.A(_0215_),
    .B(\mem[0][7] ),
    .S(_0201_),
    .Z(_0022_));
 INV_X2 _0723_ (.A(_0192_),
    .ZN(_0216_));
 NAND2_X4 _0724_ (.A1(_0191_),
    .A2(_0216_),
    .ZN(_0217_));
 BUF_X2 _0725_ (.A(_0641_),
    .Z(_0218_));
 NAND2_X2 _0726_ (.A1(_0218_),
    .A2(_0200_),
    .ZN(_0219_));
 NOR2_X4 _0727_ (.A1(_0217_),
    .A2(_0219_),
    .ZN(_0220_));
 MUX2_X1 _0728_ (.A(\mem[10][0] ),
    .B(_0197_),
    .S(_0220_),
    .Z(_0023_));
 MUX2_X1 _0729_ (.A(\mem[10][1] ),
    .B(_0203_),
    .S(_0220_),
    .Z(_0024_));
 MUX2_X1 _0730_ (.A(\mem[10][2] ),
    .B(_0205_),
    .S(_0220_),
    .Z(_0025_));
 MUX2_X1 _0731_ (.A(\mem[10][3] ),
    .B(_0207_),
    .S(_0220_),
    .Z(_0026_));
 MUX2_X1 _0732_ (.A(\mem[10][4] ),
    .B(_0209_),
    .S(_0220_),
    .Z(_0027_));
 MUX2_X1 _0733_ (.A(\mem[10][5] ),
    .B(_0211_),
    .S(_0220_),
    .Z(_0028_));
 MUX2_X1 _0734_ (.A(\mem[10][6] ),
    .B(_0213_),
    .S(_0220_),
    .Z(_0029_));
 MUX2_X1 _0735_ (.A(\mem[10][7] ),
    .B(_0215_),
    .S(_0220_),
    .Z(_0030_));
 BUF_X4 _0736_ (.A(_0645_),
    .Z(_0221_));
 NAND2_X4 _0737_ (.A1(_0221_),
    .A2(_0200_),
    .ZN(_0222_));
 NOR2_X4 _0738_ (.A1(_0217_),
    .A2(_0222_),
    .ZN(_0223_));
 MUX2_X1 _0739_ (.A(\mem[11][0] ),
    .B(_0197_),
    .S(_0223_),
    .Z(_0031_));
 MUX2_X1 _0740_ (.A(\mem[11][1] ),
    .B(_0203_),
    .S(_0223_),
    .Z(_0032_));
 MUX2_X1 _0741_ (.A(\mem[11][2] ),
    .B(_0205_),
    .S(_0223_),
    .Z(_0033_));
 MUX2_X1 _0742_ (.A(\mem[11][3] ),
    .B(_0207_),
    .S(_0223_),
    .Z(_0034_));
 MUX2_X1 _0743_ (.A(\mem[11][4] ),
    .B(_0209_),
    .S(_0223_),
    .Z(_0035_));
 MUX2_X1 _0744_ (.A(\mem[11][5] ),
    .B(_0211_),
    .S(_0223_),
    .Z(_0036_));
 MUX2_X1 _0745_ (.A(\mem[11][6] ),
    .B(_0213_),
    .S(_0223_),
    .Z(_0037_));
 MUX2_X1 _0746_ (.A(\mem[11][7] ),
    .B(_0215_),
    .S(_0223_),
    .Z(_0038_));
 BUF_X4 _0747_ (.A(_0200_),
    .Z(_0224_));
 INV_X2 _0748_ (.A(_0191_),
    .ZN(_0225_));
 NOR2_X4 _0749_ (.A1(_0225_),
    .A2(_0216_),
    .ZN(_0226_));
 NAND3_X4 _0750_ (.A1(_0190_),
    .A2(_0224_),
    .A3(_0226_),
    .ZN(_0227_));
 MUX2_X1 _0751_ (.A(_0197_),
    .B(\mem[12][0] ),
    .S(_0227_),
    .Z(_0039_));
 MUX2_X1 _0752_ (.A(_0203_),
    .B(\mem[12][1] ),
    .S(_0227_),
    .Z(_0040_));
 MUX2_X1 _0753_ (.A(_0205_),
    .B(\mem[12][2] ),
    .S(_0227_),
    .Z(_0041_));
 MUX2_X1 _0754_ (.A(_0207_),
    .B(\mem[12][3] ),
    .S(_0227_),
    .Z(_0042_));
 MUX2_X1 _0755_ (.A(_0209_),
    .B(\mem[12][4] ),
    .S(_0227_),
    .Z(_0043_));
 MUX2_X1 _0756_ (.A(_0211_),
    .B(\mem[12][5] ),
    .S(_0227_),
    .Z(_0044_));
 MUX2_X1 _0757_ (.A(_0213_),
    .B(\mem[12][6] ),
    .S(_0227_),
    .Z(_0045_));
 MUX2_X1 _0758_ (.A(_0215_),
    .B(\mem[12][7] ),
    .S(_0227_),
    .Z(_0046_));
 BUF_X2 _0759_ (.A(_0643_),
    .Z(_0228_));
 NAND3_X4 _0760_ (.A1(_0228_),
    .A2(_0224_),
    .A3(_0226_),
    .ZN(_0229_));
 MUX2_X1 _0761_ (.A(_0196_),
    .B(\mem[13][0] ),
    .S(_0229_),
    .Z(_0047_));
 MUX2_X1 _0762_ (.A(_0202_),
    .B(\mem[13][1] ),
    .S(_0229_),
    .Z(_0048_));
 MUX2_X1 _0763_ (.A(_0204_),
    .B(\mem[13][2] ),
    .S(_0229_),
    .Z(_0049_));
 MUX2_X1 _0764_ (.A(_0206_),
    .B(\mem[13][3] ),
    .S(_0229_),
    .Z(_0050_));
 MUX2_X1 _0765_ (.A(_0208_),
    .B(\mem[13][4] ),
    .S(_0229_),
    .Z(_0051_));
 MUX2_X1 _0766_ (.A(_0210_),
    .B(\mem[13][5] ),
    .S(_0229_),
    .Z(_0052_));
 MUX2_X1 _0767_ (.A(_0212_),
    .B(\mem[13][6] ),
    .S(_0229_),
    .Z(_0053_));
 MUX2_X1 _0768_ (.A(_0214_),
    .B(\mem[13][7] ),
    .S(_0229_),
    .Z(_0054_));
 NAND3_X4 _0769_ (.A1(_0218_),
    .A2(_0224_),
    .A3(_0226_),
    .ZN(_0230_));
 MUX2_X1 _0770_ (.A(_0196_),
    .B(\mem[14][0] ),
    .S(_0230_),
    .Z(_0055_));
 MUX2_X1 _0771_ (.A(_0202_),
    .B(\mem[14][1] ),
    .S(_0230_),
    .Z(_0056_));
 MUX2_X1 _0772_ (.A(_0204_),
    .B(\mem[14][2] ),
    .S(_0230_),
    .Z(_0057_));
 MUX2_X1 _0773_ (.A(_0206_),
    .B(\mem[14][3] ),
    .S(_0230_),
    .Z(_0058_));
 MUX2_X1 _0774_ (.A(_0208_),
    .B(\mem[14][4] ),
    .S(_0230_),
    .Z(_0059_));
 MUX2_X1 _0775_ (.A(_0210_),
    .B(\mem[14][5] ),
    .S(_0230_),
    .Z(_0060_));
 MUX2_X1 _0776_ (.A(_0212_),
    .B(\mem[14][6] ),
    .S(_0230_),
    .Z(_0061_));
 MUX2_X1 _0777_ (.A(_0214_),
    .B(\mem[14][7] ),
    .S(_0230_),
    .Z(_0062_));
 NAND3_X4 _0778_ (.A1(_0221_),
    .A2(_0200_),
    .A3(_0226_),
    .ZN(_0231_));
 MUX2_X1 _0779_ (.A(_0196_),
    .B(\mem[15][0] ),
    .S(_0231_),
    .Z(_0063_));
 MUX2_X1 _0780_ (.A(_0202_),
    .B(\mem[15][1] ),
    .S(_0231_),
    .Z(_0064_));
 MUX2_X1 _0781_ (.A(_0204_),
    .B(\mem[15][2] ),
    .S(_0231_),
    .Z(_0065_));
 MUX2_X1 _0782_ (.A(_0206_),
    .B(\mem[15][3] ),
    .S(_0231_),
    .Z(_0066_));
 MUX2_X1 _0783_ (.A(_0208_),
    .B(\mem[15][4] ),
    .S(_0231_),
    .Z(_0067_));
 MUX2_X1 _0784_ (.A(_0210_),
    .B(\mem[15][5] ),
    .S(_0231_),
    .Z(_0068_));
 MUX2_X1 _0785_ (.A(_0212_),
    .B(\mem[15][6] ),
    .S(_0231_),
    .Z(_0069_));
 MUX2_X1 _0786_ (.A(_0214_),
    .B(\mem[15][7] ),
    .S(_0231_),
    .Z(_0070_));
 NAND3_X4 _0787_ (.A1(_0228_),
    .A2(_0193_),
    .A3(_0200_),
    .ZN(_0232_));
 MUX2_X1 _0788_ (.A(_0196_),
    .B(\mem[1][0] ),
    .S(_0232_),
    .Z(_0071_));
 MUX2_X1 _0789_ (.A(_0202_),
    .B(\mem[1][1] ),
    .S(_0232_),
    .Z(_0072_));
 MUX2_X1 _0790_ (.A(_0204_),
    .B(\mem[1][2] ),
    .S(_0232_),
    .Z(_0073_));
 MUX2_X1 _0791_ (.A(_0206_),
    .B(\mem[1][3] ),
    .S(_0232_),
    .Z(_0074_));
 MUX2_X1 _0792_ (.A(_0208_),
    .B(\mem[1][4] ),
    .S(_0232_),
    .Z(_0075_));
 MUX2_X1 _0793_ (.A(_0210_),
    .B(\mem[1][5] ),
    .S(_0232_),
    .Z(_0076_));
 MUX2_X1 _0794_ (.A(_0212_),
    .B(\mem[1][6] ),
    .S(_0232_),
    .Z(_0077_));
 MUX2_X1 _0795_ (.A(_0214_),
    .B(\mem[1][7] ),
    .S(_0232_),
    .Z(_0078_));
 NAND3_X4 _0796_ (.A1(_0218_),
    .A2(_0193_),
    .A3(_0200_),
    .ZN(_0233_));
 MUX2_X1 _0797_ (.A(_0196_),
    .B(\mem[2][0] ),
    .S(_0233_),
    .Z(_0079_));
 MUX2_X1 _0798_ (.A(_0202_),
    .B(\mem[2][1] ),
    .S(_0233_),
    .Z(_0080_));
 MUX2_X1 _0799_ (.A(_0204_),
    .B(\mem[2][2] ),
    .S(_0233_),
    .Z(_0081_));
 MUX2_X1 _0800_ (.A(_0206_),
    .B(\mem[2][3] ),
    .S(_0233_),
    .Z(_0082_));
 MUX2_X1 _0801_ (.A(_0208_),
    .B(\mem[2][4] ),
    .S(_0233_),
    .Z(_0083_));
 MUX2_X1 _0802_ (.A(_0210_),
    .B(\mem[2][5] ),
    .S(_0233_),
    .Z(_0084_));
 MUX2_X1 _0803_ (.A(_0212_),
    .B(\mem[2][6] ),
    .S(_0233_),
    .Z(_0085_));
 MUX2_X1 _0804_ (.A(_0214_),
    .B(\mem[2][7] ),
    .S(_0233_),
    .Z(_0086_));
 NAND3_X4 _0805_ (.A1(_0221_),
    .A2(_0193_),
    .A3(_0200_),
    .ZN(_0234_));
 MUX2_X1 _0806_ (.A(_0196_),
    .B(\mem[3][0] ),
    .S(_0234_),
    .Z(_0087_));
 MUX2_X1 _0807_ (.A(_0202_),
    .B(\mem[3][1] ),
    .S(_0234_),
    .Z(_0088_));
 MUX2_X1 _0808_ (.A(_0204_),
    .B(\mem[3][2] ),
    .S(_0234_),
    .Z(_0089_));
 MUX2_X1 _0809_ (.A(_0206_),
    .B(\mem[3][3] ),
    .S(_0234_),
    .Z(_0090_));
 MUX2_X1 _0810_ (.A(_0208_),
    .B(\mem[3][4] ),
    .S(_0234_),
    .Z(_0091_));
 MUX2_X1 _0811_ (.A(_0210_),
    .B(\mem[3][5] ),
    .S(_0234_),
    .Z(_0092_));
 MUX2_X1 _0812_ (.A(_0212_),
    .B(\mem[3][6] ),
    .S(_0234_),
    .Z(_0093_));
 MUX2_X1 _0813_ (.A(_0214_),
    .B(\mem[3][7] ),
    .S(_0234_),
    .Z(_0094_));
 NAND2_X2 _0814_ (.A1(_0190_),
    .A2(_0200_),
    .ZN(_0235_));
 NAND2_X4 _0815_ (.A1(_0225_),
    .A2(_0192_),
    .ZN(_0236_));
 NOR2_X4 _0816_ (.A1(_0235_),
    .A2(_0236_),
    .ZN(_0237_));
 MUX2_X1 _0817_ (.A(\mem[4][0] ),
    .B(_0197_),
    .S(_0237_),
    .Z(_0095_));
 MUX2_X1 _0818_ (.A(\mem[4][1] ),
    .B(_0203_),
    .S(_0237_),
    .Z(_0096_));
 MUX2_X1 _0819_ (.A(\mem[4][2] ),
    .B(_0205_),
    .S(_0237_),
    .Z(_0097_));
 MUX2_X1 _0820_ (.A(\mem[4][3] ),
    .B(_0207_),
    .S(_0237_),
    .Z(_0098_));
 MUX2_X1 _0821_ (.A(\mem[4][4] ),
    .B(_0209_),
    .S(_0237_),
    .Z(_0099_));
 MUX2_X1 _0822_ (.A(\mem[4][5] ),
    .B(_0211_),
    .S(_0237_),
    .Z(_0100_));
 MUX2_X1 _0823_ (.A(\mem[4][6] ),
    .B(_0213_),
    .S(_0237_),
    .Z(_0101_));
 MUX2_X1 _0824_ (.A(\mem[4][7] ),
    .B(_0215_),
    .S(_0237_),
    .Z(_0102_));
 NAND2_X2 _0825_ (.A1(_0228_),
    .A2(_0200_),
    .ZN(_0238_));
 NOR2_X4 _0826_ (.A1(_0238_),
    .A2(_0236_),
    .ZN(_0239_));
 MUX2_X1 _0827_ (.A(\mem[5][0] ),
    .B(_0197_),
    .S(_0239_),
    .Z(_0103_));
 MUX2_X1 _0828_ (.A(\mem[5][1] ),
    .B(_0203_),
    .S(_0239_),
    .Z(_0104_));
 MUX2_X1 _0829_ (.A(\mem[5][2] ),
    .B(_0205_),
    .S(_0239_),
    .Z(_0105_));
 MUX2_X1 _0830_ (.A(\mem[5][3] ),
    .B(_0207_),
    .S(_0239_),
    .Z(_0106_));
 MUX2_X1 _0831_ (.A(\mem[5][4] ),
    .B(_0209_),
    .S(_0239_),
    .Z(_0107_));
 MUX2_X1 _0832_ (.A(\mem[5][5] ),
    .B(_0211_),
    .S(_0239_),
    .Z(_0108_));
 MUX2_X1 _0833_ (.A(\mem[5][6] ),
    .B(_0213_),
    .S(_0239_),
    .Z(_0109_));
 MUX2_X1 _0834_ (.A(\mem[5][7] ),
    .B(_0215_),
    .S(_0239_),
    .Z(_0110_));
 NOR2_X4 _0835_ (.A1(_0219_),
    .A2(_0236_),
    .ZN(_0240_));
 MUX2_X1 _0836_ (.A(\mem[6][0] ),
    .B(_0197_),
    .S(_0240_),
    .Z(_0111_));
 MUX2_X1 _0837_ (.A(\mem[6][1] ),
    .B(_0203_),
    .S(_0240_),
    .Z(_0112_));
 MUX2_X1 _0838_ (.A(\mem[6][2] ),
    .B(_0205_),
    .S(_0240_),
    .Z(_0113_));
 MUX2_X1 _0839_ (.A(\mem[6][3] ),
    .B(_0207_),
    .S(_0240_),
    .Z(_0114_));
 MUX2_X1 _0840_ (.A(\mem[6][4] ),
    .B(_0209_),
    .S(_0240_),
    .Z(_0115_));
 MUX2_X1 _0841_ (.A(\mem[6][5] ),
    .B(_0211_),
    .S(_0240_),
    .Z(_0116_));
 MUX2_X1 _0842_ (.A(\mem[6][6] ),
    .B(_0213_),
    .S(_0240_),
    .Z(_0117_));
 MUX2_X1 _0843_ (.A(\mem[6][7] ),
    .B(_0215_),
    .S(_0240_),
    .Z(_0118_));
 NOR2_X4 _0844_ (.A1(_0222_),
    .A2(_0236_),
    .ZN(_0241_));
 MUX2_X1 _0845_ (.A(\mem[7][0] ),
    .B(_0197_),
    .S(_0241_),
    .Z(_0119_));
 MUX2_X1 _0846_ (.A(\mem[7][1] ),
    .B(_0203_),
    .S(_0241_),
    .Z(_0120_));
 MUX2_X1 _0847_ (.A(\mem[7][2] ),
    .B(_0205_),
    .S(_0241_),
    .Z(_0121_));
 MUX2_X1 _0848_ (.A(\mem[7][3] ),
    .B(_0207_),
    .S(_0241_),
    .Z(_0122_));
 MUX2_X1 _0849_ (.A(\mem[7][4] ),
    .B(_0209_),
    .S(_0241_),
    .Z(_0123_));
 MUX2_X1 _0850_ (.A(\mem[7][5] ),
    .B(_0211_),
    .S(_0241_),
    .Z(_0124_));
 MUX2_X1 _0851_ (.A(\mem[7][6] ),
    .B(_0213_),
    .S(_0241_),
    .Z(_0125_));
 MUX2_X1 _0852_ (.A(\mem[7][7] ),
    .B(_0215_),
    .S(_0241_),
    .Z(_0126_));
 NOR2_X4 _0853_ (.A1(_0235_),
    .A2(_0217_),
    .ZN(_0242_));
 MUX2_X1 _0854_ (.A(\mem[8][0] ),
    .B(_0197_),
    .S(_0242_),
    .Z(_0127_));
 MUX2_X1 _0855_ (.A(\mem[8][1] ),
    .B(_0203_),
    .S(_0242_),
    .Z(_0128_));
 MUX2_X1 _0856_ (.A(\mem[8][2] ),
    .B(_0205_),
    .S(_0242_),
    .Z(_0129_));
 MUX2_X1 _0857_ (.A(\mem[8][3] ),
    .B(_0207_),
    .S(_0242_),
    .Z(_0130_));
 MUX2_X1 _0858_ (.A(\mem[8][4] ),
    .B(_0209_),
    .S(_0242_),
    .Z(_0131_));
 MUX2_X1 _0859_ (.A(\mem[8][5] ),
    .B(_0211_),
    .S(_0242_),
    .Z(_0132_));
 MUX2_X1 _0860_ (.A(\mem[8][6] ),
    .B(_0213_),
    .S(_0242_),
    .Z(_0133_));
 MUX2_X1 _0861_ (.A(\mem[8][7] ),
    .B(_0215_),
    .S(_0242_),
    .Z(_0134_));
 NOR2_X4 _0862_ (.A1(_0217_),
    .A2(_0238_),
    .ZN(_0243_));
 MUX2_X1 _0863_ (.A(\mem[9][0] ),
    .B(_0197_),
    .S(_0243_),
    .Z(_0135_));
 MUX2_X1 _0864_ (.A(\mem[9][1] ),
    .B(_0203_),
    .S(_0243_),
    .Z(_0136_));
 MUX2_X1 _0865_ (.A(\mem[9][2] ),
    .B(_0205_),
    .S(_0243_),
    .Z(_0137_));
 MUX2_X1 _0866_ (.A(\mem[9][3] ),
    .B(_0207_),
    .S(_0243_),
    .Z(_0138_));
 MUX2_X1 _0867_ (.A(\mem[9][4] ),
    .B(_0209_),
    .S(_0243_),
    .Z(_0139_));
 MUX2_X1 _0868_ (.A(\mem[9][5] ),
    .B(_0211_),
    .S(_0243_),
    .Z(_0140_));
 MUX2_X1 _0869_ (.A(\mem[9][6] ),
    .B(_0213_),
    .S(_0243_),
    .Z(_0141_));
 MUX2_X1 _0870_ (.A(\mem[9][7] ),
    .B(_0215_),
    .S(_0243_),
    .Z(_0142_));
 BUF_X4 _0871_ (.A(\rd_ptr_bin[2] ),
    .Z(_0244_));
 MUX2_X1 _0872_ (.A(\mem[1][0] ),
    .B(\mem[5][0] ),
    .S(_0244_),
    .Z(_0245_));
 MUX2_X1 _0873_ (.A(\mem[3][0] ),
    .B(\mem[7][0] ),
    .S(_0244_),
    .Z(_0246_));
 BUF_X2 _0874_ (.A(\rd_ptr_bin[1] ),
    .Z(_0247_));
 CLKBUF_X3 _0875_ (.A(_0247_),
    .Z(_0248_));
 MUX2_X1 _0876_ (.A(_0245_),
    .B(_0246_),
    .S(_0248_),
    .Z(_0249_));
 MUX2_X1 _0877_ (.A(\mem[0][0] ),
    .B(\mem[4][0] ),
    .S(_0244_),
    .Z(_0250_));
 BUF_X8 _0878_ (.A(_0244_),
    .Z(_0251_));
 MUX2_X1 _0879_ (.A(\mem[2][0] ),
    .B(\mem[6][0] ),
    .S(_0251_),
    .Z(_0252_));
 MUX2_X1 _0880_ (.A(_0250_),
    .B(_0252_),
    .S(_0248_),
    .Z(_0253_));
 BUF_X2 _0881_ (.A(\rd_ptr_bin[0] ),
    .Z(_0254_));
 BUF_X4 _0882_ (.A(_0254_),
    .Z(_0255_));
 INV_X1 _0883_ (.A(_0255_),
    .ZN(_0256_));
 MUX2_X1 _0884_ (.A(_0249_),
    .B(_0253_),
    .S(_0256_),
    .Z(_0257_));
 CLKBUF_X3 _0885_ (.A(_0255_),
    .Z(_0258_));
 CLKBUF_X3 _0886_ (.A(_0251_),
    .Z(_0259_));
 INV_X1 _0887_ (.A(_0259_),
    .ZN(_0260_));
 MUX2_X1 _0888_ (.A(\mem[12][0] ),
    .B(\mem[14][0] ),
    .S(_0247_),
    .Z(_0261_));
 NOR3_X1 _0889_ (.A1(_0258_),
    .A2(_0260_),
    .A3(_0261_),
    .ZN(_0262_));
 MUX2_X1 _0890_ (.A(\mem[9][0] ),
    .B(\mem[11][0] ),
    .S(_0247_),
    .Z(_0263_));
 NOR3_X1 _0891_ (.A1(_0256_),
    .A2(_0259_),
    .A3(_0263_),
    .ZN(_0264_));
 MUX2_X1 _0892_ (.A(\mem[8][0] ),
    .B(\mem[10][0] ),
    .S(_0247_),
    .Z(_0265_));
 NOR3_X1 _0893_ (.A1(_0255_),
    .A2(_0259_),
    .A3(_0265_),
    .ZN(_0266_));
 MUX2_X1 _0894_ (.A(\mem[13][0] ),
    .B(\mem[15][0] ),
    .S(_0247_),
    .Z(_0267_));
 NOR3_X1 _0895_ (.A1(_0256_),
    .A2(_0260_),
    .A3(_0267_),
    .ZN(_0268_));
 NOR4_X1 _0896_ (.A1(_0262_),
    .A2(_0264_),
    .A3(_0266_),
    .A4(_0268_),
    .ZN(_0269_));
 BUF_X4 _0897_ (.A(\rd_ptr_bin[3] ),
    .Z(_0270_));
 MUX2_X1 _0898_ (.A(_0257_),
    .B(_0269_),
    .S(_0270_),
    .Z(_0271_));
 INV_X1 _0899_ (.A(net9),
    .ZN(_0272_));
 NAND2_X2 _0900_ (.A1(net2),
    .A2(_0272_),
    .ZN(_0273_));
 CLKBUF_X3 _0901_ (.A(_0273_),
    .Z(_0274_));
 CLKBUF_X3 _0902_ (.A(_0274_),
    .Z(_0275_));
 MUX2_X1 _0903_ (.A(_0271_),
    .B(net17),
    .S(_0275_),
    .Z(_0143_));
 CLKBUF_X3 _0904_ (.A(_0251_),
    .Z(_0276_));
 AND3_X2 _0905_ (.A1(_0248_),
    .A2(_0276_),
    .A3(_0270_),
    .ZN(_0277_));
 CLKBUF_X3 _0906_ (.A(_0254_),
    .Z(_0278_));
 MUX2_X1 _0907_ (.A(\mem[14][1] ),
    .B(\mem[15][1] ),
    .S(_0278_),
    .Z(_0279_));
 INV_X1 _0908_ (.A(_0247_),
    .ZN(_0280_));
 AND3_X2 _0909_ (.A1(_0280_),
    .A2(_0259_),
    .A3(_0270_),
    .ZN(_0281_));
 MUX2_X1 _0910_ (.A(\mem[12][1] ),
    .B(\mem[13][1] ),
    .S(_0278_),
    .Z(_0282_));
 AOI221_X1 _0911_ (.A(_0274_),
    .B1(_0277_),
    .B2(_0279_),
    .C1(_0281_),
    .C2(_0282_),
    .ZN(_0283_));
 BUF_X4 _0912_ (.A(_0247_),
    .Z(_0284_));
 MUX2_X1 _0913_ (.A(\mem[8][1] ),
    .B(\mem[10][1] ),
    .S(_0284_),
    .Z(_0285_));
 MUX2_X1 _0914_ (.A(\mem[9][1] ),
    .B(\mem[11][1] ),
    .S(_0284_),
    .Z(_0286_));
 MUX2_X1 _0915_ (.A(_0285_),
    .B(_0286_),
    .S(_0258_),
    .Z(_0287_));
 AND2_X2 _0916_ (.A1(_0260_),
    .A2(_0270_),
    .ZN(_0288_));
 NAND2_X1 _0917_ (.A1(_0287_),
    .A2(_0288_),
    .ZN(_0289_));
 NOR2_X4 _0918_ (.A1(_0280_),
    .A2(_0270_),
    .ZN(_0290_));
 CLKBUF_X3 _0919_ (.A(_0251_),
    .Z(_0291_));
 MUX2_X1 _0920_ (.A(\mem[2][1] ),
    .B(\mem[6][1] ),
    .S(_0291_),
    .Z(_0292_));
 MUX2_X1 _0921_ (.A(\mem[3][1] ),
    .B(\mem[7][1] ),
    .S(_0259_),
    .Z(_0293_));
 CLKBUF_X3 _0922_ (.A(_0278_),
    .Z(_0294_));
 MUX2_X1 _0923_ (.A(_0292_),
    .B(_0293_),
    .S(_0294_),
    .Z(_0295_));
 MUX2_X1 _0924_ (.A(\mem[0][1] ),
    .B(\mem[4][1] ),
    .S(_0276_),
    .Z(_0296_));
 MUX2_X1 _0925_ (.A(\mem[1][1] ),
    .B(\mem[5][1] ),
    .S(_0276_),
    .Z(_0297_));
 MUX2_X1 _0926_ (.A(_0296_),
    .B(_0297_),
    .S(_0294_),
    .Z(_0298_));
 NOR2_X4 _0927_ (.A1(_0284_),
    .A2(_0270_),
    .ZN(_0299_));
 AOI22_X1 _0928_ (.A1(_0290_),
    .A2(_0295_),
    .B1(_0298_),
    .B2(_0299_),
    .ZN(_0300_));
 AND3_X1 _0929_ (.A1(_0283_),
    .A2(_0289_),
    .A3(_0300_),
    .ZN(_0301_));
 INV_X1 _0930_ (.A(net18),
    .ZN(_0302_));
 AOI21_X1 _0931_ (.A(_0301_),
    .B1(_0275_),
    .B2(_0302_),
    .ZN(_0144_));
 MUX2_X1 _0932_ (.A(\mem[14][2] ),
    .B(\mem[15][2] ),
    .S(_0278_),
    .Z(_0303_));
 MUX2_X1 _0933_ (.A(\mem[12][2] ),
    .B(\mem[13][2] ),
    .S(_0255_),
    .Z(_0304_));
 AOI221_X1 _0934_ (.A(_0273_),
    .B1(_0277_),
    .B2(_0303_),
    .C1(_0304_),
    .C2(_0281_),
    .ZN(_0305_));
 MUX2_X1 _0935_ (.A(\mem[8][2] ),
    .B(\mem[10][2] ),
    .S(_0248_),
    .Z(_0306_));
 MUX2_X1 _0936_ (.A(\mem[9][2] ),
    .B(\mem[11][2] ),
    .S(_0284_),
    .Z(_0307_));
 MUX2_X1 _0937_ (.A(_0306_),
    .B(_0307_),
    .S(_0258_),
    .Z(_0308_));
 NAND2_X1 _0938_ (.A1(_0288_),
    .A2(_0308_),
    .ZN(_0309_));
 MUX2_X1 _0939_ (.A(\mem[2][2] ),
    .B(\mem[6][2] ),
    .S(_0291_),
    .Z(_0310_));
 MUX2_X1 _0940_ (.A(\mem[3][2] ),
    .B(\mem[7][2] ),
    .S(_0259_),
    .Z(_0311_));
 MUX2_X1 _0941_ (.A(_0310_),
    .B(_0311_),
    .S(_0294_),
    .Z(_0312_));
 MUX2_X1 _0942_ (.A(\mem[0][2] ),
    .B(\mem[4][2] ),
    .S(_0251_),
    .Z(_0313_));
 MUX2_X1 _0943_ (.A(\mem[1][2] ),
    .B(\mem[5][2] ),
    .S(_0276_),
    .Z(_0314_));
 MUX2_X1 _0944_ (.A(_0313_),
    .B(_0314_),
    .S(_0294_),
    .Z(_0315_));
 AOI22_X1 _0945_ (.A1(_0290_),
    .A2(_0312_),
    .B1(_0315_),
    .B2(_0299_),
    .ZN(_0316_));
 AND3_X1 _0946_ (.A1(_0305_),
    .A2(_0309_),
    .A3(_0316_),
    .ZN(_0317_));
 INV_X1 _0947_ (.A(net19),
    .ZN(_0318_));
 AOI21_X1 _0948_ (.A(_0317_),
    .B1(_0275_),
    .B2(_0318_),
    .ZN(_0145_));
 MUX2_X1 _0949_ (.A(\mem[14][3] ),
    .B(\mem[15][3] ),
    .S(_0278_),
    .Z(_0319_));
 MUX2_X1 _0950_ (.A(\mem[12][3] ),
    .B(\mem[13][3] ),
    .S(_0255_),
    .Z(_0320_));
 AOI221_X1 _0951_ (.A(_0273_),
    .B1(_0277_),
    .B2(_0319_),
    .C1(_0320_),
    .C2(_0281_),
    .ZN(_0321_));
 MUX2_X1 _0952_ (.A(\mem[8][3] ),
    .B(\mem[10][3] ),
    .S(_0248_),
    .Z(_0322_));
 MUX2_X1 _0953_ (.A(\mem[9][3] ),
    .B(\mem[11][3] ),
    .S(_0284_),
    .Z(_0323_));
 MUX2_X1 _0954_ (.A(_0322_),
    .B(_0323_),
    .S(_0258_),
    .Z(_0324_));
 NAND2_X1 _0955_ (.A1(_0288_),
    .A2(_0324_),
    .ZN(_0325_));
 MUX2_X1 _0956_ (.A(\mem[2][3] ),
    .B(\mem[6][3] ),
    .S(_0291_),
    .Z(_0326_));
 MUX2_X1 _0957_ (.A(\mem[3][3] ),
    .B(\mem[7][3] ),
    .S(_0259_),
    .Z(_0327_));
 MUX2_X1 _0958_ (.A(_0326_),
    .B(_0327_),
    .S(_0294_),
    .Z(_0328_));
 MUX2_X1 _0959_ (.A(\mem[0][3] ),
    .B(\mem[4][3] ),
    .S(_0251_),
    .Z(_0329_));
 MUX2_X1 _0960_ (.A(\mem[1][3] ),
    .B(\mem[5][3] ),
    .S(_0276_),
    .Z(_0330_));
 MUX2_X1 _0961_ (.A(_0329_),
    .B(_0330_),
    .S(_0294_),
    .Z(_0331_));
 AOI22_X1 _0962_ (.A1(_0290_),
    .A2(_0328_),
    .B1(_0331_),
    .B2(_0299_),
    .ZN(_0332_));
 AND3_X1 _0963_ (.A1(_0321_),
    .A2(_0325_),
    .A3(_0332_),
    .ZN(_0333_));
 INV_X1 _0964_ (.A(net20),
    .ZN(_0334_));
 AOI21_X1 _0965_ (.A(_0333_),
    .B1(_0275_),
    .B2(_0334_),
    .ZN(_0146_));
 MUX2_X1 _0966_ (.A(\mem[14][4] ),
    .B(\mem[15][4] ),
    .S(_0278_),
    .Z(_0335_));
 MUX2_X1 _0967_ (.A(\mem[12][4] ),
    .B(\mem[13][4] ),
    .S(_0278_),
    .Z(_0336_));
 AOI221_X1 _0968_ (.A(_0273_),
    .B1(_0277_),
    .B2(_0335_),
    .C1(_0336_),
    .C2(_0281_),
    .ZN(_0337_));
 MUX2_X1 _0969_ (.A(\mem[8][4] ),
    .B(\mem[10][4] ),
    .S(_0248_),
    .Z(_0338_));
 MUX2_X1 _0970_ (.A(\mem[9][4] ),
    .B(\mem[11][4] ),
    .S(_0284_),
    .Z(_0339_));
 MUX2_X1 _0971_ (.A(_0338_),
    .B(_0339_),
    .S(_0258_),
    .Z(_0340_));
 NAND2_X1 _0972_ (.A1(_0288_),
    .A2(_0340_),
    .ZN(_0341_));
 MUX2_X1 _0973_ (.A(\mem[2][4] ),
    .B(\mem[6][4] ),
    .S(_0291_),
    .Z(_0342_));
 MUX2_X1 _0974_ (.A(\mem[3][4] ),
    .B(\mem[7][4] ),
    .S(_0291_),
    .Z(_0343_));
 MUX2_X1 _0975_ (.A(_0342_),
    .B(_0343_),
    .S(_0294_),
    .Z(_0344_));
 MUX2_X1 _0976_ (.A(\mem[0][4] ),
    .B(\mem[4][4] ),
    .S(_0251_),
    .Z(_0345_));
 MUX2_X1 _0977_ (.A(\mem[1][4] ),
    .B(\mem[5][4] ),
    .S(_0276_),
    .Z(_0346_));
 MUX2_X1 _0978_ (.A(_0345_),
    .B(_0346_),
    .S(_0255_),
    .Z(_0347_));
 AOI22_X1 _0979_ (.A1(_0290_),
    .A2(_0344_),
    .B1(_0347_),
    .B2(_0299_),
    .ZN(_0348_));
 AND3_X1 _0980_ (.A1(_0337_),
    .A2(_0341_),
    .A3(_0348_),
    .ZN(_0349_));
 INV_X1 _0981_ (.A(net21),
    .ZN(_0350_));
 AOI21_X1 _0982_ (.A(_0349_),
    .B1(_0275_),
    .B2(_0350_),
    .ZN(_0147_));
 MUX2_X1 _0983_ (.A(\mem[14][5] ),
    .B(\mem[15][5] ),
    .S(_0254_),
    .Z(_0351_));
 MUX2_X1 _0984_ (.A(\mem[12][5] ),
    .B(\mem[13][5] ),
    .S(_0278_),
    .Z(_0352_));
 AOI221_X1 _0985_ (.A(_0273_),
    .B1(_0277_),
    .B2(_0351_),
    .C1(_0352_),
    .C2(_0281_),
    .ZN(_0353_));
 MUX2_X1 _0986_ (.A(\mem[8][5] ),
    .B(\mem[10][5] ),
    .S(_0248_),
    .Z(_0354_));
 MUX2_X1 _0987_ (.A(\mem[9][5] ),
    .B(\mem[11][5] ),
    .S(_0284_),
    .Z(_0355_));
 MUX2_X1 _0988_ (.A(_0354_),
    .B(_0355_),
    .S(_0258_),
    .Z(_0356_));
 NAND2_X1 _0989_ (.A1(_0288_),
    .A2(_0356_),
    .ZN(_0357_));
 MUX2_X1 _0990_ (.A(\mem[2][5] ),
    .B(\mem[6][5] ),
    .S(_0291_),
    .Z(_0358_));
 MUX2_X1 _0991_ (.A(\mem[3][5] ),
    .B(\mem[7][5] ),
    .S(_0291_),
    .Z(_0359_));
 MUX2_X1 _0992_ (.A(_0358_),
    .B(_0359_),
    .S(_0294_),
    .Z(_0360_));
 MUX2_X1 _0993_ (.A(\mem[0][5] ),
    .B(\mem[4][5] ),
    .S(_0251_),
    .Z(_0361_));
 MUX2_X1 _0994_ (.A(\mem[1][5] ),
    .B(\mem[5][5] ),
    .S(_0276_),
    .Z(_0362_));
 MUX2_X1 _0995_ (.A(_0361_),
    .B(_0362_),
    .S(_0255_),
    .Z(_0363_));
 AOI22_X1 _0996_ (.A1(_0290_),
    .A2(_0360_),
    .B1(_0363_),
    .B2(_0299_),
    .ZN(_0364_));
 AND3_X1 _0997_ (.A1(_0353_),
    .A2(_0357_),
    .A3(_0364_),
    .ZN(_0365_));
 INV_X1 _0998_ (.A(net22),
    .ZN(_0366_));
 AOI21_X1 _0999_ (.A(_0365_),
    .B1(_0275_),
    .B2(_0366_),
    .ZN(_0148_));
 MUX2_X1 _1000_ (.A(\mem[14][6] ),
    .B(\mem[15][6] ),
    .S(_0254_),
    .Z(_0367_));
 MUX2_X1 _1001_ (.A(\mem[12][6] ),
    .B(\mem[13][6] ),
    .S(_0278_),
    .Z(_0368_));
 AOI221_X1 _1002_ (.A(_0273_),
    .B1(_0277_),
    .B2(_0367_),
    .C1(_0368_),
    .C2(_0281_),
    .ZN(_0369_));
 MUX2_X1 _1003_ (.A(\mem[8][6] ),
    .B(\mem[10][6] ),
    .S(_0248_),
    .Z(_0370_));
 MUX2_X1 _1004_ (.A(\mem[9][6] ),
    .B(\mem[11][6] ),
    .S(_0284_),
    .Z(_0371_));
 MUX2_X1 _1005_ (.A(_0370_),
    .B(_0371_),
    .S(_0258_),
    .Z(_0372_));
 NAND2_X1 _1006_ (.A1(_0288_),
    .A2(_0372_),
    .ZN(_0373_));
 MUX2_X1 _1007_ (.A(\mem[2][6] ),
    .B(\mem[6][6] ),
    .S(_0291_),
    .Z(_0374_));
 MUX2_X1 _1008_ (.A(\mem[3][6] ),
    .B(\mem[7][6] ),
    .S(_0291_),
    .Z(_0375_));
 MUX2_X1 _1009_ (.A(_0374_),
    .B(_0375_),
    .S(_0294_),
    .Z(_0376_));
 MUX2_X1 _1010_ (.A(\mem[0][6] ),
    .B(\mem[4][6] ),
    .S(_0251_),
    .Z(_0377_));
 MUX2_X1 _1011_ (.A(\mem[1][6] ),
    .B(\mem[5][6] ),
    .S(_0276_),
    .Z(_0378_));
 MUX2_X1 _1012_ (.A(_0377_),
    .B(_0378_),
    .S(_0255_),
    .Z(_0379_));
 AOI22_X1 _1013_ (.A1(_0290_),
    .A2(_0376_),
    .B1(_0379_),
    .B2(_0299_),
    .ZN(_0380_));
 AND3_X1 _1014_ (.A1(_0369_),
    .A2(_0373_),
    .A3(_0380_),
    .ZN(_0381_));
 INV_X1 _1015_ (.A(net23),
    .ZN(_0382_));
 AOI21_X1 _1016_ (.A(_0381_),
    .B1(_0275_),
    .B2(_0382_),
    .ZN(_0149_));
 MUX2_X1 _1017_ (.A(\mem[14][7] ),
    .B(\mem[15][7] ),
    .S(_0254_),
    .Z(_0383_));
 MUX2_X1 _1018_ (.A(\mem[12][7] ),
    .B(\mem[13][7] ),
    .S(_0278_),
    .Z(_0384_));
 AOI221_X1 _1019_ (.A(_0273_),
    .B1(_0277_),
    .B2(_0383_),
    .C1(_0384_),
    .C2(_0281_),
    .ZN(_0385_));
 MUX2_X1 _1020_ (.A(\mem[8][7] ),
    .B(\mem[10][7] ),
    .S(_0248_),
    .Z(_0386_));
 MUX2_X1 _1021_ (.A(\mem[9][7] ),
    .B(\mem[11][7] ),
    .S(_0248_),
    .Z(_0387_));
 MUX2_X1 _1022_ (.A(_0386_),
    .B(_0387_),
    .S(_0258_),
    .Z(_0388_));
 NAND2_X1 _1023_ (.A1(_0288_),
    .A2(_0388_),
    .ZN(_0389_));
 MUX2_X1 _1024_ (.A(\mem[2][7] ),
    .B(\mem[6][7] ),
    .S(_0276_),
    .Z(_0390_));
 MUX2_X1 _1025_ (.A(\mem[3][7] ),
    .B(\mem[7][7] ),
    .S(_0291_),
    .Z(_0391_));
 MUX2_X1 _1026_ (.A(_0390_),
    .B(_0391_),
    .S(_0294_),
    .Z(_0392_));
 MUX2_X1 _1027_ (.A(\mem[0][7] ),
    .B(\mem[4][7] ),
    .S(_0251_),
    .Z(_0393_));
 MUX2_X1 _1028_ (.A(\mem[1][7] ),
    .B(\mem[5][7] ),
    .S(_0276_),
    .Z(_0394_));
 MUX2_X1 _1029_ (.A(_0393_),
    .B(_0394_),
    .S(_0255_),
    .Z(_0395_));
 AOI22_X1 _1030_ (.A1(_0290_),
    .A2(_0392_),
    .B1(_0395_),
    .B2(_0299_),
    .ZN(_0396_));
 AND3_X1 _1031_ (.A1(_0385_),
    .A2(_0389_),
    .A3(_0396_),
    .ZN(_0397_));
 INV_X1 _1032_ (.A(net24),
    .ZN(_0398_));
 AOI21_X1 _1033_ (.A(_0397_),
    .B1(_0275_),
    .B2(_0398_),
    .ZN(_0150_));
 MUX2_X1 _1034_ (.A(_0013_),
    .B(_0258_),
    .S(_0274_),
    .Z(_0151_));
 MUX2_X1 _1035_ (.A(_0014_),
    .B(_0284_),
    .S(_0274_),
    .Z(_0152_));
 NAND2_X1 _1036_ (.A1(_0259_),
    .A2(_0275_),
    .ZN(_0399_));
 XOR2_X2 _1037_ (.A(_0639_),
    .B(_0611_),
    .Z(_0400_));
 OAI21_X1 _1038_ (.A(_0399_),
    .B1(_0400_),
    .B2(_0275_),
    .ZN(_0153_));
 NAND3_X1 _1039_ (.A1(_0255_),
    .A2(_0284_),
    .A3(_0259_),
    .ZN(_0401_));
 XOR2_X2 _1040_ (.A(_0601_),
    .B(_0401_),
    .Z(_0402_));
 MUX2_X1 _1041_ (.A(_0402_),
    .B(_0270_),
    .S(_0274_),
    .Z(_0154_));
 XNOR2_X1 _1042_ (.A(_0258_),
    .B(_0014_),
    .ZN(_0403_));
 MUX2_X1 _1043_ (.A(_0403_),
    .B(\rd_ptr_gray[0] ),
    .S(_0274_),
    .Z(_0155_));
 XNOR2_X1 _1044_ (.A(_0014_),
    .B(_0400_),
    .ZN(_0404_));
 MUX2_X1 _1045_ (.A(_0404_),
    .B(\rd_ptr_gray[1] ),
    .S(_0274_),
    .Z(_0156_));
 XNOR2_X1 _1046_ (.A(_0400_),
    .B(_0402_),
    .ZN(_0405_));
 MUX2_X1 _1047_ (.A(_0405_),
    .B(\rd_ptr_gray[2] ),
    .S(_0274_),
    .Z(_0157_));
 NAND3_X1 _1048_ (.A1(_0259_),
    .A2(_0270_),
    .A3(_0639_),
    .ZN(_0406_));
 XOR2_X1 _1049_ (.A(\rd_ptr_bin[4] ),
    .B(_0406_),
    .Z(_0407_));
 XNOR2_X1 _1050_ (.A(_0402_),
    .B(_0407_),
    .ZN(_0408_));
 MUX2_X1 _1051_ (.A(_0408_),
    .B(\rd_ptr_gray[3] ),
    .S(_0274_),
    .Z(_0158_));
 NOR2_X1 _1052_ (.A1(_0274_),
    .A2(_0406_),
    .ZN(_0409_));
 XOR2_X1 _1053_ (.A(\rd_ptr_bin[4] ),
    .B(_0409_),
    .Z(_0159_));
 MUX2_X1 _1054_ (.A(\wr_ptr_bin[0] ),
    .B(_0011_),
    .S(_0224_),
    .Z(_0160_));
 MUX2_X1 _1055_ (.A(\wr_ptr_bin[1] ),
    .B(_0012_),
    .S(_0224_),
    .Z(_0161_));
 XNOR2_X1 _1056_ (.A(_0192_),
    .B(_0222_),
    .ZN(_0162_));
 NAND4_X1 _1057_ (.A1(_0192_),
    .A2(\wr_ptr_bin[1] ),
    .A3(\wr_ptr_bin[0] ),
    .A4(_0224_),
    .ZN(_0410_));
 XNOR2_X1 _1058_ (.A(_0191_),
    .B(_0410_),
    .ZN(_0163_));
 XNOR2_X1 _1059_ (.A(\wr_ptr_bin[0] ),
    .B(_0012_),
    .ZN(_0411_));
 MUX2_X1 _1060_ (.A(\wr_ptr_gray[0] ),
    .B(_0411_),
    .S(_0224_),
    .Z(_0164_));
 XNOR2_X1 _1061_ (.A(_0221_),
    .B(_0012_),
    .ZN(_0412_));
 XNOR2_X1 _1062_ (.A(_0192_),
    .B(_0412_),
    .ZN(_0413_));
 MUX2_X1 _1063_ (.A(\wr_ptr_gray[1] ),
    .B(_0413_),
    .S(_0224_),
    .Z(_0165_));
 XOR2_X1 _1064_ (.A(_0191_),
    .B(_0221_),
    .Z(_0414_));
 NAND2_X1 _1065_ (.A1(\wr_ptr_bin[1] ),
    .A2(\wr_ptr_bin[0] ),
    .ZN(_0415_));
 NAND2_X1 _1066_ (.A1(_0192_),
    .A2(_0415_),
    .ZN(_0416_));
 XNOR2_X1 _1067_ (.A(_0414_),
    .B(_0416_),
    .ZN(_0417_));
 MUX2_X1 _1068_ (.A(\wr_ptr_gray[2] ),
    .B(_0417_),
    .S(_0224_),
    .Z(_0166_));
 INV_X1 _1069_ (.A(_0221_),
    .ZN(_0418_));
 OAI21_X1 _1070_ (.A(_0191_),
    .B1(_0216_),
    .B2(_0418_),
    .ZN(_0419_));
 NOR3_X1 _1071_ (.A1(_0225_),
    .A2(_0216_),
    .A3(_0415_),
    .ZN(_0420_));
 AOI221_X2 _1072_ (.A(_0193_),
    .B1(_0415_),
    .B2(_0419_),
    .C1(_0420_),
    .C2(_0418_),
    .ZN(_0421_));
 XOR2_X1 _1073_ (.A(\wr_ptr_bin[4] ),
    .B(_0421_),
    .Z(_0422_));
 MUX2_X1 _1074_ (.A(\wr_ptr_gray[3] ),
    .B(_0422_),
    .S(_0224_),
    .Z(_0167_));
 XNOR2_X1 _1075_ (.A(\wr_ptr_bin[4] ),
    .B(_0231_),
    .ZN(_0168_));
 AND2_X1 _1076_ (.A1(net12),
    .A2(net13),
    .ZN(_0423_));
 NOR4_X1 _1077_ (.A1(net16),
    .A2(net14),
    .A3(net15),
    .A4(_0423_),
    .ZN(net7));
 XOR2_X1 _1078_ (.A(_0182_),
    .B(_0600_),
    .Z(net28));
 NAND2_X1 _1079_ (.A1(net27),
    .A2(net28),
    .ZN(_0424_));
 OAI21_X1 _1080_ (.A(_0188_),
    .B1(_0424_),
    .B2(_0184_),
    .ZN(net8));
 FA_X1 _1081_ (.A(_0595_),
    .B(\wr_ptr_sync[1] ),
    .CI(_0596_),
    .CO(_0597_),
    .S(net13));
 FA_X1 _1082_ (.A(_0598_),
    .B(\wr_ptr_bin[1] ),
    .CI(_0599_),
    .CO(_0600_),
    .S(net27));
 HA_X1 _1083_ (.A(_0601_),
    .B(\wr_ptr_sync[3] ),
    .CO(_0602_),
    .S(_0603_));
 HA_X1 _1084_ (.A(\rd_ptr_bin[4] ),
    .B(_0605_),
    .CO(_0606_),
    .S(_0607_));
 HA_X1 _1085_ (.A(_0595_),
    .B(\wr_ptr_sync[1] ),
    .CO(_0608_),
    .S(_0609_));
 HA_X1 _1086_ (.A(_0611_),
    .B(\wr_ptr_sync[2] ),
    .CO(_0612_),
    .S(_0613_));
 HA_X1 _1087_ (.A(_0013_),
    .B(\wr_ptr_sync[0] ),
    .CO(_0615_),
    .S(_0616_));
 HA_X1 _1088_ (.A(\rd_ptr_bin[0] ),
    .B(_0617_),
    .CO(_0618_),
    .S(_0619_));
 HA_X1 _1089_ (.A(_0621_),
    .B(\wr_ptr_bin[0] ),
    .CO(_0622_),
    .S(_0623_));
 HA_X1 _1090_ (.A(\rd_ptr_sync[0] ),
    .B(_0011_),
    .CO(_0624_),
    .S(_0625_));
 HA_X1 _1091_ (.A(_0598_),
    .B(\wr_ptr_bin[1] ),
    .CO(_0626_),
    .S(_0620_));
 HA_X1 _1092_ (.A(_0628_),
    .B(\wr_ptr_bin[2] ),
    .CO(_0629_),
    .S(_0630_));
 HA_X1 _1093_ (.A(_0632_),
    .B(\wr_ptr_bin[3] ),
    .CO(_0633_),
    .S(_0634_));
 HA_X1 _1094_ (.A(\rd_ptr_sync[4] ),
    .B(_0636_),
    .CO(_0637_),
    .S(_0638_));
 HA_X1 _1095_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .CO(_0639_),
    .S(_0014_));
 HA_X1 _1096_ (.A(_0011_),
    .B(_0627_),
    .CO(_0640_),
    .S(_0012_));
 HA_X1 _1097_ (.A(_0011_),
    .B(\wr_ptr_bin[1] ),
    .CO(_0641_),
    .S(_0642_));
 HA_X1 _1098_ (.A(\wr_ptr_bin[0] ),
    .B(_0627_),
    .CO(_0643_),
    .S(_0644_));
 HA_X1 _1099_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .CO(_0645_),
    .S(_0646_));
 FILLCELL_X32 FILLER_0_1 ();
 DFFS_X1 \empty_reg$_DFF_PN1_  (.D(_0000_),
    .SN(net3),
    .CK(net1),
    .Q(net9),
    .QN(_0571_));
 DFFR_X1 \full_reg$_DFF_PN0_  (.D(_0001_),
    .RN(net6),
    .CK(net4),
    .Q(net10),
    .QN(_0570_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0015_),
    .CK(net4),
    .Q(\mem[0][0] ),
    .QN(_0569_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0016_),
    .CK(net4),
    .Q(\mem[0][1] ),
    .QN(_0568_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0017_),
    .CK(net4),
    .Q(\mem[0][2] ),
    .QN(_0567_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0018_),
    .CK(net4),
    .Q(\mem[0][3] ),
    .QN(_0566_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0019_),
    .CK(net4),
    .Q(\mem[0][4] ),
    .QN(_0565_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0020_),
    .CK(net4),
    .Q(\mem[0][5] ),
    .QN(_0564_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0021_),
    .CK(net4),
    .Q(\mem[0][6] ),
    .QN(_0563_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0022_),
    .CK(net4),
    .Q(\mem[0][7] ),
    .QN(_0562_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0023_),
    .CK(net4),
    .Q(\mem[10][0] ),
    .QN(_0561_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0024_),
    .CK(net4),
    .Q(\mem[10][1] ),
    .QN(_0560_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0025_),
    .CK(net4),
    .Q(\mem[10][2] ),
    .QN(_0559_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0026_),
    .CK(net4),
    .Q(\mem[10][3] ),
    .QN(_0558_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0027_),
    .CK(net4),
    .Q(\mem[10][4] ),
    .QN(_0557_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0028_),
    .CK(net4),
    .Q(\mem[10][5] ),
    .QN(_0556_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0029_),
    .CK(net4),
    .Q(\mem[10][6] ),
    .QN(_0555_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0030_),
    .CK(net4),
    .Q(\mem[10][7] ),
    .QN(_0554_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0031_),
    .CK(net4),
    .Q(\mem[11][0] ),
    .QN(_0553_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0032_),
    .CK(net4),
    .Q(\mem[11][1] ),
    .QN(_0552_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0033_),
    .CK(net4),
    .Q(\mem[11][2] ),
    .QN(_0551_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0034_),
    .CK(net4),
    .Q(\mem[11][3] ),
    .QN(_0550_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0035_),
    .CK(net4),
    .Q(\mem[11][4] ),
    .QN(_0549_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0036_),
    .CK(net4),
    .Q(\mem[11][5] ),
    .QN(_0548_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0037_),
    .CK(net4),
    .Q(\mem[11][6] ),
    .QN(_0547_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0038_),
    .CK(net4),
    .Q(\mem[11][7] ),
    .QN(_0546_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0039_),
    .CK(net4),
    .Q(\mem[12][0] ),
    .QN(_0545_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0040_),
    .CK(net4),
    .Q(\mem[12][1] ),
    .QN(_0544_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0041_),
    .CK(net4),
    .Q(\mem[12][2] ),
    .QN(_0543_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0042_),
    .CK(net4),
    .Q(\mem[12][3] ),
    .QN(_0542_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0043_),
    .CK(net4),
    .Q(\mem[12][4] ),
    .QN(_0541_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0044_),
    .CK(net4),
    .Q(\mem[12][5] ),
    .QN(_0540_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0045_),
    .CK(net4),
    .Q(\mem[12][6] ),
    .QN(_0539_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0046_),
    .CK(net4),
    .Q(\mem[12][7] ),
    .QN(_0538_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0047_),
    .CK(net4),
    .Q(\mem[13][0] ),
    .QN(_0537_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0048_),
    .CK(net4),
    .Q(\mem[13][1] ),
    .QN(_0536_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0049_),
    .CK(net4),
    .Q(\mem[13][2] ),
    .QN(_0535_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0050_),
    .CK(net4),
    .Q(\mem[13][3] ),
    .QN(_0534_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0051_),
    .CK(net4),
    .Q(\mem[13][4] ),
    .QN(_0533_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0052_),
    .CK(net4),
    .Q(\mem[13][5] ),
    .QN(_0532_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0053_),
    .CK(net4),
    .Q(\mem[13][6] ),
    .QN(_0531_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0054_),
    .CK(net4),
    .Q(\mem[13][7] ),
    .QN(_0530_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0055_),
    .CK(net4),
    .Q(\mem[14][0] ),
    .QN(_0529_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0056_),
    .CK(net4),
    .Q(\mem[14][1] ),
    .QN(_0528_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0057_),
    .CK(net4),
    .Q(\mem[14][2] ),
    .QN(_0527_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0058_),
    .CK(net4),
    .Q(\mem[14][3] ),
    .QN(_0526_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0059_),
    .CK(net4),
    .Q(\mem[14][4] ),
    .QN(_0525_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0060_),
    .CK(net4),
    .Q(\mem[14][5] ),
    .QN(_0524_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0061_),
    .CK(net4),
    .Q(\mem[14][6] ),
    .QN(_0523_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0062_),
    .CK(net4),
    .Q(\mem[14][7] ),
    .QN(_0522_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0063_),
    .CK(net4),
    .Q(\mem[15][0] ),
    .QN(_0521_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0064_),
    .CK(net4),
    .Q(\mem[15][1] ),
    .QN(_0520_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0065_),
    .CK(net4),
    .Q(\mem[15][2] ),
    .QN(_0519_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0066_),
    .CK(net4),
    .Q(\mem[15][3] ),
    .QN(_0518_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0067_),
    .CK(net4),
    .Q(\mem[15][4] ),
    .QN(_0517_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0068_),
    .CK(net4),
    .Q(\mem[15][5] ),
    .QN(_0516_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0069_),
    .CK(net4),
    .Q(\mem[15][6] ),
    .QN(_0515_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0070_),
    .CK(net4),
    .Q(\mem[15][7] ),
    .QN(_0514_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0071_),
    .CK(net4),
    .Q(\mem[1][0] ),
    .QN(_0513_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0072_),
    .CK(net4),
    .Q(\mem[1][1] ),
    .QN(_0512_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0073_),
    .CK(net4),
    .Q(\mem[1][2] ),
    .QN(_0511_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0074_),
    .CK(net4),
    .Q(\mem[1][3] ),
    .QN(_0510_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0075_),
    .CK(net4),
    .Q(\mem[1][4] ),
    .QN(_0509_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0076_),
    .CK(net4),
    .Q(\mem[1][5] ),
    .QN(_0508_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0077_),
    .CK(net4),
    .Q(\mem[1][6] ),
    .QN(_0507_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0078_),
    .CK(net4),
    .Q(\mem[1][7] ),
    .QN(_0506_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0079_),
    .CK(net4),
    .Q(\mem[2][0] ),
    .QN(_0505_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0080_),
    .CK(net4),
    .Q(\mem[2][1] ),
    .QN(_0504_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0081_),
    .CK(net4),
    .Q(\mem[2][2] ),
    .QN(_0503_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0082_),
    .CK(net4),
    .Q(\mem[2][3] ),
    .QN(_0502_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0083_),
    .CK(net4),
    .Q(\mem[2][4] ),
    .QN(_0501_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0084_),
    .CK(net4),
    .Q(\mem[2][5] ),
    .QN(_0500_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0085_),
    .CK(net4),
    .Q(\mem[2][6] ),
    .QN(_0499_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0086_),
    .CK(net4),
    .Q(\mem[2][7] ),
    .QN(_0498_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0087_),
    .CK(net4),
    .Q(\mem[3][0] ),
    .QN(_0497_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0088_),
    .CK(net4),
    .Q(\mem[3][1] ),
    .QN(_0496_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0089_),
    .CK(net4),
    .Q(\mem[3][2] ),
    .QN(_0495_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0090_),
    .CK(net4),
    .Q(\mem[3][3] ),
    .QN(_0494_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0091_),
    .CK(net4),
    .Q(\mem[3][4] ),
    .QN(_0493_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0092_),
    .CK(net4),
    .Q(\mem[3][5] ),
    .QN(_0492_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0093_),
    .CK(net4),
    .Q(\mem[3][6] ),
    .QN(_0491_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0094_),
    .CK(net4),
    .Q(\mem[3][7] ),
    .QN(_0490_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0095_),
    .CK(net4),
    .Q(\mem[4][0] ),
    .QN(_0489_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0096_),
    .CK(net4),
    .Q(\mem[4][1] ),
    .QN(_0488_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0097_),
    .CK(net4),
    .Q(\mem[4][2] ),
    .QN(_0487_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0098_),
    .CK(net4),
    .Q(\mem[4][3] ),
    .QN(_0486_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0099_),
    .CK(net4),
    .Q(\mem[4][4] ),
    .QN(_0485_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0100_),
    .CK(net4),
    .Q(\mem[4][5] ),
    .QN(_0484_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0101_),
    .CK(net4),
    .Q(\mem[4][6] ),
    .QN(_0483_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0102_),
    .CK(net4),
    .Q(\mem[4][7] ),
    .QN(_0482_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0103_),
    .CK(net4),
    .Q(\mem[5][0] ),
    .QN(_0481_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0104_),
    .CK(net4),
    .Q(\mem[5][1] ),
    .QN(_0480_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0105_),
    .CK(net4),
    .Q(\mem[5][2] ),
    .QN(_0479_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0106_),
    .CK(net4),
    .Q(\mem[5][3] ),
    .QN(_0478_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0107_),
    .CK(net4),
    .Q(\mem[5][4] ),
    .QN(_0477_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0108_),
    .CK(net4),
    .Q(\mem[5][5] ),
    .QN(_0476_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0109_),
    .CK(net4),
    .Q(\mem[5][6] ),
    .QN(_0475_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0110_),
    .CK(net4),
    .Q(\mem[5][7] ),
    .QN(_0474_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0111_),
    .CK(net4),
    .Q(\mem[6][0] ),
    .QN(_0473_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0112_),
    .CK(net4),
    .Q(\mem[6][1] ),
    .QN(_0472_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0113_),
    .CK(net4),
    .Q(\mem[6][2] ),
    .QN(_0471_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0114_),
    .CK(net4),
    .Q(\mem[6][3] ),
    .QN(_0470_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0115_),
    .CK(net4),
    .Q(\mem[6][4] ),
    .QN(_0469_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0116_),
    .CK(net4),
    .Q(\mem[6][5] ),
    .QN(_0468_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0117_),
    .CK(net4),
    .Q(\mem[6][6] ),
    .QN(_0467_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0118_),
    .CK(net4),
    .Q(\mem[6][7] ),
    .QN(_0466_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0119_),
    .CK(net4),
    .Q(\mem[7][0] ),
    .QN(_0465_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0120_),
    .CK(net4),
    .Q(\mem[7][1] ),
    .QN(_0464_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0121_),
    .CK(net4),
    .Q(\mem[7][2] ),
    .QN(_0463_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0122_),
    .CK(net4),
    .Q(\mem[7][3] ),
    .QN(_0462_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0123_),
    .CK(net4),
    .Q(\mem[7][4] ),
    .QN(_0461_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0124_),
    .CK(net4),
    .Q(\mem[7][5] ),
    .QN(_0460_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0125_),
    .CK(net4),
    .Q(\mem[7][6] ),
    .QN(_0459_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0126_),
    .CK(net4),
    .Q(\mem[7][7] ),
    .QN(_0458_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0127_),
    .CK(net4),
    .Q(\mem[8][0] ),
    .QN(_0457_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0128_),
    .CK(net4),
    .Q(\mem[8][1] ),
    .QN(_0456_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0129_),
    .CK(net4),
    .Q(\mem[8][2] ),
    .QN(_0455_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0130_),
    .CK(net4),
    .Q(\mem[8][3] ),
    .QN(_0454_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0131_),
    .CK(net4),
    .Q(\mem[8][4] ),
    .QN(_0453_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0132_),
    .CK(net4),
    .Q(\mem[8][5] ),
    .QN(_0452_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0133_),
    .CK(net4),
    .Q(\mem[8][6] ),
    .QN(_0451_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0134_),
    .CK(net4),
    .Q(\mem[8][7] ),
    .QN(_0450_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0135_),
    .CK(net4),
    .Q(\mem[9][0] ),
    .QN(_0449_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0136_),
    .CK(net4),
    .Q(\mem[9][1] ),
    .QN(_0448_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0137_),
    .CK(net4),
    .Q(\mem[9][2] ),
    .QN(_0447_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0138_),
    .CK(net4),
    .Q(\mem[9][3] ),
    .QN(_0446_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0139_),
    .CK(net4),
    .Q(\mem[9][4] ),
    .QN(_0445_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0140_),
    .CK(net4),
    .Q(\mem[9][5] ),
    .QN(_0444_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0141_),
    .CK(net4),
    .Q(\mem[9][6] ),
    .QN(_0443_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0142_),
    .CK(net4),
    .Q(\mem[9][7] ),
    .QN(_0572_));
 DFFR_X1 \pointer_wraparound_error$_DFF_PN0_  (.D(_0010_),
    .RN(net6),
    .CK(net4),
    .Q(net11),
    .QN(_0442_));
 DFFR_X1 \rd_data_reg[0]$_DFFE_PN0P_  (.D(_0143_),
    .RN(net3),
    .CK(net1),
    .Q(net17),
    .QN(_0441_));
 DFFR_X1 \rd_data_reg[1]$_DFFE_PN0P_  (.D(_0144_),
    .RN(net3),
    .CK(net1),
    .Q(net18),
    .QN(_0440_));
 DFFR_X1 \rd_data_reg[2]$_DFFE_PN0P_  (.D(_0145_),
    .RN(net3),
    .CK(net1),
    .Q(net19),
    .QN(_0439_));
 DFFR_X1 \rd_data_reg[3]$_DFFE_PN0P_  (.D(_0146_),
    .RN(net3),
    .CK(net1),
    .Q(net20),
    .QN(_0438_));
 DFFR_X1 \rd_data_reg[4]$_DFFE_PN0P_  (.D(_0147_),
    .RN(net3),
    .CK(net1),
    .Q(net21),
    .QN(_0437_));
 DFFR_X1 \rd_data_reg[5]$_DFFE_PN0P_  (.D(_0148_),
    .RN(net3),
    .CK(net1),
    .Q(net22),
    .QN(_0436_));
 DFFR_X1 \rd_data_reg[6]$_DFFE_PN0P_  (.D(_0149_),
    .RN(net3),
    .CK(net1),
    .Q(net23),
    .QN(_0435_));
 DFFR_X1 \rd_data_reg[7]$_DFFE_PN0P_  (.D(_0150_),
    .RN(net3),
    .CK(net1),
    .Q(net24),
    .QN(_0434_));
 DFFR_X2 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_0151_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[0] ),
    .QN(_0013_));
 DFFR_X2 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_0152_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[1] ),
    .QN(_0595_));
 DFFR_X2 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_0153_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[2] ),
    .QN(_0611_));
 DFFR_X2 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_0154_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[3] ),
    .QN(_0601_));
 DFFR_X1 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_0155_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[0] ),
    .QN(_0433_));
 DFFR_X1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_0156_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[1] ),
    .QN(_0432_));
 DFFR_X1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_0157_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[2] ),
    .QN(_0431_));
 DFFR_X1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_0158_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[3] ),
    .QN(_0430_));
 DFFR_X2 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_0159_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[4] ),
    .QN(_0573_));
 DFFR_X1 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[0] ),
    .QN(_0574_));
 DFFR_X1 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[1] ),
    .QN(_0575_));
 DFFR_X1 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[2] ),
    .QN(_0576_));
 DFFR_X1 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[3] ),
    .QN(_0577_));
 DFFR_X1 \rd_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[4] ),
    .QN(_0578_));
 DFFR_X1 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[0] ),
    .QN(_0579_));
 DFFR_X1 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[1] ),
    .QN(_0580_));
 DFFR_X1 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[2] ),
    .QN(_0581_));
 DFFR_X1 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[3] ),
    .QN(_0582_));
 DFFR_X1 \rd_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[4] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[4] ),
    .QN(_0583_));
 DFFR_X1 \rd_ptr_sync[0]$_DFF_PN0_  (.D(_0006_),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_sync[0] ),
    .QN(_0621_));
 DFFR_X1 \rd_ptr_sync[1]$_DFF_PN0_  (.D(_0007_),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_sync[1] ),
    .QN(_0598_));
 DFFR_X1 \rd_ptr_sync[2]$_DFF_PN0_  (.D(_0008_),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_sync[2] ),
    .QN(_0628_));
 DFFR_X1 \rd_ptr_sync[3]$_DFF_PN0_  (.D(_0009_),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_sync[3] ),
    .QN(_0632_));
 DFFR_X1 \rd_ptr_sync[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync2[4] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_sync[4] ),
    .QN(_0584_));
 DFFR_X1 \sync_error$_DFF_PN0_  (.D(net31),
    .RN(net3),
    .CK(net1),
    .Q(net25),
    .QN(_0429_));
 DFFR_X2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_0160_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[0] ),
    .QN(_0011_));
 DFFR_X2 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_0161_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[1] ),
    .QN(_0627_));
 DFFR_X1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_0162_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[2] ),
    .QN(_0631_));
 DFFR_X1 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_0163_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[3] ),
    .QN(_0635_));
 DFFR_X1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_0164_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[0] ),
    .QN(_0428_));
 DFFR_X1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_0165_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[1] ),
    .QN(_0427_));
 DFFR_X1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_0166_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[2] ),
    .QN(_0426_));
 DFFR_X1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_0167_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[3] ),
    .QN(_0425_));
 DFFR_X2 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_0168_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[4] ),
    .QN(_0636_));
 DFFR_X1 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[0] ),
    .QN(_0585_));
 DFFR_X1 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[1] ),
    .QN(_0586_));
 DFFR_X1 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[2] ),
    .QN(_0587_));
 DFFR_X1 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[3] ),
    .QN(_0588_));
 DFFR_X1 \wr_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[4] ),
    .QN(_0589_));
 DFFR_X1 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[0] ),
    .QN(_0590_));
 DFFR_X1 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[1] ),
    .QN(_0591_));
 DFFR_X1 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[2] ),
    .QN(_0592_));
 DFFR_X1 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[3] ),
    .QN(_0593_));
 DFFR_X1 \wr_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[4] ),
    .QN(_0594_));
 DFFR_X1 \wr_ptr_sync[0]$_DFF_PN0_  (.D(_0002_),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_sync[0] ),
    .QN(_0617_));
 DFFR_X1 \wr_ptr_sync[1]$_DFF_PN0_  (.D(_0003_),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_sync[1] ),
    .QN(_0610_));
 DFFR_X1 \wr_ptr_sync[2]$_DFF_PN0_  (.D(_0004_),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_sync[2] ),
    .QN(_0614_));
 DFFR_X1 \wr_ptr_sync[3]$_DFF_PN0_  (.D(_0005_),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_sync[3] ),
    .QN(_0604_));
 DFFR_X1 \wr_ptr_sync[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync2[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_sync[4] ),
    .QN(_0605_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_75 ();
 BUF_X4 input1 (.A(rd_clk),
    .Z(net1));
 BUF_X1 input2 (.A(rd_en),
    .Z(net2));
 BUF_X8 input3 (.A(rd_rst_n),
    .Z(net3));
 BUF_X32 input4 (.A(wr_clk),
    .Z(net4));
 BUF_X1 input5 (.A(wr_en),
    .Z(net5));
 BUF_X8 input6 (.A(wr_rst_n),
    .Z(net6));
 BUF_X1 output7 (.A(net7),
    .Z(almost_empty));
 BUF_X1 output8 (.A(net8),
    .Z(almost_full));
 BUF_X1 output9 (.A(net9),
    .Z(empty));
 BUF_X1 output10 (.A(net10),
    .Z(full));
 BUF_X1 output11 (.A(net11),
    .Z(pointer_wraparound_flag));
 BUF_X1 output12 (.A(net12),
    .Z(rd_count[0]));
 BUF_X1 output13 (.A(net13),
    .Z(rd_count[1]));
 BUF_X1 output14 (.A(net14),
    .Z(rd_count[2]));
 BUF_X1 output15 (.A(net15),
    .Z(rd_count[3]));
 BUF_X1 output16 (.A(net16),
    .Z(rd_count[4]));
 BUF_X1 output17 (.A(net17),
    .Z(rd_data[0]));
 BUF_X1 output18 (.A(net18),
    .Z(rd_data[1]));
 BUF_X1 output19 (.A(net19),
    .Z(rd_data[2]));
 BUF_X1 output20 (.A(net20),
    .Z(rd_data[3]));
 BUF_X1 output21 (.A(net21),
    .Z(rd_data[4]));
 BUF_X1 output22 (.A(net22),
    .Z(rd_data[5]));
 BUF_X1 output23 (.A(net23),
    .Z(rd_data[6]));
 BUF_X1 output24 (.A(net24),
    .Z(rd_data[7]));
 BUF_X1 output25 (.A(net25),
    .Z(sync_error_flag));
 BUF_X1 output26 (.A(net26),
    .Z(wr_count[0]));
 BUF_X1 output27 (.A(net27),
    .Z(wr_count[1]));
 BUF_X1 output28 (.A(net28),
    .Z(wr_count[2]));
 BUF_X1 output29 (.A(net29),
    .Z(wr_count[3]));
 BUF_X1 output30 (.A(net30),
    .Z(wr_count[4]));
 LOGIC1_X1 \sync_error$_DFF_PN0__31  (.Z(net31));
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_90 ();
 FILLCELL_X2 FILLER_0_122 ();
 FILLCELL_X32 FILLER_0_141 ();
 FILLCELL_X2 FILLER_0_173 ();
 FILLCELL_X8 FILLER_0_192 ();
 FILLCELL_X4 FILLER_0_200 ();
 FILLCELL_X2 FILLER_0_204 ();
 FILLCELL_X1 FILLER_0_206 ();
 FILLCELL_X16 FILLER_0_212 ();
 FILLCELL_X8 FILLER_0_228 ();
 FILLCELL_X4 FILLER_0_236 ();
 FILLCELL_X1 FILLER_0_269 ();
 FILLCELL_X8 FILLER_0_273 ();
 FILLCELL_X1 FILLER_0_281 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X1 FILLER_1_41 ();
 FILLCELL_X4 FILLER_1_90 ();
 FILLCELL_X2 FILLER_1_94 ();
 FILLCELL_X2 FILLER_1_103 ();
 FILLCELL_X4 FILLER_1_122 ();
 FILLCELL_X2 FILLER_1_126 ();
 FILLCELL_X8 FILLER_1_145 ();
 FILLCELL_X1 FILLER_1_153 ();
 FILLCELL_X2 FILLER_1_171 ();
 FILLCELL_X1 FILLER_1_173 ();
 FILLCELL_X4 FILLER_1_191 ();
 FILLCELL_X4 FILLER_1_234 ();
 FILLCELL_X2 FILLER_1_238 ();
 FILLCELL_X1 FILLER_1_240 ();
 FILLCELL_X1 FILLER_1_265 ();
 FILLCELL_X4 FILLER_1_276 ();
 FILLCELL_X2 FILLER_1_280 ();
 FILLCELL_X4 FILLER_2_1 ();
 FILLCELL_X2 FILLER_2_5 ();
 FILLCELL_X1 FILLER_2_41 ();
 FILLCELL_X16 FILLER_2_66 ();
 FILLCELL_X2 FILLER_2_120 ();
 FILLCELL_X2 FILLER_2_136 ();
 FILLCELL_X1 FILLER_2_145 ();
 FILLCELL_X2 FILLER_2_163 ();
 FILLCELL_X2 FILLER_2_172 ();
 FILLCELL_X8 FILLER_2_188 ();
 FILLCELL_X16 FILLER_2_223 ();
 FILLCELL_X2 FILLER_2_239 ();
 FILLCELL_X1 FILLER_2_241 ();
 FILLCELL_X1 FILLER_2_262 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X4 FILLER_3_17 ();
 FILLCELL_X4 FILLER_3_42 ();
 FILLCELL_X1 FILLER_3_46 ();
 FILLCELL_X1 FILLER_3_54 ();
 FILLCELL_X16 FILLER_3_93 ();
 FILLCELL_X1 FILLER_3_109 ();
 FILLCELL_X4 FILLER_3_117 ();
 FILLCELL_X8 FILLER_3_145 ();
 FILLCELL_X4 FILLER_3_153 ();
 FILLCELL_X1 FILLER_3_157 ();
 FILLCELL_X2 FILLER_3_172 ();
 FILLCELL_X1 FILLER_3_174 ();
 FILLCELL_X8 FILLER_3_182 ();
 FILLCELL_X4 FILLER_3_190 ();
 FILLCELL_X4 FILLER_3_200 ();
 FILLCELL_X1 FILLER_3_204 ();
 FILLCELL_X4 FILLER_3_236 ();
 FILLCELL_X1 FILLER_3_240 ();
 FILLCELL_X4 FILLER_3_243 ();
 FILLCELL_X2 FILLER_3_268 ();
 FILLCELL_X1 FILLER_3_270 ();
 FILLCELL_X4 FILLER_3_273 ();
 FILLCELL_X1 FILLER_3_277 ();
 FILLCELL_X2 FILLER_3_280 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X4 FILLER_4_17 ();
 FILLCELL_X16 FILLER_4_45 ();
 FILLCELL_X4 FILLER_4_61 ();
 FILLCELL_X1 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_90 ();
 FILLCELL_X2 FILLER_4_122 ();
 FILLCELL_X1 FILLER_4_124 ();
 FILLCELL_X32 FILLER_4_142 ();
 FILLCELL_X1 FILLER_4_174 ();
 FILLCELL_X16 FILLER_4_182 ();
 FILLCELL_X4 FILLER_4_198 ();
 FILLCELL_X2 FILLER_4_202 ();
 FILLCELL_X2 FILLER_4_209 ();
 FILLCELL_X1 FILLER_4_211 ();
 FILLCELL_X16 FILLER_4_219 ();
 FILLCELL_X4 FILLER_4_235 ();
 FILLCELL_X2 FILLER_4_239 ();
 FILLCELL_X4 FILLER_4_251 ();
 FILLCELL_X2 FILLER_4_265 ();
 FILLCELL_X1 FILLER_4_267 ();
 FILLCELL_X1 FILLER_4_281 ();
 FILLCELL_X8 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_9 ();
 FILLCELL_X2 FILLER_5_13 ();
 FILLCELL_X16 FILLER_5_46 ();
 FILLCELL_X8 FILLER_5_62 ();
 FILLCELL_X4 FILLER_5_70 ();
 FILLCELL_X2 FILLER_5_74 ();
 FILLCELL_X1 FILLER_5_76 ();
 FILLCELL_X4 FILLER_5_84 ();
 FILLCELL_X16 FILLER_5_95 ();
 FILLCELL_X4 FILLER_5_111 ();
 FILLCELL_X2 FILLER_5_115 ();
 FILLCELL_X4 FILLER_5_120 ();
 FILLCELL_X2 FILLER_5_124 ();
 FILLCELL_X4 FILLER_5_140 ();
 FILLCELL_X1 FILLER_5_144 ();
 FILLCELL_X8 FILLER_5_152 ();
 FILLCELL_X2 FILLER_5_160 ();
 FILLCELL_X4 FILLER_5_182 ();
 FILLCELL_X1 FILLER_5_186 ();
 FILLCELL_X2 FILLER_5_201 ();
 FILLCELL_X1 FILLER_5_203 ();
 FILLCELL_X2 FILLER_5_214 ();
 FILLCELL_X1 FILLER_5_216 ();
 FILLCELL_X2 FILLER_5_279 ();
 FILLCELL_X1 FILLER_5_281 ();
 FILLCELL_X16 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_17 ();
 FILLCELL_X2 FILLER_6_21 ();
 FILLCELL_X1 FILLER_6_23 ();
 FILLCELL_X8 FILLER_6_31 ();
 FILLCELL_X4 FILLER_6_39 ();
 FILLCELL_X1 FILLER_6_43 ();
 FILLCELL_X16 FILLER_6_61 ();
 FILLCELL_X4 FILLER_6_77 ();
 FILLCELL_X8 FILLER_6_88 ();
 FILLCELL_X2 FILLER_6_113 ();
 FILLCELL_X1 FILLER_6_115 ();
 FILLCELL_X4 FILLER_6_119 ();
 FILLCELL_X2 FILLER_6_123 ();
 FILLCELL_X8 FILLER_6_145 ();
 FILLCELL_X2 FILLER_6_153 ();
 FILLCELL_X1 FILLER_6_155 ();
 FILLCELL_X4 FILLER_6_163 ();
 FILLCELL_X1 FILLER_6_167 ();
 FILLCELL_X1 FILLER_6_185 ();
 FILLCELL_X16 FILLER_6_224 ();
 FILLCELL_X4 FILLER_6_240 ();
 FILLCELL_X2 FILLER_6_244 ();
 FILLCELL_X1 FILLER_6_246 ();
 FILLCELL_X2 FILLER_6_253 ();
 FILLCELL_X4 FILLER_6_275 ();
 FILLCELL_X2 FILLER_6_279 ();
 FILLCELL_X1 FILLER_6_281 ();
 FILLCELL_X8 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_9 ();
 FILLCELL_X4 FILLER_7_49 ();
 FILLCELL_X4 FILLER_7_60 ();
 FILLCELL_X2 FILLER_7_71 ();
 FILLCELL_X1 FILLER_7_73 ();
 FILLCELL_X4 FILLER_7_91 ();
 FILLCELL_X2 FILLER_7_95 ();
 FILLCELL_X4 FILLER_7_104 ();
 FILLCELL_X2 FILLER_7_108 ();
 FILLCELL_X8 FILLER_7_117 ();
 FILLCELL_X1 FILLER_7_125 ();
 FILLCELL_X2 FILLER_7_150 ();
 FILLCELL_X1 FILLER_7_152 ();
 FILLCELL_X2 FILLER_7_156 ();
 FILLCELL_X2 FILLER_7_167 ();
 FILLCELL_X1 FILLER_7_189 ();
 FILLCELL_X4 FILLER_7_213 ();
 FILLCELL_X8 FILLER_7_237 ();
 FILLCELL_X4 FILLER_7_245 ();
 FILLCELL_X2 FILLER_7_249 ();
 FILLCELL_X1 FILLER_7_251 ();
 FILLCELL_X4 FILLER_7_277 ();
 FILLCELL_X1 FILLER_7_281 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_17 ();
 FILLCELL_X2 FILLER_8_25 ();
 FILLCELL_X4 FILLER_8_44 ();
 FILLCELL_X2 FILLER_8_48 ();
 FILLCELL_X8 FILLER_8_67 ();
 FILLCELL_X2 FILLER_8_82 ();
 FILLCELL_X1 FILLER_8_91 ();
 FILLCELL_X1 FILLER_8_116 ();
 FILLCELL_X8 FILLER_8_124 ();
 FILLCELL_X4 FILLER_8_132 ();
 FILLCELL_X1 FILLER_8_136 ();
 FILLCELL_X4 FILLER_8_151 ();
 FILLCELL_X2 FILLER_8_155 ();
 FILLCELL_X1 FILLER_8_157 ();
 FILLCELL_X2 FILLER_8_188 ();
 FILLCELL_X1 FILLER_8_209 ();
 FILLCELL_X8 FILLER_8_222 ();
 FILLCELL_X4 FILLER_8_250 ();
 FILLCELL_X2 FILLER_8_254 ();
 FILLCELL_X16 FILLER_8_265 ();
 FILLCELL_X1 FILLER_8_281 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X4 FILLER_9_25 ();
 FILLCELL_X1 FILLER_9_29 ();
 FILLCELL_X16 FILLER_9_47 ();
 FILLCELL_X4 FILLER_9_63 ();
 FILLCELL_X1 FILLER_9_67 ();
 FILLCELL_X16 FILLER_9_92 ();
 FILLCELL_X8 FILLER_9_108 ();
 FILLCELL_X4 FILLER_9_116 ();
 FILLCELL_X2 FILLER_9_120 ();
 FILLCELL_X1 FILLER_9_122 ();
 FILLCELL_X2 FILLER_9_126 ();
 FILLCELL_X8 FILLER_9_135 ();
 FILLCELL_X2 FILLER_9_143 ();
 FILLCELL_X1 FILLER_9_163 ();
 FILLCELL_X4 FILLER_9_174 ();
 FILLCELL_X2 FILLER_9_187 ();
 FILLCELL_X1 FILLER_9_215 ();
 FILLCELL_X32 FILLER_9_222 ();
 FILLCELL_X4 FILLER_9_254 ();
 FILLCELL_X2 FILLER_9_258 ();
 FILLCELL_X2 FILLER_9_280 ();
 FILLCELL_X2 FILLER_10_25 ();
 FILLCELL_X1 FILLER_10_27 ();
 FILLCELL_X4 FILLER_10_42 ();
 FILLCELL_X2 FILLER_10_46 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X8 FILLER_10_97 ();
 FILLCELL_X4 FILLER_10_105 ();
 FILLCELL_X2 FILLER_10_109 ();
 FILLCELL_X1 FILLER_10_111 ();
 FILLCELL_X4 FILLER_10_115 ();
 FILLCELL_X2 FILLER_10_119 ();
 FILLCELL_X1 FILLER_10_121 ();
 FILLCELL_X2 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_150 ();
 FILLCELL_X2 FILLER_10_160 ();
 FILLCELL_X2 FILLER_10_175 ();
 FILLCELL_X2 FILLER_10_190 ();
 FILLCELL_X1 FILLER_10_192 ();
 FILLCELL_X2 FILLER_10_214 ();
 FILLCELL_X1 FILLER_10_216 ();
 FILLCELL_X8 FILLER_10_237 ();
 FILLCELL_X4 FILLER_10_245 ();
 FILLCELL_X4 FILLER_10_272 ();
 FILLCELL_X2 FILLER_10_276 ();
 FILLCELL_X1 FILLER_10_278 ();
 FILLCELL_X2 FILLER_11_42 ();
 FILLCELL_X1 FILLER_11_44 ();
 FILLCELL_X32 FILLER_11_76 ();
 FILLCELL_X2 FILLER_11_108 ();
 FILLCELL_X1 FILLER_11_110 ();
 FILLCELL_X2 FILLER_11_135 ();
 FILLCELL_X8 FILLER_11_233 ();
 FILLCELL_X1 FILLER_11_241 ();
 FILLCELL_X8 FILLER_11_271 ();
 FILLCELL_X2 FILLER_11_279 ();
 FILLCELL_X1 FILLER_11_281 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_17 ();
 FILLCELL_X1 FILLER_12_25 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X4 FILLER_12_49 ();
 FILLCELL_X4 FILLER_12_67 ();
 FILLCELL_X1 FILLER_12_71 ();
 FILLCELL_X2 FILLER_12_79 ();
 FILLCELL_X2 FILLER_12_88 ();
 FILLCELL_X1 FILLER_12_90 ();
 FILLCELL_X8 FILLER_12_108 ();
 FILLCELL_X4 FILLER_12_116 ();
 FILLCELL_X1 FILLER_12_120 ();
 FILLCELL_X1 FILLER_12_135 ();
 FILLCELL_X16 FILLER_12_143 ();
 FILLCELL_X4 FILLER_12_159 ();
 FILLCELL_X2 FILLER_12_163 ();
 FILLCELL_X8 FILLER_12_169 ();
 FILLCELL_X2 FILLER_12_177 ();
 FILLCELL_X4 FILLER_12_192 ();
 FILLCELL_X1 FILLER_12_208 ();
 FILLCELL_X1 FILLER_12_215 ();
 FILLCELL_X1 FILLER_12_245 ();
 FILLCELL_X4 FILLER_12_256 ();
 FILLCELL_X2 FILLER_12_280 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_9 ();
 FILLCELL_X4 FILLER_13_35 ();
 FILLCELL_X2 FILLER_13_46 ();
 FILLCELL_X1 FILLER_13_48 ();
 FILLCELL_X8 FILLER_13_66 ();
 FILLCELL_X8 FILLER_13_98 ();
 FILLCELL_X4 FILLER_13_106 ();
 FILLCELL_X8 FILLER_13_134 ();
 FILLCELL_X2 FILLER_13_142 ();
 FILLCELL_X8 FILLER_13_161 ();
 FILLCELL_X2 FILLER_13_169 ();
 FILLCELL_X1 FILLER_13_178 ();
 FILLCELL_X8 FILLER_13_195 ();
 FILLCELL_X2 FILLER_13_203 ();
 FILLCELL_X16 FILLER_13_239 ();
 FILLCELL_X8 FILLER_13_255 ();
 FILLCELL_X4 FILLER_13_263 ();
 FILLCELL_X4 FILLER_13_276 ();
 FILLCELL_X2 FILLER_13_280 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X2 FILLER_14_25 ();
 FILLCELL_X1 FILLER_14_34 ();
 FILLCELL_X16 FILLER_14_59 ();
 FILLCELL_X8 FILLER_14_75 ();
 FILLCELL_X2 FILLER_14_83 ();
 FILLCELL_X16 FILLER_14_109 ();
 FILLCELL_X8 FILLER_14_125 ();
 FILLCELL_X4 FILLER_14_140 ();
 FILLCELL_X8 FILLER_14_158 ();
 FILLCELL_X4 FILLER_14_166 ();
 FILLCELL_X4 FILLER_14_204 ();
 FILLCELL_X4 FILLER_14_228 ();
 FILLCELL_X1 FILLER_14_232 ();
 FILLCELL_X8 FILLER_14_253 ();
 FILLCELL_X1 FILLER_14_261 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_21 ();
 FILLCELL_X16 FILLER_15_29 ();
 FILLCELL_X4 FILLER_15_45 ();
 FILLCELL_X1 FILLER_15_49 ();
 FILLCELL_X2 FILLER_15_57 ();
 FILLCELL_X16 FILLER_15_76 ();
 FILLCELL_X2 FILLER_15_92 ();
 FILLCELL_X2 FILLER_15_101 ();
 FILLCELL_X1 FILLER_15_103 ();
 FILLCELL_X8 FILLER_15_121 ();
 FILLCELL_X2 FILLER_15_129 ();
 FILLCELL_X1 FILLER_15_131 ();
 FILLCELL_X1 FILLER_15_146 ();
 FILLCELL_X16 FILLER_15_164 ();
 FILLCELL_X8 FILLER_15_194 ();
 FILLCELL_X32 FILLER_15_222 ();
 FILLCELL_X8 FILLER_15_254 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X1 FILLER_16_9 ();
 FILLCELL_X16 FILLER_16_14 ();
 FILLCELL_X2 FILLER_16_30 ();
 FILLCELL_X2 FILLER_16_36 ();
 FILLCELL_X2 FILLER_16_55 ();
 FILLCELL_X1 FILLER_16_57 ();
 FILLCELL_X4 FILLER_16_65 ();
 FILLCELL_X2 FILLER_16_69 ();
 FILLCELL_X16 FILLER_16_78 ();
 FILLCELL_X2 FILLER_16_94 ();
 FILLCELL_X1 FILLER_16_120 ();
 FILLCELL_X2 FILLER_16_172 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X1 FILLER_16_225 ();
 FILLCELL_X16 FILLER_16_266 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_5 ();
 FILLCELL_X1 FILLER_17_7 ();
 FILLCELL_X8 FILLER_17_32 ();
 FILLCELL_X1 FILLER_17_40 ();
 FILLCELL_X4 FILLER_17_55 ();
 FILLCELL_X2 FILLER_17_59 ();
 FILLCELL_X4 FILLER_17_85 ();
 FILLCELL_X1 FILLER_17_89 ();
 FILLCELL_X4 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_157 ();
 FILLCELL_X2 FILLER_17_172 ();
 FILLCELL_X2 FILLER_17_188 ();
 FILLCELL_X1 FILLER_17_190 ();
 FILLCELL_X4 FILLER_17_198 ();
 FILLCELL_X2 FILLER_17_202 ();
 FILLCELL_X1 FILLER_17_204 ();
 FILLCELL_X32 FILLER_17_212 ();
 FILLCELL_X4 FILLER_17_244 ();
 FILLCELL_X1 FILLER_17_248 ();
 FILLCELL_X8 FILLER_17_269 ();
 FILLCELL_X4 FILLER_17_277 ();
 FILLCELL_X1 FILLER_17_281 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_3 ();
 FILLCELL_X4 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_32 ();
 FILLCELL_X4 FILLER_18_50 ();
 FILLCELL_X2 FILLER_18_54 ();
 FILLCELL_X2 FILLER_18_63 ();
 FILLCELL_X32 FILLER_18_72 ();
 FILLCELL_X4 FILLER_18_104 ();
 FILLCELL_X2 FILLER_18_108 ();
 FILLCELL_X1 FILLER_18_110 ();
 FILLCELL_X8 FILLER_18_125 ();
 FILLCELL_X2 FILLER_18_133 ();
 FILLCELL_X1 FILLER_18_135 ();
 FILLCELL_X8 FILLER_18_141 ();
 FILLCELL_X4 FILLER_18_149 ();
 FILLCELL_X1 FILLER_18_153 ();
 FILLCELL_X2 FILLER_18_171 ();
 FILLCELL_X2 FILLER_18_180 ();
 FILLCELL_X1 FILLER_18_182 ();
 FILLCELL_X1 FILLER_18_200 ();
 FILLCELL_X1 FILLER_18_221 ();
 FILLCELL_X8 FILLER_18_242 ();
 FILLCELL_X2 FILLER_18_250 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X1 FILLER_19_13 ();
 FILLCELL_X4 FILLER_19_35 ();
 FILLCELL_X8 FILLER_19_46 ();
 FILLCELL_X4 FILLER_19_54 ();
 FILLCELL_X2 FILLER_19_58 ();
 FILLCELL_X1 FILLER_19_72 ();
 FILLCELL_X8 FILLER_19_78 ();
 FILLCELL_X2 FILLER_19_86 ();
 FILLCELL_X1 FILLER_19_88 ();
 FILLCELL_X16 FILLER_19_96 ();
 FILLCELL_X2 FILLER_19_112 ();
 FILLCELL_X1 FILLER_19_128 ();
 FILLCELL_X8 FILLER_19_134 ();
 FILLCELL_X1 FILLER_19_142 ();
 FILLCELL_X32 FILLER_19_150 ();
 FILLCELL_X16 FILLER_19_182 ();
 FILLCELL_X4 FILLER_19_198 ();
 FILLCELL_X4 FILLER_19_209 ();
 FILLCELL_X2 FILLER_19_213 ();
 FILLCELL_X8 FILLER_19_242 ();
 FILLCELL_X2 FILLER_19_250 ();
 FILLCELL_X4 FILLER_19_272 ();
 FILLCELL_X2 FILLER_19_276 ();
 FILLCELL_X1 FILLER_19_278 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_5 ();
 FILLCELL_X1 FILLER_20_7 ();
 FILLCELL_X8 FILLER_20_12 ();
 FILLCELL_X1 FILLER_20_20 ();
 FILLCELL_X1 FILLER_20_38 ();
 FILLCELL_X4 FILLER_20_56 ();
 FILLCELL_X2 FILLER_20_88 ();
 FILLCELL_X4 FILLER_20_107 ();
 FILLCELL_X1 FILLER_20_111 ();
 FILLCELL_X8 FILLER_20_125 ();
 FILLCELL_X2 FILLER_20_133 ();
 FILLCELL_X1 FILLER_20_135 ();
 FILLCELL_X2 FILLER_20_143 ();
 FILLCELL_X4 FILLER_20_162 ();
 FILLCELL_X2 FILLER_20_166 ();
 FILLCELL_X1 FILLER_20_168 ();
 FILLCELL_X16 FILLER_20_176 ();
 FILLCELL_X2 FILLER_20_192 ();
 FILLCELL_X1 FILLER_20_194 ();
 FILLCELL_X16 FILLER_20_204 ();
 FILLCELL_X2 FILLER_20_220 ();
 FILLCELL_X16 FILLER_20_229 ();
 FILLCELL_X4 FILLER_20_245 ();
 FILLCELL_X2 FILLER_20_249 ();
 FILLCELL_X1 FILLER_20_251 ();
 FILLCELL_X1 FILLER_20_278 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_26 ();
 FILLCELL_X2 FILLER_21_34 ();
 FILLCELL_X4 FILLER_21_43 ();
 FILLCELL_X2 FILLER_21_47 ();
 FILLCELL_X4 FILLER_21_63 ();
 FILLCELL_X8 FILLER_21_98 ();
 FILLCELL_X2 FILLER_21_106 ();
 FILLCELL_X1 FILLER_21_108 ();
 FILLCELL_X4 FILLER_21_116 ();
 FILLCELL_X2 FILLER_21_120 ();
 FILLCELL_X2 FILLER_21_134 ();
 FILLCELL_X1 FILLER_21_136 ();
 FILLCELL_X2 FILLER_21_154 ();
 FILLCELL_X1 FILLER_21_156 ();
 FILLCELL_X4 FILLER_21_164 ();
 FILLCELL_X2 FILLER_21_168 ();
 FILLCELL_X4 FILLER_21_187 ();
 FILLCELL_X2 FILLER_21_191 ();
 FILLCELL_X4 FILLER_21_197 ();
 FILLCELL_X2 FILLER_21_201 ();
 FILLCELL_X1 FILLER_21_203 ();
 FILLCELL_X16 FILLER_21_210 ();
 FILLCELL_X2 FILLER_21_226 ();
 FILLCELL_X8 FILLER_21_248 ();
 FILLCELL_X2 FILLER_21_256 ();
 FILLCELL_X1 FILLER_21_258 ();
 FILLCELL_X4 FILLER_21_263 ();
 FILLCELL_X2 FILLER_21_267 ();
 FILLCELL_X4 FILLER_21_278 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_33 ();
 FILLCELL_X16 FILLER_22_54 ();
 FILLCELL_X16 FILLER_22_77 ();
 FILLCELL_X8 FILLER_22_93 ();
 FILLCELL_X2 FILLER_22_101 ();
 FILLCELL_X1 FILLER_22_135 ();
 FILLCELL_X4 FILLER_22_138 ();
 FILLCELL_X4 FILLER_22_149 ();
 FILLCELL_X2 FILLER_22_153 ();
 FILLCELL_X1 FILLER_22_155 ();
 FILLCELL_X8 FILLER_22_180 ();
 FILLCELL_X2 FILLER_22_188 ();
 FILLCELL_X4 FILLER_22_218 ();
 FILLCELL_X2 FILLER_22_222 ();
 FILLCELL_X1 FILLER_22_224 ();
 FILLCELL_X16 FILLER_22_252 ();
 FILLCELL_X1 FILLER_22_268 ();
 FILLCELL_X2 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_3 ();
 FILLCELL_X8 FILLER_23_28 ();
 FILLCELL_X4 FILLER_23_36 ();
 FILLCELL_X1 FILLER_23_40 ();
 FILLCELL_X16 FILLER_23_48 ();
 FILLCELL_X4 FILLER_23_64 ();
 FILLCELL_X1 FILLER_23_68 ();
 FILLCELL_X32 FILLER_23_74 ();
 FILLCELL_X4 FILLER_23_106 ();
 FILLCELL_X2 FILLER_23_110 ();
 FILLCELL_X1 FILLER_23_112 ();
 FILLCELL_X2 FILLER_23_123 ();
 FILLCELL_X16 FILLER_23_131 ();
 FILLCELL_X8 FILLER_23_147 ();
 FILLCELL_X4 FILLER_23_155 ();
 FILLCELL_X2 FILLER_23_159 ();
 FILLCELL_X1 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_169 ();
 FILLCELL_X4 FILLER_23_177 ();
 FILLCELL_X2 FILLER_23_185 ();
 FILLCELL_X1 FILLER_23_187 ();
 FILLCELL_X1 FILLER_23_195 ();
 FILLCELL_X4 FILLER_23_231 ();
 FILLCELL_X1 FILLER_23_235 ();
 FILLCELL_X2 FILLER_24_1 ();
 FILLCELL_X1 FILLER_24_3 ();
 FILLCELL_X2 FILLER_24_21 ();
 FILLCELL_X1 FILLER_24_23 ();
 FILLCELL_X8 FILLER_24_41 ();
 FILLCELL_X1 FILLER_24_49 ();
 FILLCELL_X8 FILLER_24_74 ();
 FILLCELL_X1 FILLER_24_82 ();
 FILLCELL_X2 FILLER_24_114 ();
 FILLCELL_X8 FILLER_24_140 ();
 FILLCELL_X4 FILLER_24_148 ();
 FILLCELL_X16 FILLER_24_169 ();
 FILLCELL_X2 FILLER_24_185 ();
 FILLCELL_X1 FILLER_24_187 ();
 FILLCELL_X2 FILLER_24_227 ();
 FILLCELL_X16 FILLER_24_249 ();
 FILLCELL_X8 FILLER_24_265 ();
 FILLCELL_X4 FILLER_24_273 ();
 FILLCELL_X2 FILLER_24_277 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_9 ();
 FILLCELL_X1 FILLER_25_18 ();
 FILLCELL_X4 FILLER_25_26 ();
 FILLCELL_X8 FILLER_25_44 ();
 FILLCELL_X1 FILLER_25_52 ();
 FILLCELL_X8 FILLER_25_71 ();
 FILLCELL_X1 FILLER_25_79 ();
 FILLCELL_X2 FILLER_25_104 ();
 FILLCELL_X1 FILLER_25_106 ();
 FILLCELL_X4 FILLER_25_114 ();
 FILLCELL_X1 FILLER_25_118 ();
 FILLCELL_X2 FILLER_25_126 ();
 FILLCELL_X4 FILLER_25_135 ();
 FILLCELL_X1 FILLER_25_139 ();
 FILLCELL_X8 FILLER_25_164 ();
 FILLCELL_X2 FILLER_25_172 ();
 FILLCELL_X8 FILLER_25_178 ();
 FILLCELL_X4 FILLER_25_186 ();
 FILLCELL_X2 FILLER_25_190 ();
 FILLCELL_X2 FILLER_25_196 ();
 FILLCELL_X1 FILLER_25_198 ();
 FILLCELL_X16 FILLER_25_227 ();
 FILLCELL_X4 FILLER_25_243 ();
 FILLCELL_X8 FILLER_25_267 ();
 FILLCELL_X4 FILLER_25_275 ();
 FILLCELL_X2 FILLER_25_279 ();
 FILLCELL_X1 FILLER_25_281 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_17 ();
 FILLCELL_X8 FILLER_26_43 ();
 FILLCELL_X2 FILLER_26_51 ();
 FILLCELL_X2 FILLER_26_77 ();
 FILLCELL_X4 FILLER_26_103 ();
 FILLCELL_X2 FILLER_26_107 ();
 FILLCELL_X1 FILLER_26_128 ();
 FILLCELL_X2 FILLER_26_146 ();
 FILLCELL_X2 FILLER_26_155 ();
 FILLCELL_X2 FILLER_26_164 ();
 FILLCELL_X1 FILLER_26_166 ();
 FILLCELL_X8 FILLER_26_198 ();
 FILLCELL_X4 FILLER_26_206 ();
 FILLCELL_X2 FILLER_26_210 ();
 FILLCELL_X1 FILLER_26_212 ();
 FILLCELL_X4 FILLER_26_244 ();
 FILLCELL_X1 FILLER_26_248 ();
 FILLCELL_X4 FILLER_26_278 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X8 FILLER_27_81 ();
 FILLCELL_X4 FILLER_27_89 ();
 FILLCELL_X8 FILLER_27_100 ();
 FILLCELL_X4 FILLER_27_108 ();
 FILLCELL_X2 FILLER_27_112 ();
 FILLCELL_X1 FILLER_27_114 ();
 FILLCELL_X16 FILLER_27_139 ();
 FILLCELL_X8 FILLER_27_155 ();
 FILLCELL_X1 FILLER_27_163 ();
 FILLCELL_X2 FILLER_27_186 ();
 FILLCELL_X1 FILLER_27_188 ();
 FILLCELL_X8 FILLER_27_194 ();
 FILLCELL_X4 FILLER_27_202 ();
 FILLCELL_X1 FILLER_27_206 ();
 FILLCELL_X8 FILLER_27_232 ();
 FILLCELL_X2 FILLER_27_240 ();
 FILLCELL_X1 FILLER_27_242 ();
 FILLCELL_X8 FILLER_27_252 ();
 FILLCELL_X4 FILLER_27_260 ();
 FILLCELL_X1 FILLER_27_264 ();
 FILLCELL_X4 FILLER_27_275 ();
 FILLCELL_X2 FILLER_27_279 ();
 FILLCELL_X1 FILLER_27_281 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_29 ();
 FILLCELL_X16 FILLER_28_61 ();
 FILLCELL_X2 FILLER_28_77 ();
 FILLCELL_X1 FILLER_28_79 ();
 FILLCELL_X32 FILLER_28_104 ();
 FILLCELL_X32 FILLER_28_136 ();
 FILLCELL_X4 FILLER_28_168 ();
 FILLCELL_X2 FILLER_28_172 ();
 FILLCELL_X1 FILLER_28_174 ();
 FILLCELL_X16 FILLER_28_188 ();
 FILLCELL_X8 FILLER_28_204 ();
 FILLCELL_X2 FILLER_28_212 ();
 FILLCELL_X1 FILLER_28_214 ();
 FILLCELL_X1 FILLER_28_227 ();
 FILLCELL_X4 FILLER_28_278 ();
 FILLCELL_X1 FILLER_29_18 ();
 FILLCELL_X2 FILLER_29_26 ();
 FILLCELL_X1 FILLER_29_28 ();
 FILLCELL_X4 FILLER_29_36 ();
 FILLCELL_X2 FILLER_29_40 ();
 FILLCELL_X2 FILLER_29_49 ();
 FILLCELL_X4 FILLER_29_75 ();
 FILLCELL_X4 FILLER_29_103 ();
 FILLCELL_X2 FILLER_29_107 ();
 FILLCELL_X8 FILLER_29_157 ();
 FILLCELL_X1 FILLER_29_165 ();
 FILLCELL_X16 FILLER_29_197 ();
 FILLCELL_X1 FILLER_29_213 ();
 FILLCELL_X8 FILLER_29_256 ();
 FILLCELL_X4 FILLER_29_264 ();
 FILLCELL_X1 FILLER_29_268 ();
 FILLCELL_X1 FILLER_29_281 ();
 FILLCELL_X2 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_3 ();
 FILLCELL_X1 FILLER_30_28 ();
 FILLCELL_X2 FILLER_30_77 ();
 FILLCELL_X1 FILLER_30_93 ();
 FILLCELL_X1 FILLER_30_101 ();
 FILLCELL_X1 FILLER_30_109 ();
 FILLCELL_X1 FILLER_30_134 ();
 FILLCELL_X4 FILLER_30_142 ();
 FILLCELL_X1 FILLER_30_146 ();
 FILLCELL_X8 FILLER_30_154 ();
 FILLCELL_X4 FILLER_30_162 ();
 FILLCELL_X2 FILLER_30_166 ();
 FILLCELL_X1 FILLER_30_168 ();
 FILLCELL_X8 FILLER_30_186 ();
 FILLCELL_X4 FILLER_30_194 ();
 FILLCELL_X2 FILLER_30_202 ();
 FILLCELL_X1 FILLER_30_204 ();
 FILLCELL_X32 FILLER_30_207 ();
 FILLCELL_X8 FILLER_30_239 ();
 FILLCELL_X4 FILLER_30_247 ();
 FILLCELL_X1 FILLER_30_251 ();
 FILLCELL_X1 FILLER_30_275 ();
 FILLCELL_X8 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_9 ();
 FILLCELL_X1 FILLER_31_18 ();
 FILLCELL_X2 FILLER_31_26 ();
 FILLCELL_X4 FILLER_31_35 ();
 FILLCELL_X4 FILLER_31_46 ();
 FILLCELL_X2 FILLER_31_50 ();
 FILLCELL_X1 FILLER_31_52 ();
 FILLCELL_X16 FILLER_31_96 ();
 FILLCELL_X8 FILLER_31_112 ();
 FILLCELL_X1 FILLER_31_120 ();
 FILLCELL_X2 FILLER_31_126 ();
 FILLCELL_X2 FILLER_31_134 ();
 FILLCELL_X1 FILLER_31_136 ();
 FILLCELL_X4 FILLER_31_159 ();
 FILLCELL_X2 FILLER_31_163 ();
 FILLCELL_X1 FILLER_31_165 ();
 FILLCELL_X2 FILLER_31_185 ();
 FILLCELL_X1 FILLER_31_187 ();
 FILLCELL_X2 FILLER_31_192 ();
 FILLCELL_X1 FILLER_31_194 ();
 FILLCELL_X16 FILLER_31_215 ();
 FILLCELL_X2 FILLER_31_231 ();
 FILLCELL_X8 FILLER_31_243 ();
 FILLCELL_X2 FILLER_31_251 ();
 FILLCELL_X1 FILLER_31_267 ();
 FILLCELL_X4 FILLER_32_1 ();
 FILLCELL_X2 FILLER_32_5 ();
 FILLCELL_X2 FILLER_32_18 ();
 FILLCELL_X16 FILLER_32_44 ();
 FILLCELL_X4 FILLER_32_60 ();
 FILLCELL_X2 FILLER_32_64 ();
 FILLCELL_X1 FILLER_32_66 ();
 FILLCELL_X16 FILLER_32_91 ();
 FILLCELL_X8 FILLER_32_107 ();
 FILLCELL_X1 FILLER_32_115 ();
 FILLCELL_X4 FILLER_32_121 ();
 FILLCELL_X1 FILLER_32_125 ();
 FILLCELL_X16 FILLER_32_132 ();
 FILLCELL_X2 FILLER_32_148 ();
 FILLCELL_X1 FILLER_32_150 ();
 FILLCELL_X4 FILLER_32_164 ();
 FILLCELL_X32 FILLER_32_175 ();
 FILLCELL_X8 FILLER_32_207 ();
 FILLCELL_X4 FILLER_32_215 ();
 FILLCELL_X4 FILLER_32_249 ();
 FILLCELL_X2 FILLER_32_253 ();
 FILLCELL_X1 FILLER_32_255 ();
 FILLCELL_X1 FILLER_32_278 ();
 FILLCELL_X2 FILLER_33_1 ();
 FILLCELL_X1 FILLER_33_3 ();
 FILLCELL_X8 FILLER_33_25 ();
 FILLCELL_X2 FILLER_33_33 ();
 FILLCELL_X8 FILLER_33_49 ();
 FILLCELL_X4 FILLER_33_57 ();
 FILLCELL_X2 FILLER_33_68 ();
 FILLCELL_X2 FILLER_33_84 ();
 FILLCELL_X1 FILLER_33_86 ();
 FILLCELL_X8 FILLER_33_94 ();
 FILLCELL_X4 FILLER_33_102 ();
 FILLCELL_X2 FILLER_33_106 ();
 FILLCELL_X1 FILLER_33_108 ();
 FILLCELL_X4 FILLER_33_116 ();
 FILLCELL_X4 FILLER_33_127 ();
 FILLCELL_X1 FILLER_33_131 ();
 FILLCELL_X2 FILLER_33_143 ();
 FILLCELL_X2 FILLER_33_166 ();
 FILLCELL_X16 FILLER_33_185 ();
 FILLCELL_X8 FILLER_33_201 ();
 FILLCELL_X2 FILLER_33_209 ();
 FILLCELL_X1 FILLER_33_211 ();
 FILLCELL_X8 FILLER_33_232 ();
 FILLCELL_X4 FILLER_33_240 ();
 FILLCELL_X1 FILLER_33_244 ();
 FILLCELL_X2 FILLER_33_251 ();
 FILLCELL_X1 FILLER_33_253 ();
 FILLCELL_X4 FILLER_33_275 ();
 FILLCELL_X16 FILLER_34_1 ();
 FILLCELL_X16 FILLER_34_82 ();
 FILLCELL_X4 FILLER_34_98 ();
 FILLCELL_X2 FILLER_34_102 ();
 FILLCELL_X1 FILLER_34_104 ();
 FILLCELL_X8 FILLER_34_122 ();
 FILLCELL_X1 FILLER_34_130 ();
 FILLCELL_X1 FILLER_34_148 ();
 FILLCELL_X4 FILLER_34_166 ();
 FILLCELL_X1 FILLER_34_195 ();
 FILLCELL_X16 FILLER_34_200 ();
 FILLCELL_X8 FILLER_34_216 ();
 FILLCELL_X1 FILLER_34_224 ();
 FILLCELL_X2 FILLER_34_245 ();
 FILLCELL_X8 FILLER_34_267 ();
 FILLCELL_X4 FILLER_34_275 ();
 FILLCELL_X2 FILLER_34_279 ();
 FILLCELL_X1 FILLER_34_281 ();
 FILLCELL_X1 FILLER_35_1 ();
 FILLCELL_X16 FILLER_35_6 ();
 FILLCELL_X4 FILLER_35_22 ();
 FILLCELL_X1 FILLER_35_26 ();
 FILLCELL_X4 FILLER_35_61 ();
 FILLCELL_X4 FILLER_35_82 ();
 FILLCELL_X16 FILLER_35_100 ();
 FILLCELL_X8 FILLER_35_178 ();
 FILLCELL_X2 FILLER_35_186 ();
 FILLCELL_X2 FILLER_35_210 ();
 FILLCELL_X1 FILLER_35_212 ();
 FILLCELL_X4 FILLER_35_215 ();
 FILLCELL_X2 FILLER_35_219 ();
 FILLCELL_X1 FILLER_35_221 ();
 FILLCELL_X2 FILLER_35_242 ();
 FILLCELL_X4 FILLER_35_253 ();
 FILLCELL_X2 FILLER_35_257 ();
 FILLCELL_X1 FILLER_35_259 ();
 FILLCELL_X2 FILLER_35_280 ();
 FILLCELL_X2 FILLER_36_50 ();
 FILLCELL_X1 FILLER_36_52 ();
 FILLCELL_X2 FILLER_36_67 ();
 FILLCELL_X4 FILLER_36_76 ();
 FILLCELL_X4 FILLER_36_87 ();
 FILLCELL_X4 FILLER_36_108 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X16 FILLER_36_161 ();
 FILLCELL_X8 FILLER_36_177 ();
 FILLCELL_X2 FILLER_36_185 ();
 FILLCELL_X1 FILLER_36_187 ();
 FILLCELL_X4 FILLER_36_210 ();
 FILLCELL_X1 FILLER_36_217 ();
 FILLCELL_X8 FILLER_36_225 ();
 FILLCELL_X4 FILLER_36_233 ();
 FILLCELL_X1 FILLER_36_237 ();
 FILLCELL_X1 FILLER_36_258 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X1 FILLER_37_65 ();
 FILLCELL_X8 FILLER_37_69 ();
 FILLCELL_X4 FILLER_37_77 ();
 FILLCELL_X2 FILLER_37_81 ();
 FILLCELL_X16 FILLER_37_100 ();
 FILLCELL_X8 FILLER_37_116 ();
 FILLCELL_X4 FILLER_37_124 ();
 FILLCELL_X1 FILLER_37_128 ();
 FILLCELL_X32 FILLER_37_133 ();
 FILLCELL_X16 FILLER_37_165 ();
 FILLCELL_X8 FILLER_37_181 ();
 FILLCELL_X4 FILLER_37_221 ();
 FILLCELL_X2 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_230 ();
 FILLCELL_X16 FILLER_37_264 ();
 FILLCELL_X2 FILLER_37_280 ();
endmodule
