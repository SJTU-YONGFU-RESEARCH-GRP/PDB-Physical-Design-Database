module axi_lite_master (arready,
    arvalid,
    awready,
    awvalid,
    bready,
    bvalid,
    clk,
    read_done,
    read_req,
    rready,
    rst_n,
    rvalid,
    wready,
    write_done,
    write_req,
    wvalid,
    araddr,
    awaddr,
    bresp,
    rdata,
    read_addr,
    read_data,
    rresp,
    wdata,
    write_addr,
    write_data,
    write_strb,
    wstrb);
 input arready;
 output arvalid;
 input awready;
 output awvalid;
 output bready;
 input bvalid;
 input clk;
 output read_done;
 input read_req;
 output rready;
 input rst_n;
 input rvalid;
 input wready;
 output write_done;
 input write_req;
 output wvalid;
 output [31:0] araddr;
 output [31:0] awaddr;
 input [1:0] bresp;
 input [31:0] rdata;
 input [31:0] read_addr;
 output [31:0] read_data;
 input [1:0] rresp;
 output [31:0] wdata;
 input [31:0] write_addr;
 input [31:0] write_data;
 input [3:0] write_strb;
 output [3:0] wstrb;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire _494_;
 wire _495_;
 wire _496_;
 wire _497_;
 wire _498_;
 wire _499_;
 wire _500_;
 wire _501_;
 wire _502_;
 wire _503_;
 wire _504_;
 wire _505_;
 wire _506_;
 wire _507_;
 wire _508_;
 wire _509_;
 wire _510_;
 wire _511_;
 wire _512_;
 wire \state_r[0] ;
 wire \state_r[1] ;
 wire \state_r[2] ;
 wire \state_r[3] ;
 wire \state_r[4] ;
 wire \state_r[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X2 _513_ (.A(rst_n),
    .Z(_146_));
 CLKBUF_X3 _514_ (.A(_146_),
    .Z(_147_));
 CLKBUF_X2 _515_ (.A(_147_),
    .Z(_148_));
 BUF_X4 _516_ (.A(\state_r[1] ),
    .Z(_149_));
 INV_X1 _517_ (.A(_149_),
    .ZN(_150_));
 AND2_X1 _518_ (.A1(net170),
    .A2(net1),
    .ZN(_151_));
 BUF_X1 _519_ (.A(read_req),
    .Z(_152_));
 CLKBUF_X3 _520_ (.A(\state_r[0] ),
    .Z(_153_));
 NAND2_X2 _521_ (.A1(_152_),
    .A2(_153_),
    .ZN(_154_));
 CLKBUF_X3 _522_ (.A(_154_),
    .Z(_155_));
 CLKBUF_X2 _523_ (.A(write_req),
    .Z(_156_));
 OAI22_X1 _524_ (.A1(_150_),
    .A2(_151_),
    .B1(_155_),
    .B2(_156_),
    .ZN(_157_));
 AND2_X1 _525_ (.A1(_148_),
    .A2(_157_),
    .ZN(_001_));
 CLKBUF_X3 _526_ (.A(\state_r[5] ),
    .Z(_158_));
 NAND3_X1 _527_ (.A1(_158_),
    .A2(net204),
    .A3(net3),
    .ZN(_159_));
 BUF_X4 _528_ (.A(\state_r[4] ),
    .Z(_160_));
 CLKBUF_X2 _529_ (.A(net238),
    .Z(_161_));
 NAND3_X4 _530_ (.A1(_160_),
    .A2(_161_),
    .A3(net68),
    .ZN(_162_));
 BUF_X4 _531_ (.A(_162_),
    .Z(_163_));
 INV_X1 _532_ (.A(_146_),
    .ZN(_164_));
 CLKBUF_X3 _533_ (.A(_164_),
    .Z(_165_));
 NOR2_X1 _534_ (.A1(_152_),
    .A2(_156_),
    .ZN(_166_));
 AOI21_X1 _535_ (.A(_165_),
    .B1(_153_),
    .B2(_166_),
    .ZN(_167_));
 NAND3_X1 _536_ (.A1(_159_),
    .A2(_163_),
    .A3(_167_),
    .ZN(_000_));
 CLKBUF_X3 _537_ (.A(\state_r[2] ),
    .Z(_168_));
 NAND2_X1 _538_ (.A1(net276),
    .A2(net69),
    .ZN(_169_));
 AND2_X1 _539_ (.A1(net203),
    .A2(net2),
    .ZN(_170_));
 BUF_X2 _540_ (.A(\state_r[3] ),
    .Z(_171_));
 AOI22_X1 _541_ (.A1(_168_),
    .A2(_169_),
    .B1(_170_),
    .B2(_171_),
    .ZN(_172_));
 NOR2_X1 _542_ (.A1(_165_),
    .A2(_172_),
    .ZN(_002_));
 NAND2_X2 _543_ (.A1(_156_),
    .A2(_153_),
    .ZN(_173_));
 BUF_X4 _544_ (.A(_173_),
    .Z(_174_));
 BUF_X4 _545_ (.A(_174_),
    .Z(_175_));
 NAND2_X1 _546_ (.A1(net203),
    .A2(net2),
    .ZN(_176_));
 NAND2_X1 _547_ (.A1(_171_),
    .A2(_176_),
    .ZN(_177_));
 AOI21_X1 _548_ (.A(_165_),
    .B1(_175_),
    .B2(_177_),
    .ZN(_003_));
 NAND2_X1 _549_ (.A1(_161_),
    .A2(net68),
    .ZN(_178_));
 AOI22_X1 _550_ (.A1(_149_),
    .A2(_151_),
    .B1(_178_),
    .B2(_160_),
    .ZN(_179_));
 NOR2_X1 _551_ (.A1(_165_),
    .A2(_179_),
    .ZN(_004_));
 NAND2_X1 _552_ (.A1(net204),
    .A2(net3),
    .ZN(_180_));
 AND2_X1 _553_ (.A1(net276),
    .A2(net69),
    .ZN(_181_));
 AOI22_X1 _554_ (.A1(_158_),
    .A2(_180_),
    .B1(_181_),
    .B2(_168_),
    .ZN(_182_));
 NOR2_X1 _555_ (.A1(_165_),
    .A2(_182_),
    .ZN(_005_));
 MUX2_X1 _556_ (.A(net36),
    .B(net138),
    .S(_155_),
    .Z(_183_));
 AND2_X1 _557_ (.A1(_148_),
    .A2(_183_),
    .ZN(_007_));
 MUX2_X1 _558_ (.A(net37),
    .B(net139),
    .S(_155_),
    .Z(_184_));
 AND2_X1 _559_ (.A1(_148_),
    .A2(_184_),
    .ZN(_008_));
 MUX2_X1 _560_ (.A(net38),
    .B(net140),
    .S(_155_),
    .Z(_185_));
 AND2_X1 _561_ (.A1(_148_),
    .A2(_185_),
    .ZN(_009_));
 MUX2_X1 _562_ (.A(net39),
    .B(net141),
    .S(_155_),
    .Z(_186_));
 AND2_X1 _563_ (.A1(_148_),
    .A2(_186_),
    .ZN(_010_));
 MUX2_X1 _564_ (.A(net40),
    .B(net142),
    .S(_155_),
    .Z(_187_));
 AND2_X1 _565_ (.A1(_148_),
    .A2(_187_),
    .ZN(_011_));
 MUX2_X1 _566_ (.A(net41),
    .B(net143),
    .S(_155_),
    .Z(_188_));
 AND2_X1 _567_ (.A1(_148_),
    .A2(_188_),
    .ZN(_012_));
 MUX2_X1 _568_ (.A(net42),
    .B(net144),
    .S(_155_),
    .Z(_189_));
 AND2_X1 _569_ (.A1(_148_),
    .A2(_189_),
    .ZN(_013_));
 MUX2_X1 _570_ (.A(net43),
    .B(net145),
    .S(_155_),
    .Z(_190_));
 AND2_X1 _571_ (.A1(_148_),
    .A2(_190_),
    .ZN(_014_));
 MUX2_X1 _572_ (.A(net44),
    .B(net146),
    .S(_155_),
    .Z(_191_));
 AND2_X1 _573_ (.A1(_148_),
    .A2(_191_),
    .ZN(_015_));
 CLKBUF_X2 _574_ (.A(_147_),
    .Z(_192_));
 CLKBUF_X3 _575_ (.A(_154_),
    .Z(_193_));
 MUX2_X1 _576_ (.A(net45),
    .B(net147),
    .S(_193_),
    .Z(_194_));
 AND2_X1 _577_ (.A1(_192_),
    .A2(_194_),
    .ZN(_016_));
 MUX2_X1 _578_ (.A(net46),
    .B(net148),
    .S(_193_),
    .Z(_195_));
 AND2_X1 _579_ (.A1(_192_),
    .A2(_195_),
    .ZN(_017_));
 MUX2_X1 _580_ (.A(net47),
    .B(net149),
    .S(_193_),
    .Z(_196_));
 AND2_X1 _581_ (.A1(_192_),
    .A2(_196_),
    .ZN(_018_));
 MUX2_X1 _582_ (.A(net48),
    .B(net150),
    .S(_193_),
    .Z(_197_));
 AND2_X1 _583_ (.A1(_192_),
    .A2(_197_),
    .ZN(_019_));
 MUX2_X1 _584_ (.A(net49),
    .B(net151),
    .S(_193_),
    .Z(_198_));
 AND2_X1 _585_ (.A1(_192_),
    .A2(_198_),
    .ZN(_020_));
 MUX2_X1 _586_ (.A(net50),
    .B(net152),
    .S(_193_),
    .Z(_199_));
 AND2_X1 _587_ (.A1(_192_),
    .A2(_199_),
    .ZN(_021_));
 MUX2_X1 _588_ (.A(net51),
    .B(net153),
    .S(_193_),
    .Z(_200_));
 AND2_X1 _589_ (.A1(_192_),
    .A2(_200_),
    .ZN(_022_));
 MUX2_X1 _590_ (.A(net52),
    .B(net154),
    .S(_193_),
    .Z(_201_));
 AND2_X1 _591_ (.A1(_192_),
    .A2(_201_),
    .ZN(_023_));
 MUX2_X1 _592_ (.A(net53),
    .B(net155),
    .S(_193_),
    .Z(_202_));
 AND2_X1 _593_ (.A1(_192_),
    .A2(_202_),
    .ZN(_024_));
 MUX2_X1 _594_ (.A(net54),
    .B(net156),
    .S(_193_),
    .Z(_203_));
 AND2_X1 _595_ (.A1(_192_),
    .A2(_203_),
    .ZN(_025_));
 CLKBUF_X2 _596_ (.A(_147_),
    .Z(_204_));
 CLKBUF_X3 _597_ (.A(_154_),
    .Z(_205_));
 MUX2_X1 _598_ (.A(net55),
    .B(net157),
    .S(_205_),
    .Z(_206_));
 AND2_X1 _599_ (.A1(_204_),
    .A2(_206_),
    .ZN(_026_));
 MUX2_X1 _600_ (.A(net56),
    .B(net158),
    .S(_205_),
    .Z(_207_));
 AND2_X1 _601_ (.A1(_204_),
    .A2(_207_),
    .ZN(_027_));
 MUX2_X1 _602_ (.A(net57),
    .B(net159),
    .S(_205_),
    .Z(_208_));
 AND2_X1 _603_ (.A1(_204_),
    .A2(_208_),
    .ZN(_028_));
 MUX2_X1 _604_ (.A(net58),
    .B(net160),
    .S(_205_),
    .Z(_209_));
 AND2_X1 _605_ (.A1(_204_),
    .A2(_209_),
    .ZN(_029_));
 MUX2_X1 _606_ (.A(net59),
    .B(net161),
    .S(_205_),
    .Z(_210_));
 AND2_X1 _607_ (.A1(_204_),
    .A2(_210_),
    .ZN(_030_));
 MUX2_X1 _608_ (.A(net60),
    .B(net162),
    .S(_205_),
    .Z(_211_));
 AND2_X1 _609_ (.A1(_204_),
    .A2(_211_),
    .ZN(_031_));
 MUX2_X1 _610_ (.A(net61),
    .B(net163),
    .S(_205_),
    .Z(_212_));
 AND2_X1 _611_ (.A1(_204_),
    .A2(_212_),
    .ZN(_032_));
 MUX2_X1 _612_ (.A(net62),
    .B(net164),
    .S(_205_),
    .Z(_213_));
 AND2_X1 _613_ (.A1(_204_),
    .A2(_213_),
    .ZN(_033_));
 MUX2_X1 _614_ (.A(net63),
    .B(net165),
    .S(_205_),
    .Z(_214_));
 AND2_X1 _615_ (.A1(_204_),
    .A2(_214_),
    .ZN(_034_));
 MUX2_X1 _616_ (.A(net64),
    .B(net166),
    .S(_205_),
    .Z(_215_));
 AND2_X1 _617_ (.A1(_204_),
    .A2(_215_),
    .ZN(_035_));
 CLKBUF_X2 _618_ (.A(_147_),
    .Z(_216_));
 MUX2_X1 _619_ (.A(net65),
    .B(net167),
    .S(_154_),
    .Z(_217_));
 AND2_X1 _620_ (.A1(_216_),
    .A2(_217_),
    .ZN(_036_));
 MUX2_X1 _621_ (.A(net66),
    .B(net168),
    .S(_154_),
    .Z(_218_));
 AND2_X1 _622_ (.A1(_216_),
    .A2(_218_),
    .ZN(_037_));
 MUX2_X1 _623_ (.A(net67),
    .B(net169),
    .S(_154_),
    .Z(_219_));
 AND2_X1 _624_ (.A1(_216_),
    .A2(_219_),
    .ZN(_038_));
 INV_X1 _625_ (.A(_153_),
    .ZN(_220_));
 OR4_X1 _626_ (.A1(_171_),
    .A2(_158_),
    .A3(_168_),
    .A4(_160_),
    .ZN(_221_));
 NAND2_X1 _627_ (.A1(net170),
    .A2(net1),
    .ZN(_222_));
 AOI21_X1 _628_ (.A(_221_),
    .B1(_222_),
    .B2(_149_),
    .ZN(_223_));
 NOR4_X2 _629_ (.A1(_171_),
    .A2(_158_),
    .A3(_168_),
    .A4(_160_),
    .ZN(_224_));
 OAI211_X2 _630_ (.A(_152_),
    .B(_224_),
    .C1(_151_),
    .C2(_150_),
    .ZN(_225_));
 INV_X1 _631_ (.A(net170),
    .ZN(_226_));
 AOI221_X1 _632_ (.A(_165_),
    .B1(_220_),
    .B2(_223_),
    .C1(_225_),
    .C2(_226_),
    .ZN(_039_));
 MUX2_X1 _633_ (.A(net70),
    .B(net171),
    .S(_175_),
    .Z(_227_));
 AND2_X1 _634_ (.A1(_216_),
    .A2(_227_),
    .ZN(_040_));
 MUX2_X1 _635_ (.A(net71),
    .B(net172),
    .S(_175_),
    .Z(_228_));
 AND2_X1 _636_ (.A1(_216_),
    .A2(_228_),
    .ZN(_041_));
 MUX2_X1 _637_ (.A(net72),
    .B(net173),
    .S(_175_),
    .Z(_229_));
 AND2_X1 _638_ (.A1(_216_),
    .A2(_229_),
    .ZN(_042_));
 MUX2_X1 _639_ (.A(net73),
    .B(net174),
    .S(_175_),
    .Z(_230_));
 AND2_X1 _640_ (.A1(_216_),
    .A2(_230_),
    .ZN(_043_));
 MUX2_X1 _641_ (.A(net74),
    .B(net175),
    .S(_175_),
    .Z(_231_));
 AND2_X1 _642_ (.A1(_216_),
    .A2(_231_),
    .ZN(_044_));
 MUX2_X1 _643_ (.A(net75),
    .B(net176),
    .S(_175_),
    .Z(_232_));
 AND2_X1 _644_ (.A1(_216_),
    .A2(_232_),
    .ZN(_045_));
 MUX2_X1 _645_ (.A(net76),
    .B(net177),
    .S(_175_),
    .Z(_233_));
 AND2_X1 _646_ (.A1(_216_),
    .A2(_233_),
    .ZN(_046_));
 CLKBUF_X2 _647_ (.A(_147_),
    .Z(_234_));
 MUX2_X1 _648_ (.A(net77),
    .B(net178),
    .S(_175_),
    .Z(_235_));
 AND2_X1 _649_ (.A1(_234_),
    .A2(_235_),
    .ZN(_047_));
 MUX2_X1 _650_ (.A(net78),
    .B(net179),
    .S(_175_),
    .Z(_236_));
 AND2_X1 _651_ (.A1(_234_),
    .A2(_236_),
    .ZN(_048_));
 CLKBUF_X3 _652_ (.A(_173_),
    .Z(_237_));
 MUX2_X1 _653_ (.A(net79),
    .B(net180),
    .S(_237_),
    .Z(_238_));
 AND2_X1 _654_ (.A1(_234_),
    .A2(_238_),
    .ZN(_049_));
 MUX2_X1 _655_ (.A(net80),
    .B(net181),
    .S(_237_),
    .Z(_239_));
 AND2_X1 _656_ (.A1(_234_),
    .A2(_239_),
    .ZN(_050_));
 MUX2_X1 _657_ (.A(net81),
    .B(net182),
    .S(_237_),
    .Z(_240_));
 AND2_X1 _658_ (.A1(_234_),
    .A2(_240_),
    .ZN(_051_));
 MUX2_X1 _659_ (.A(net82),
    .B(net183),
    .S(_237_),
    .Z(_241_));
 AND2_X1 _660_ (.A1(_234_),
    .A2(_241_),
    .ZN(_052_));
 MUX2_X1 _661_ (.A(net83),
    .B(net184),
    .S(_237_),
    .Z(_242_));
 AND2_X1 _662_ (.A1(_234_),
    .A2(_242_),
    .ZN(_053_));
 MUX2_X1 _663_ (.A(net84),
    .B(net185),
    .S(_237_),
    .Z(_243_));
 AND2_X1 _664_ (.A1(_234_),
    .A2(_243_),
    .ZN(_054_));
 MUX2_X1 _665_ (.A(net85),
    .B(net186),
    .S(_237_),
    .Z(_244_));
 AND2_X1 _666_ (.A1(_234_),
    .A2(_244_),
    .ZN(_055_));
 MUX2_X1 _667_ (.A(net86),
    .B(net187),
    .S(_237_),
    .Z(_245_));
 AND2_X1 _668_ (.A1(_234_),
    .A2(_245_),
    .ZN(_056_));
 CLKBUF_X2 _669_ (.A(_147_),
    .Z(_246_));
 MUX2_X1 _670_ (.A(net87),
    .B(net188),
    .S(_237_),
    .Z(_247_));
 AND2_X1 _671_ (.A1(_246_),
    .A2(_247_),
    .ZN(_057_));
 MUX2_X1 _672_ (.A(net88),
    .B(net189),
    .S(_237_),
    .Z(_248_));
 AND2_X1 _673_ (.A1(_246_),
    .A2(_248_),
    .ZN(_058_));
 CLKBUF_X3 _674_ (.A(_173_),
    .Z(_249_));
 MUX2_X1 _675_ (.A(net89),
    .B(net190),
    .S(_249_),
    .Z(_250_));
 AND2_X1 _676_ (.A1(_246_),
    .A2(_250_),
    .ZN(_059_));
 MUX2_X1 _677_ (.A(net90),
    .B(net191),
    .S(_249_),
    .Z(_251_));
 AND2_X1 _678_ (.A1(_246_),
    .A2(_251_),
    .ZN(_060_));
 MUX2_X1 _679_ (.A(net91),
    .B(net192),
    .S(_249_),
    .Z(_252_));
 AND2_X1 _680_ (.A1(_246_),
    .A2(_252_),
    .ZN(_061_));
 MUX2_X1 _681_ (.A(net92),
    .B(net193),
    .S(_249_),
    .Z(_253_));
 AND2_X1 _682_ (.A1(_246_),
    .A2(_253_),
    .ZN(_062_));
 MUX2_X1 _683_ (.A(net93),
    .B(net194),
    .S(_249_),
    .Z(_254_));
 AND2_X1 _684_ (.A1(_246_),
    .A2(_254_),
    .ZN(_063_));
 MUX2_X1 _685_ (.A(net94),
    .B(net195),
    .S(_249_),
    .Z(_255_));
 AND2_X1 _686_ (.A1(_246_),
    .A2(_255_),
    .ZN(_064_));
 MUX2_X1 _687_ (.A(net95),
    .B(net196),
    .S(_249_),
    .Z(_256_));
 AND2_X1 _688_ (.A1(_246_),
    .A2(_256_),
    .ZN(_065_));
 MUX2_X1 _689_ (.A(net96),
    .B(net197),
    .S(_249_),
    .Z(_257_));
 AND2_X1 _690_ (.A1(_246_),
    .A2(_257_),
    .ZN(_066_));
 BUF_X2 _691_ (.A(_147_),
    .Z(_258_));
 MUX2_X1 _692_ (.A(net97),
    .B(net198),
    .S(_249_),
    .Z(_259_));
 AND2_X1 _693_ (.A1(_258_),
    .A2(_259_),
    .ZN(_067_));
 MUX2_X1 _694_ (.A(net98),
    .B(net199),
    .S(_249_),
    .Z(_260_));
 AND2_X1 _695_ (.A1(_258_),
    .A2(_260_),
    .ZN(_068_));
 CLKBUF_X3 _696_ (.A(_173_),
    .Z(_261_));
 MUX2_X1 _697_ (.A(net99),
    .B(net200),
    .S(_261_),
    .Z(_262_));
 AND2_X1 _698_ (.A1(_258_),
    .A2(_262_),
    .ZN(_069_));
 MUX2_X1 _699_ (.A(net100),
    .B(net201),
    .S(_261_),
    .Z(_263_));
 AND2_X1 _700_ (.A1(_258_),
    .A2(_263_),
    .ZN(_070_));
 MUX2_X1 _701_ (.A(net101),
    .B(net202),
    .S(_261_),
    .Z(_264_));
 AND2_X1 _702_ (.A1(_258_),
    .A2(_264_),
    .ZN(_071_));
 OR4_X1 _703_ (.A1(_149_),
    .A2(_158_),
    .A3(_168_),
    .A4(\state_r[4] ),
    .ZN(_265_));
 AOI21_X1 _704_ (.A(_265_),
    .B1(_176_),
    .B2(_171_),
    .ZN(_266_));
 NOR4_X2 _705_ (.A1(_149_),
    .A2(_158_),
    .A3(_168_),
    .A4(_160_),
    .ZN(_267_));
 INV_X1 _706_ (.A(_171_),
    .ZN(_268_));
 OAI211_X2 _707_ (.A(_156_),
    .B(_267_),
    .C1(_170_),
    .C2(_268_),
    .ZN(_269_));
 INV_X1 _708_ (.A(net203),
    .ZN(_270_));
 AOI221_X1 _709_ (.A(_165_),
    .B1(_220_),
    .B2(_266_),
    .C1(_269_),
    .C2(_270_),
    .ZN(_072_));
 INV_X1 _710_ (.A(_168_),
    .ZN(_271_));
 OR4_X1 _711_ (.A1(_171_),
    .A2(_153_),
    .A3(_149_),
    .A4(\state_r[4] ),
    .ZN(_272_));
 AOI21_X1 _712_ (.A(_006_),
    .B1(net204),
    .B2(net3),
    .ZN(_273_));
 NOR2_X1 _713_ (.A1(_272_),
    .A2(_273_),
    .ZN(_274_));
 OR3_X1 _714_ (.A1(_169_),
    .A2(_272_),
    .A3(_273_),
    .ZN(_275_));
 INV_X1 _715_ (.A(net204),
    .ZN(_276_));
 AOI221_X1 _716_ (.A(_165_),
    .B1(_271_),
    .B2(_274_),
    .C1(_275_),
    .C2(_276_),
    .ZN(_073_));
 MUX2_X1 _717_ (.A(net4),
    .B(net205),
    .S(_163_),
    .Z(_277_));
 AND2_X1 _718_ (.A1(_258_),
    .A2(_277_),
    .ZN(_074_));
 MUX2_X1 _719_ (.A(net5),
    .B(net206),
    .S(_163_),
    .Z(_278_));
 AND2_X1 _720_ (.A1(_258_),
    .A2(_278_),
    .ZN(_075_));
 MUX2_X1 _721_ (.A(net6),
    .B(net207),
    .S(_163_),
    .Z(_279_));
 AND2_X1 _722_ (.A1(_258_),
    .A2(_279_),
    .ZN(_076_));
 MUX2_X1 _723_ (.A(net7),
    .B(net208),
    .S(_163_),
    .Z(_280_));
 AND2_X1 _724_ (.A1(_258_),
    .A2(_280_),
    .ZN(_077_));
 MUX2_X1 _725_ (.A(net8),
    .B(net209),
    .S(_163_),
    .Z(_281_));
 AND2_X1 _726_ (.A1(_258_),
    .A2(_281_),
    .ZN(_078_));
 CLKBUF_X2 _727_ (.A(_146_),
    .Z(_282_));
 MUX2_X1 _728_ (.A(net9),
    .B(net210),
    .S(_163_),
    .Z(_283_));
 AND2_X1 _729_ (.A1(_282_),
    .A2(_283_),
    .ZN(_079_));
 MUX2_X1 _730_ (.A(net10),
    .B(net211),
    .S(_163_),
    .Z(_284_));
 AND2_X1 _731_ (.A1(_282_),
    .A2(_284_),
    .ZN(_080_));
 MUX2_X1 _732_ (.A(net11),
    .B(net212),
    .S(_163_),
    .Z(_285_));
 AND2_X1 _733_ (.A1(_282_),
    .A2(_285_),
    .ZN(_081_));
 CLKBUF_X3 _734_ (.A(_162_),
    .Z(_286_));
 MUX2_X1 _735_ (.A(net12),
    .B(net213),
    .S(_286_),
    .Z(_287_));
 AND2_X1 _736_ (.A1(_282_),
    .A2(_287_),
    .ZN(_082_));
 MUX2_X1 _737_ (.A(net13),
    .B(net214),
    .S(_286_),
    .Z(_288_));
 AND2_X1 _738_ (.A1(_282_),
    .A2(_288_),
    .ZN(_083_));
 MUX2_X1 _739_ (.A(net14),
    .B(net215),
    .S(_286_),
    .Z(_289_));
 AND2_X1 _740_ (.A1(_282_),
    .A2(_289_),
    .ZN(_084_));
 MUX2_X1 _741_ (.A(net15),
    .B(net216),
    .S(_286_),
    .Z(_290_));
 AND2_X1 _742_ (.A1(_282_),
    .A2(_290_),
    .ZN(_085_));
 MUX2_X1 _743_ (.A(net16),
    .B(net217),
    .S(_286_),
    .Z(_291_));
 AND2_X1 _744_ (.A1(_282_),
    .A2(_291_),
    .ZN(_086_));
 MUX2_X1 _745_ (.A(net17),
    .B(net218),
    .S(_286_),
    .Z(_292_));
 AND2_X1 _746_ (.A1(_282_),
    .A2(_292_),
    .ZN(_087_));
 MUX2_X1 _747_ (.A(net18),
    .B(net219),
    .S(_286_),
    .Z(_293_));
 AND2_X1 _748_ (.A1(_282_),
    .A2(_293_),
    .ZN(_088_));
 CLKBUF_X2 _749_ (.A(_146_),
    .Z(_294_));
 MUX2_X1 _750_ (.A(net19),
    .B(net220),
    .S(_286_),
    .Z(_295_));
 AND2_X1 _751_ (.A1(_294_),
    .A2(_295_),
    .ZN(_089_));
 MUX2_X1 _752_ (.A(net20),
    .B(net221),
    .S(_286_),
    .Z(_296_));
 AND2_X1 _753_ (.A1(_294_),
    .A2(_296_),
    .ZN(_090_));
 MUX2_X1 _754_ (.A(net21),
    .B(net222),
    .S(_286_),
    .Z(_297_));
 AND2_X1 _755_ (.A1(_294_),
    .A2(_297_),
    .ZN(_091_));
 CLKBUF_X3 _756_ (.A(_162_),
    .Z(_298_));
 MUX2_X1 _757_ (.A(net22),
    .B(net223),
    .S(_298_),
    .Z(_299_));
 AND2_X1 _758_ (.A1(_294_),
    .A2(_299_),
    .ZN(_092_));
 MUX2_X1 _759_ (.A(net23),
    .B(net224),
    .S(_298_),
    .Z(_300_));
 AND2_X1 _760_ (.A1(_294_),
    .A2(_300_),
    .ZN(_093_));
 MUX2_X1 _761_ (.A(net24),
    .B(net225),
    .S(_298_),
    .Z(_301_));
 AND2_X1 _762_ (.A1(_294_),
    .A2(_301_),
    .ZN(_094_));
 MUX2_X1 _763_ (.A(net25),
    .B(net226),
    .S(_298_),
    .Z(_302_));
 AND2_X1 _764_ (.A1(_294_),
    .A2(_302_),
    .ZN(_095_));
 MUX2_X1 _765_ (.A(net26),
    .B(net227),
    .S(_298_),
    .Z(_303_));
 AND2_X1 _766_ (.A1(_294_),
    .A2(_303_),
    .ZN(_096_));
 MUX2_X1 _767_ (.A(net27),
    .B(net228),
    .S(_298_),
    .Z(_304_));
 AND2_X1 _768_ (.A1(_294_),
    .A2(_304_),
    .ZN(_097_));
 MUX2_X1 _769_ (.A(net28),
    .B(net229),
    .S(_298_),
    .Z(_305_));
 AND2_X1 _770_ (.A1(_294_),
    .A2(_305_),
    .ZN(_098_));
 CLKBUF_X2 _771_ (.A(_146_),
    .Z(_306_));
 MUX2_X1 _772_ (.A(net29),
    .B(net230),
    .S(_298_),
    .Z(_307_));
 AND2_X1 _773_ (.A1(_306_),
    .A2(_307_),
    .ZN(_099_));
 MUX2_X1 _774_ (.A(net30),
    .B(net231),
    .S(_298_),
    .Z(_308_));
 AND2_X1 _775_ (.A1(_306_),
    .A2(_308_),
    .ZN(_100_));
 MUX2_X1 _776_ (.A(net31),
    .B(net232),
    .S(_298_),
    .Z(_309_));
 AND2_X1 _777_ (.A1(_306_),
    .A2(_309_),
    .ZN(_101_));
 MUX2_X1 _778_ (.A(net32),
    .B(net233),
    .S(_162_),
    .Z(_310_));
 AND2_X1 _779_ (.A1(_306_),
    .A2(_310_),
    .ZN(_102_));
 MUX2_X1 _780_ (.A(net33),
    .B(net234),
    .S(_162_),
    .Z(_311_));
 AND2_X1 _781_ (.A1(_306_),
    .A2(_311_),
    .ZN(_103_));
 MUX2_X1 _782_ (.A(net34),
    .B(net235),
    .S(_162_),
    .Z(_312_));
 AND2_X1 _783_ (.A1(_306_),
    .A2(_312_),
    .ZN(_104_));
 MUX2_X1 _784_ (.A(net35),
    .B(net236),
    .S(_162_),
    .Z(_313_));
 AND2_X1 _785_ (.A1(_306_),
    .A2(_313_),
    .ZN(_105_));
 OAI21_X1 _786_ (.A(net237),
    .B1(_160_),
    .B2(_220_),
    .ZN(_314_));
 AOI21_X1 _787_ (.A(_165_),
    .B1(_163_),
    .B2(_314_),
    .ZN(_106_));
 OR4_X1 _788_ (.A1(_171_),
    .A2(_153_),
    .A3(\state_r[5] ),
    .A4(_168_),
    .ZN(_315_));
 AOI21_X1 _789_ (.A(_315_),
    .B1(_178_),
    .B2(_160_),
    .ZN(_316_));
 NOR4_X2 _790_ (.A1(_171_),
    .A2(_153_),
    .A3(_158_),
    .A4(_168_),
    .ZN(_317_));
 AND2_X1 _791_ (.A1(_161_),
    .A2(net68),
    .ZN(_318_));
 INV_X1 _792_ (.A(_160_),
    .ZN(_319_));
 OAI211_X2 _793_ (.A(_151_),
    .B(_317_),
    .C1(_318_),
    .C2(_319_),
    .ZN(_320_));
 INV_X1 _794_ (.A(_161_),
    .ZN(_321_));
 AOI221_X1 _795_ (.A(_164_),
    .B1(_150_),
    .B2(_316_),
    .C1(_320_),
    .C2(_321_),
    .ZN(_107_));
 MUX2_X1 _796_ (.A(net102),
    .B(net239),
    .S(_261_),
    .Z(_322_));
 AND2_X1 _797_ (.A1(_306_),
    .A2(_322_),
    .ZN(_108_));
 MUX2_X1 _798_ (.A(net103),
    .B(net240),
    .S(_261_),
    .Z(_323_));
 AND2_X1 _799_ (.A1(_306_),
    .A2(_323_),
    .ZN(_109_));
 MUX2_X1 _800_ (.A(net104),
    .B(net241),
    .S(_261_),
    .Z(_324_));
 AND2_X1 _801_ (.A1(_306_),
    .A2(_324_),
    .ZN(_110_));
 CLKBUF_X2 _802_ (.A(_146_),
    .Z(_325_));
 MUX2_X1 _803_ (.A(net105),
    .B(net242),
    .S(_261_),
    .Z(_326_));
 AND2_X1 _804_ (.A1(_325_),
    .A2(_326_),
    .ZN(_111_));
 MUX2_X1 _805_ (.A(net106),
    .B(net243),
    .S(_261_),
    .Z(_327_));
 AND2_X1 _806_ (.A1(_325_),
    .A2(_327_),
    .ZN(_112_));
 MUX2_X1 _807_ (.A(net107),
    .B(net244),
    .S(_261_),
    .Z(_328_));
 AND2_X1 _808_ (.A1(_325_),
    .A2(_328_),
    .ZN(_113_));
 MUX2_X1 _809_ (.A(net108),
    .B(net245),
    .S(_261_),
    .Z(_329_));
 AND2_X1 _810_ (.A1(_325_),
    .A2(_329_),
    .ZN(_114_));
 CLKBUF_X3 _811_ (.A(_173_),
    .Z(_330_));
 MUX2_X1 _812_ (.A(net109),
    .B(net246),
    .S(_330_),
    .Z(_331_));
 AND2_X1 _813_ (.A1(_325_),
    .A2(_331_),
    .ZN(_115_));
 MUX2_X1 _814_ (.A(net110),
    .B(net247),
    .S(_330_),
    .Z(_332_));
 AND2_X1 _815_ (.A1(_325_),
    .A2(_332_),
    .ZN(_116_));
 MUX2_X1 _816_ (.A(net111),
    .B(net248),
    .S(_330_),
    .Z(_333_));
 AND2_X1 _817_ (.A1(_325_),
    .A2(_333_),
    .ZN(_117_));
 MUX2_X1 _818_ (.A(net112),
    .B(net249),
    .S(_330_),
    .Z(_334_));
 AND2_X1 _819_ (.A1(_325_),
    .A2(_334_),
    .ZN(_118_));
 MUX2_X1 _820_ (.A(net113),
    .B(net250),
    .S(_330_),
    .Z(_335_));
 AND2_X1 _821_ (.A1(_325_),
    .A2(_335_),
    .ZN(_119_));
 MUX2_X1 _822_ (.A(net114),
    .B(net251),
    .S(_330_),
    .Z(_336_));
 AND2_X1 _823_ (.A1(_325_),
    .A2(_336_),
    .ZN(_120_));
 CLKBUF_X2 _824_ (.A(_146_),
    .Z(_337_));
 MUX2_X1 _825_ (.A(net115),
    .B(net252),
    .S(_330_),
    .Z(_338_));
 AND2_X1 _826_ (.A1(_337_),
    .A2(_338_),
    .ZN(_121_));
 MUX2_X1 _827_ (.A(net116),
    .B(net253),
    .S(_330_),
    .Z(_339_));
 AND2_X1 _828_ (.A1(_337_),
    .A2(_339_),
    .ZN(_122_));
 MUX2_X1 _829_ (.A(net117),
    .B(net254),
    .S(_330_),
    .Z(_340_));
 AND2_X1 _830_ (.A1(_337_),
    .A2(_340_),
    .ZN(_123_));
 MUX2_X1 _831_ (.A(net118),
    .B(net255),
    .S(_330_),
    .Z(_341_));
 AND2_X1 _832_ (.A1(_337_),
    .A2(_341_),
    .ZN(_124_));
 CLKBUF_X3 _833_ (.A(_173_),
    .Z(_342_));
 MUX2_X1 _834_ (.A(net119),
    .B(net256),
    .S(_342_),
    .Z(_343_));
 AND2_X1 _835_ (.A1(_337_),
    .A2(_343_),
    .ZN(_125_));
 MUX2_X1 _836_ (.A(net120),
    .B(net257),
    .S(_342_),
    .Z(_344_));
 AND2_X1 _837_ (.A1(_337_),
    .A2(_344_),
    .ZN(_126_));
 MUX2_X1 _838_ (.A(net121),
    .B(net258),
    .S(_342_),
    .Z(_345_));
 AND2_X1 _839_ (.A1(_337_),
    .A2(_345_),
    .ZN(_127_));
 MUX2_X1 _840_ (.A(net122),
    .B(net259),
    .S(_342_),
    .Z(_346_));
 AND2_X1 _841_ (.A1(_337_),
    .A2(_346_),
    .ZN(_128_));
 MUX2_X1 _842_ (.A(net123),
    .B(net260),
    .S(_342_),
    .Z(_347_));
 AND2_X1 _843_ (.A1(_337_),
    .A2(_347_),
    .ZN(_129_));
 MUX2_X1 _844_ (.A(net124),
    .B(net261),
    .S(_342_),
    .Z(_348_));
 AND2_X1 _845_ (.A1(_337_),
    .A2(_348_),
    .ZN(_130_));
 BUF_X2 _846_ (.A(_146_),
    .Z(_349_));
 MUX2_X1 _847_ (.A(net125),
    .B(net262),
    .S(_342_),
    .Z(_350_));
 AND2_X1 _848_ (.A1(_349_),
    .A2(_350_),
    .ZN(_131_));
 MUX2_X1 _849_ (.A(net126),
    .B(net263),
    .S(_342_),
    .Z(_351_));
 AND2_X1 _850_ (.A1(_349_),
    .A2(_351_),
    .ZN(_132_));
 MUX2_X1 _851_ (.A(net127),
    .B(net264),
    .S(_342_),
    .Z(_352_));
 AND2_X1 _852_ (.A1(_349_),
    .A2(_352_),
    .ZN(_133_));
 MUX2_X1 _853_ (.A(net128),
    .B(net265),
    .S(_342_),
    .Z(_353_));
 AND2_X1 _854_ (.A1(_349_),
    .A2(_353_),
    .ZN(_134_));
 MUX2_X1 _855_ (.A(net129),
    .B(net266),
    .S(_174_),
    .Z(_354_));
 AND2_X1 _856_ (.A1(_349_),
    .A2(_354_),
    .ZN(_135_));
 MUX2_X1 _857_ (.A(net130),
    .B(net267),
    .S(_174_),
    .Z(_355_));
 AND2_X1 _858_ (.A1(_349_),
    .A2(_355_),
    .ZN(_136_));
 MUX2_X1 _859_ (.A(net131),
    .B(net268),
    .S(_174_),
    .Z(_356_));
 AND2_X1 _860_ (.A1(_349_),
    .A2(_356_),
    .ZN(_137_));
 MUX2_X1 _861_ (.A(net132),
    .B(net269),
    .S(_174_),
    .Z(_357_));
 AND2_X1 _862_ (.A1(_349_),
    .A2(_357_),
    .ZN(_138_));
 MUX2_X1 _863_ (.A(net133),
    .B(net270),
    .S(_174_),
    .Z(_358_));
 AND2_X1 _864_ (.A1(_349_),
    .A2(_358_),
    .ZN(_139_));
 OAI21_X1 _865_ (.A(net271),
    .B1(_158_),
    .B2(_220_),
    .ZN(_359_));
 AOI21_X1 _866_ (.A(_165_),
    .B1(_159_),
    .B2(_359_),
    .ZN(_140_));
 MUX2_X1 _867_ (.A(net134),
    .B(net272),
    .S(_174_),
    .Z(_360_));
 AND2_X1 _868_ (.A1(_349_),
    .A2(_360_),
    .ZN(_141_));
 MUX2_X1 _869_ (.A(net135),
    .B(net273),
    .S(_174_),
    .Z(_361_));
 AND2_X1 _870_ (.A1(_147_),
    .A2(_361_),
    .ZN(_142_));
 MUX2_X1 _871_ (.A(net136),
    .B(net274),
    .S(_174_),
    .Z(_362_));
 AND2_X1 _872_ (.A1(_147_),
    .A2(_362_),
    .ZN(_143_));
 MUX2_X1 _873_ (.A(net137),
    .B(net275),
    .S(_174_),
    .Z(_363_));
 AND2_X1 _874_ (.A1(_147_),
    .A2(_363_),
    .ZN(_144_));
 INV_X1 _875_ (.A(net276),
    .ZN(_364_));
 NOR4_X1 _876_ (.A1(_153_),
    .A2(_149_),
    .A3(_158_),
    .A4(_160_),
    .ZN(_365_));
 OAI221_X1 _877_ (.A(_365_),
    .B1(_181_),
    .B2(_271_),
    .C1(_268_),
    .C2(_170_),
    .ZN(_366_));
 OR4_X1 _878_ (.A1(_153_),
    .A2(_149_),
    .A3(_158_),
    .A4(_160_),
    .ZN(_367_));
 AOI21_X1 _879_ (.A(_367_),
    .B1(_169_),
    .B2(_168_),
    .ZN(_368_));
 AOI221_X1 _880_ (.A(_164_),
    .B1(_364_),
    .B2(_366_),
    .C1(_368_),
    .C2(_268_),
    .ZN(_145_));
 DFF_X1 \araddr[0]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_4_14_0_clk),
    .Q(net138),
    .QN(_506_));
 DFF_X1 \araddr[10]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_4_11_0_clk),
    .Q(net139),
    .QN(_505_));
 DFF_X1 \araddr[11]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_4_11_0_clk),
    .Q(net140),
    .QN(_504_));
 DFF_X1 \araddr[12]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_4_11_0_clk),
    .Q(net141),
    .QN(_503_));
 DFF_X1 \araddr[13]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_4_14_0_clk),
    .Q(net142),
    .QN(_502_));
 DFF_X1 \araddr[14]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_4_14_0_clk),
    .Q(net143),
    .QN(_501_));
 DFF_X1 \araddr[15]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_4_11_0_clk),
    .Q(net144),
    .QN(_500_));
 DFF_X1 \araddr[16]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_4_14_0_clk),
    .Q(net145),
    .QN(_499_));
 DFF_X1 \araddr[17]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_4_14_0_clk),
    .Q(net146),
    .QN(_498_));
 DFF_X1 \araddr[18]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_4_15_0_clk),
    .Q(net147),
    .QN(_497_));
 DFF_X1 \araddr[19]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_4_15_0_clk),
    .Q(net148),
    .QN(_496_));
 DFF_X1 \araddr[1]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_4_15_0_clk),
    .Q(net149),
    .QN(_495_));
 DFF_X1 \araddr[20]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_4_15_0_clk),
    .Q(net150),
    .QN(_494_));
 DFF_X1 \araddr[21]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_4_13_0_clk),
    .Q(net151),
    .QN(_493_));
 DFF_X1 \araddr[22]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_4_15_0_clk),
    .Q(net152),
    .QN(_492_));
 DFF_X1 \araddr[23]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_4_13_0_clk),
    .Q(net153),
    .QN(_491_));
 DFF_X1 \araddr[24]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_4_13_0_clk),
    .Q(net154),
    .QN(_490_));
 DFF_X1 \araddr[25]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_4_15_0_clk),
    .Q(net155),
    .QN(_489_));
 DFF_X1 \araddr[26]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_4_13_0_clk),
    .Q(net156),
    .QN(_488_));
 DFF_X1 \araddr[27]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_4_15_0_clk),
    .Q(net157),
    .QN(_487_));
 DFF_X1 \araddr[28]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_4_15_0_clk),
    .Q(net158),
    .QN(_486_));
 DFF_X1 \araddr[29]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_4_15_0_clk),
    .Q(net159),
    .QN(_485_));
 DFF_X1 \araddr[2]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_4_15_0_clk),
    .Q(net160),
    .QN(_484_));
 DFF_X1 \araddr[30]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_4_15_0_clk),
    .Q(net161),
    .QN(_483_));
 DFF_X1 \araddr[31]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_4_15_0_clk),
    .Q(net162),
    .QN(_482_));
 DFF_X1 \araddr[3]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_4_14_0_clk),
    .Q(net163),
    .QN(_481_));
 DFF_X1 \araddr[4]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_4_14_0_clk),
    .Q(net164),
    .QN(_480_));
 DFF_X1 \araddr[5]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_4_15_0_clk),
    .Q(net165),
    .QN(_479_));
 DFF_X1 \araddr[6]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_4_14_0_clk),
    .Q(net166),
    .QN(_478_));
 DFF_X1 \araddr[7]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_4_13_0_clk),
    .Q(net167),
    .QN(_477_));
 DFF_X1 \araddr[8]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_4_13_0_clk),
    .Q(net168),
    .QN(_476_));
 DFF_X1 \araddr[9]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_4_13_0_clk),
    .Q(net169),
    .QN(_475_));
 DFF_X1 \arvalid$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_4_9_0_clk),
    .Q(net170),
    .QN(_474_));
 DFF_X1 \awaddr[0]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_4_6_0_clk),
    .Q(net171),
    .QN(_473_));
 DFF_X1 \awaddr[10]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_4_13_0_clk),
    .Q(net172),
    .QN(_472_));
 DFF_X1 \awaddr[11]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_4_13_0_clk),
    .Q(net173),
    .QN(_471_));
 DFF_X1 \awaddr[12]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_4_7_0_clk),
    .Q(net174),
    .QN(_470_));
 DFF_X1 \awaddr[13]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_4_6_0_clk),
    .Q(net175),
    .QN(_469_));
 DFF_X1 \awaddr[14]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_4_6_0_clk),
    .Q(net176),
    .QN(_468_));
 DFF_X1 \awaddr[15]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_4_7_0_clk),
    .Q(net177),
    .QN(_467_));
 DFF_X1 \awaddr[16]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_4_7_0_clk),
    .Q(net178),
    .QN(_466_));
 DFF_X1 \awaddr[17]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_4_7_0_clk),
    .Q(net179),
    .QN(_465_));
 DFF_X1 \awaddr[18]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_4_5_0_clk),
    .Q(net180),
    .QN(_464_));
 DFF_X1 \awaddr[19]$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_4_5_0_clk),
    .Q(net181),
    .QN(_463_));
 DFF_X1 \awaddr[1]$_SDFFE_PN0P_  (.D(_051_),
    .CK(clknet_4_5_0_clk),
    .Q(net182),
    .QN(_462_));
 DFF_X1 \awaddr[20]$_SDFFE_PN0P_  (.D(_052_),
    .CK(clknet_4_5_0_clk),
    .Q(net183),
    .QN(_461_));
 DFF_X1 \awaddr[21]$_SDFFE_PN0P_  (.D(_053_),
    .CK(clknet_4_7_0_clk),
    .Q(net184),
    .QN(_460_));
 DFF_X1 \awaddr[22]$_SDFFE_PN0P_  (.D(_054_),
    .CK(clknet_4_5_0_clk),
    .Q(net185),
    .QN(_459_));
 DFF_X1 \awaddr[23]$_SDFFE_PN0P_  (.D(_055_),
    .CK(clknet_4_5_0_clk),
    .Q(net186),
    .QN(_458_));
 DFF_X1 \awaddr[24]$_SDFFE_PN0P_  (.D(_056_),
    .CK(clknet_4_7_0_clk),
    .Q(net187),
    .QN(_457_));
 DFF_X1 \awaddr[25]$_SDFFE_PN0P_  (.D(_057_),
    .CK(clknet_4_5_0_clk),
    .Q(net188),
    .QN(_456_));
 DFF_X1 \awaddr[26]$_SDFFE_PN0P_  (.D(_058_),
    .CK(clknet_4_5_0_clk),
    .Q(net189),
    .QN(_455_));
 DFF_X1 \awaddr[27]$_SDFFE_PN0P_  (.D(_059_),
    .CK(clknet_4_5_0_clk),
    .Q(net190),
    .QN(_454_));
 DFF_X1 \awaddr[28]$_SDFFE_PN0P_  (.D(_060_),
    .CK(clknet_4_5_0_clk),
    .Q(net191),
    .QN(_453_));
 DFF_X1 \awaddr[29]$_SDFFE_PN0P_  (.D(_061_),
    .CK(clknet_4_5_0_clk),
    .Q(net192),
    .QN(_452_));
 DFF_X1 \awaddr[2]$_SDFFE_PN0P_  (.D(_062_),
    .CK(clknet_4_5_0_clk),
    .Q(net193),
    .QN(_451_));
 DFF_X1 \awaddr[30]$_SDFFE_PN0P_  (.D(_063_),
    .CK(clknet_4_4_0_clk),
    .Q(net194),
    .QN(_450_));
 DFF_X1 \awaddr[31]$_SDFFE_PN0P_  (.D(_064_),
    .CK(clknet_4_7_0_clk),
    .Q(net195),
    .QN(_449_));
 DFF_X1 \awaddr[3]$_SDFFE_PN0P_  (.D(_065_),
    .CK(clknet_4_4_0_clk),
    .Q(net196),
    .QN(_448_));
 DFF_X1 \awaddr[4]$_SDFFE_PN0P_  (.D(_066_),
    .CK(clknet_4_4_0_clk),
    .Q(net197),
    .QN(_447_));
 DFF_X1 \awaddr[5]$_SDFFE_PN0P_  (.D(_067_),
    .CK(clknet_4_4_0_clk),
    .Q(net198),
    .QN(_446_));
 DFF_X1 \awaddr[6]$_SDFFE_PN0P_  (.D(_068_),
    .CK(clknet_4_4_0_clk),
    .Q(net199),
    .QN(_445_));
 DFF_X1 \awaddr[7]$_SDFFE_PN0P_  (.D(_069_),
    .CK(clknet_4_2_0_clk),
    .Q(net200),
    .QN(_444_));
 DFF_X1 \awaddr[8]$_SDFFE_PN0P_  (.D(_070_),
    .CK(clknet_4_3_0_clk),
    .Q(net201),
    .QN(_443_));
 DFF_X1 \awaddr[9]$_SDFFE_PN0P_  (.D(_071_),
    .CK(clknet_4_3_0_clk),
    .Q(net202),
    .QN(_442_));
 DFF_X1 \awvalid$_SDFFE_PN0P_  (.D(_072_),
    .CK(clknet_4_12_0_clk),
    .Q(net203),
    .QN(_441_));
 DFF_X2 \bready$_SDFFE_PN0P_  (.D(_073_),
    .CK(clknet_4_12_0_clk),
    .Q(net204),
    .QN(_440_));
 DFF_X1 \read_data[0]$_SDFFE_PN0P_  (.D(_074_),
    .CK(clknet_4_0_0_clk),
    .Q(net205),
    .QN(_439_));
 DFF_X1 \read_data[10]$_SDFFE_PN0P_  (.D(_075_),
    .CK(clknet_4_3_0_clk),
    .Q(net206),
    .QN(_438_));
 DFF_X1 \read_data[11]$_SDFFE_PN0P_  (.D(_076_),
    .CK(clknet_4_0_0_clk),
    .Q(net207),
    .QN(_437_));
 DFF_X1 \read_data[12]$_SDFFE_PN0P_  (.D(_077_),
    .CK(clknet_4_1_0_clk),
    .Q(net208),
    .QN(_436_));
 DFF_X1 \read_data[13]$_SDFFE_PN0P_  (.D(_078_),
    .CK(clknet_4_1_0_clk),
    .Q(net209),
    .QN(_435_));
 DFF_X1 \read_data[14]$_SDFFE_PN0P_  (.D(_079_),
    .CK(clknet_4_9_0_clk),
    .Q(net210),
    .QN(_434_));
 DFF_X1 \read_data[15]$_SDFFE_PN0P_  (.D(_080_),
    .CK(clknet_4_9_0_clk),
    .Q(net211),
    .QN(_433_));
 DFF_X1 \read_data[16]$_SDFFE_PN0P_  (.D(_081_),
    .CK(clknet_4_9_0_clk),
    .Q(net212),
    .QN(_432_));
 DFF_X1 \read_data[17]$_SDFFE_PN0P_  (.D(_082_),
    .CK(clknet_4_11_0_clk),
    .Q(net213),
    .QN(_431_));
 DFF_X1 \read_data[18]$_SDFFE_PN0P_  (.D(_083_),
    .CK(clknet_4_10_0_clk),
    .Q(net214),
    .QN(_430_));
 DFF_X1 \read_data[19]$_SDFFE_PN0P_  (.D(_084_),
    .CK(clknet_4_11_0_clk),
    .Q(net215),
    .QN(_429_));
 DFF_X1 \read_data[1]$_SDFFE_PN0P_  (.D(_085_),
    .CK(clknet_4_11_0_clk),
    .Q(net216),
    .QN(_428_));
 DFF_X1 \read_data[20]$_SDFFE_PN0P_  (.D(_086_),
    .CK(clknet_4_10_0_clk),
    .Q(net217),
    .QN(_427_));
 DFF_X1 \read_data[21]$_SDFFE_PN0P_  (.D(_087_),
    .CK(clknet_4_10_0_clk),
    .Q(net218),
    .QN(_426_));
 DFF_X1 \read_data[22]$_SDFFE_PN0P_  (.D(_088_),
    .CK(clknet_4_10_0_clk),
    .Q(net219),
    .QN(_425_));
 DFF_X1 \read_data[23]$_SDFFE_PN0P_  (.D(_089_),
    .CK(clknet_4_10_0_clk),
    .Q(net220),
    .QN(_424_));
 DFF_X1 \read_data[24]$_SDFFE_PN0P_  (.D(_090_),
    .CK(clknet_4_10_0_clk),
    .Q(net221),
    .QN(_423_));
 DFF_X1 \read_data[25]$_SDFFE_PN0P_  (.D(_091_),
    .CK(clknet_4_10_0_clk),
    .Q(net222),
    .QN(_422_));
 DFF_X1 \read_data[26]$_SDFFE_PN0P_  (.D(_092_),
    .CK(clknet_4_10_0_clk),
    .Q(net223),
    .QN(_421_));
 DFF_X1 \read_data[27]$_SDFFE_PN0P_  (.D(_093_),
    .CK(clknet_4_10_0_clk),
    .Q(net224),
    .QN(_420_));
 DFF_X1 \read_data[28]$_SDFFE_PN0P_  (.D(_094_),
    .CK(clknet_4_8_0_clk),
    .Q(net225),
    .QN(_419_));
 DFF_X1 \read_data[29]$_SDFFE_PN0P_  (.D(_095_),
    .CK(clknet_4_10_0_clk),
    .Q(net226),
    .QN(_418_));
 DFF_X1 \read_data[2]$_SDFFE_PN0P_  (.D(_096_),
    .CK(clknet_4_10_0_clk),
    .Q(net227),
    .QN(_417_));
 DFF_X1 \read_data[30]$_SDFFE_PN0P_  (.D(_097_),
    .CK(clknet_4_10_0_clk),
    .Q(net228),
    .QN(_416_));
 DFF_X1 \read_data[31]$_SDFFE_PN0P_  (.D(_098_),
    .CK(clknet_4_10_0_clk),
    .Q(net229),
    .QN(_415_));
 DFF_X1 \read_data[3]$_SDFFE_PN0P_  (.D(_099_),
    .CK(clknet_4_8_0_clk),
    .Q(net230),
    .QN(_414_));
 DFF_X1 \read_data[4]$_SDFFE_PN0P_  (.D(_100_),
    .CK(clknet_4_8_0_clk),
    .Q(net231),
    .QN(_413_));
 DFF_X1 \read_data[5]$_SDFFE_PN0P_  (.D(_101_),
    .CK(clknet_4_8_0_clk),
    .Q(net232),
    .QN(_412_));
 DFF_X1 \read_data[6]$_SDFFE_PN0P_  (.D(_102_),
    .CK(clknet_4_8_0_clk),
    .Q(net233),
    .QN(_411_));
 DFF_X1 \read_data[7]$_SDFFE_PN0P_  (.D(_103_),
    .CK(clknet_4_8_0_clk),
    .Q(net234),
    .QN(_410_));
 DFF_X1 \read_data[8]$_SDFFE_PN0P_  (.D(_104_),
    .CK(clknet_4_8_0_clk),
    .Q(net235),
    .QN(_409_));
 DFF_X1 \read_data[9]$_SDFFE_PN0P_  (.D(_105_),
    .CK(clknet_4_8_0_clk),
    .Q(net236),
    .QN(_408_));
 DFF_X1 \read_done_r$_SDFFE_PN0P_  (.D(_106_),
    .CK(clknet_4_9_0_clk),
    .Q(net237),
    .QN(_407_));
 DFF_X1 \rready$_SDFFE_PN0P_  (.D(_107_),
    .CK(clknet_4_9_0_clk),
    .Q(net238),
    .QN(_507_));
 DFF_X1 \state_r[0]$_DFF_P_  (.D(_000_),
    .CK(clknet_4_6_0_clk),
    .Q(\state_r[0] ),
    .QN(_508_));
 DFF_X1 \state_r[1]$_DFF_P_  (.D(_001_),
    .CK(clknet_4_11_0_clk),
    .Q(\state_r[1] ),
    .QN(_509_));
 DFF_X1 \state_r[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_4_12_0_clk),
    .Q(\state_r[2] ),
    .QN(_510_));
 DFF_X1 \state_r[3]$_DFF_P_  (.D(_003_),
    .CK(clknet_4_12_0_clk),
    .Q(\state_r[3] ),
    .QN(_511_));
 DFF_X1 \state_r[4]$_DFF_P_  (.D(_004_),
    .CK(clknet_4_12_0_clk),
    .Q(\state_r[4] ),
    .QN(_512_));
 DFF_X1 \state_r[5]$_DFF_P_  (.D(_005_),
    .CK(clknet_4_12_0_clk),
    .Q(\state_r[5] ),
    .QN(_006_));
 DFF_X1 \wdata[0]$_SDFFE_PN0P_  (.D(_108_),
    .CK(clknet_4_2_0_clk),
    .Q(net239),
    .QN(_406_));
 DFF_X1 \wdata[10]$_SDFFE_PN0P_  (.D(_109_),
    .CK(clknet_4_2_0_clk),
    .Q(net240),
    .QN(_405_));
 DFF_X1 \wdata[11]$_SDFFE_PN0P_  (.D(_110_),
    .CK(clknet_4_2_0_clk),
    .Q(net241),
    .QN(_404_));
 DFF_X1 \wdata[12]$_SDFFE_PN0P_  (.D(_111_),
    .CK(clknet_4_3_0_clk),
    .Q(net242),
    .QN(_403_));
 DFF_X1 \wdata[13]$_SDFFE_PN0P_  (.D(_112_),
    .CK(clknet_4_2_0_clk),
    .Q(net243),
    .QN(_402_));
 DFF_X1 \wdata[14]$_SDFFE_PN0P_  (.D(_113_),
    .CK(clknet_4_2_0_clk),
    .Q(net244),
    .QN(_401_));
 DFF_X1 \wdata[15]$_SDFFE_PN0P_  (.D(_114_),
    .CK(clknet_4_3_0_clk),
    .Q(net245),
    .QN(_400_));
 DFF_X1 \wdata[16]$_SDFFE_PN0P_  (.D(_115_),
    .CK(clknet_4_0_0_clk),
    .Q(net246),
    .QN(_399_));
 DFF_X1 \wdata[17]$_SDFFE_PN0P_  (.D(_116_),
    .CK(clknet_4_0_0_clk),
    .Q(net247),
    .QN(_398_));
 DFF_X1 \wdata[18]$_SDFFE_PN0P_  (.D(_117_),
    .CK(clknet_4_0_0_clk),
    .Q(net248),
    .QN(_397_));
 DFF_X1 \wdata[19]$_SDFFE_PN0P_  (.D(_118_),
    .CK(clknet_4_0_0_clk),
    .Q(net249),
    .QN(_396_));
 DFF_X1 \wdata[1]$_SDFFE_PN0P_  (.D(_119_),
    .CK(clknet_4_0_0_clk),
    .Q(net250),
    .QN(_395_));
 DFF_X1 \wdata[20]$_SDFFE_PN0P_  (.D(_120_),
    .CK(clknet_4_3_0_clk),
    .Q(net251),
    .QN(_394_));
 DFF_X1 \wdata[21]$_SDFFE_PN0P_  (.D(_121_),
    .CK(clknet_4_3_0_clk),
    .Q(net252),
    .QN(_393_));
 DFF_X1 \wdata[22]$_SDFFE_PN0P_  (.D(_122_),
    .CK(clknet_4_0_0_clk),
    .Q(net253),
    .QN(_392_));
 DFF_X1 \wdata[23]$_SDFFE_PN0P_  (.D(_123_),
    .CK(clknet_4_0_0_clk),
    .Q(net254),
    .QN(_391_));
 DFF_X1 \wdata[24]$_SDFFE_PN0P_  (.D(_124_),
    .CK(clknet_4_3_0_clk),
    .Q(net255),
    .QN(_390_));
 DFF_X1 \wdata[25]$_SDFFE_PN0P_  (.D(_125_),
    .CK(clknet_4_0_0_clk),
    .Q(net256),
    .QN(_389_));
 DFF_X1 \wdata[26]$_SDFFE_PN0P_  (.D(_126_),
    .CK(clknet_4_1_0_clk),
    .Q(net257),
    .QN(_388_));
 DFF_X1 \wdata[27]$_SDFFE_PN0P_  (.D(_127_),
    .CK(clknet_4_3_0_clk),
    .Q(net258),
    .QN(_387_));
 DFF_X1 \wdata[28]$_SDFFE_PN0P_  (.D(_128_),
    .CK(clknet_4_0_0_clk),
    .Q(net259),
    .QN(_386_));
 DFF_X1 \wdata[29]$_SDFFE_PN0P_  (.D(_129_),
    .CK(clknet_4_1_0_clk),
    .Q(net260),
    .QN(_385_));
 DFF_X1 \wdata[2]$_SDFFE_PN0P_  (.D(_130_),
    .CK(clknet_4_0_0_clk),
    .Q(net261),
    .QN(_384_));
 DFF_X1 \wdata[30]$_SDFFE_PN0P_  (.D(_131_),
    .CK(clknet_4_1_0_clk),
    .Q(net262),
    .QN(_383_));
 DFF_X1 \wdata[31]$_SDFFE_PN0P_  (.D(_132_),
    .CK(clknet_4_1_0_clk),
    .Q(net263),
    .QN(_382_));
 DFF_X1 \wdata[3]$_SDFFE_PN0P_  (.D(_133_),
    .CK(clknet_4_1_0_clk),
    .Q(net264),
    .QN(_381_));
 DFF_X1 \wdata[4]$_SDFFE_PN0P_  (.D(_134_),
    .CK(clknet_4_1_0_clk),
    .Q(net265),
    .QN(_380_));
 DFF_X1 \wdata[5]$_SDFFE_PN0P_  (.D(_135_),
    .CK(clknet_4_5_0_clk),
    .Q(net266),
    .QN(_379_));
 DFF_X1 \wdata[6]$_SDFFE_PN0P_  (.D(_136_),
    .CK(clknet_4_4_0_clk),
    .Q(net267),
    .QN(_378_));
 DFF_X1 \wdata[7]$_SDFFE_PN0P_  (.D(_137_),
    .CK(clknet_4_4_0_clk),
    .Q(net268),
    .QN(_377_));
 DFF_X1 \wdata[8]$_SDFFE_PN0P_  (.D(_138_),
    .CK(clknet_4_4_0_clk),
    .Q(net269),
    .QN(_376_));
 DFF_X1 \wdata[9]$_SDFFE_PN0P_  (.D(_139_),
    .CK(clknet_4_4_0_clk),
    .Q(net270),
    .QN(_375_));
 DFF_X1 \write_done_r$_SDFFE_PN0P_  (.D(_140_),
    .CK(clknet_4_6_0_clk),
    .Q(net271),
    .QN(_374_));
 DFF_X1 \wstrb[0]$_SDFFE_PN0P_  (.D(_141_),
    .CK(clknet_4_1_0_clk),
    .Q(net272),
    .QN(_373_));
 DFF_X1 \wstrb[1]$_SDFFE_PN0P_  (.D(_142_),
    .CK(clknet_4_6_0_clk),
    .Q(net273),
    .QN(_372_));
 DFF_X1 \wstrb[2]$_SDFFE_PN0P_  (.D(_143_),
    .CK(clknet_4_4_0_clk),
    .Q(net274),
    .QN(_371_));
 DFF_X1 \wstrb[3]$_SDFFE_PN0P_  (.D(_144_),
    .CK(clknet_4_7_0_clk),
    .Q(net275),
    .QN(_370_));
 DFF_X1 \wvalid$_SDFFE_PN0P_  (.D(_145_),
    .CK(clknet_4_14_0_clk),
    .Q(net276),
    .QN(_369_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_67 ();
 BUF_X1 input1 (.A(arready),
    .Z(net1));
 BUF_X1 input2 (.A(awready),
    .Z(net2));
 BUF_X1 input3 (.A(bvalid),
    .Z(net3));
 BUF_X1 input4 (.A(rdata[0]),
    .Z(net4));
 BUF_X1 input5 (.A(rdata[10]),
    .Z(net5));
 BUF_X1 input6 (.A(rdata[11]),
    .Z(net6));
 BUF_X1 input7 (.A(rdata[12]),
    .Z(net7));
 BUF_X1 input8 (.A(rdata[13]),
    .Z(net8));
 BUF_X1 input9 (.A(rdata[14]),
    .Z(net9));
 BUF_X1 input10 (.A(rdata[15]),
    .Z(net10));
 BUF_X1 input11 (.A(rdata[16]),
    .Z(net11));
 BUF_X1 input12 (.A(rdata[17]),
    .Z(net12));
 BUF_X1 input13 (.A(rdata[18]),
    .Z(net13));
 BUF_X1 input14 (.A(rdata[19]),
    .Z(net14));
 BUF_X1 input15 (.A(rdata[1]),
    .Z(net15));
 BUF_X1 input16 (.A(rdata[20]),
    .Z(net16));
 BUF_X1 input17 (.A(rdata[21]),
    .Z(net17));
 BUF_X1 input18 (.A(rdata[22]),
    .Z(net18));
 BUF_X1 input19 (.A(rdata[23]),
    .Z(net19));
 BUF_X1 input20 (.A(rdata[24]),
    .Z(net20));
 BUF_X1 input21 (.A(rdata[25]),
    .Z(net21));
 BUF_X1 input22 (.A(rdata[26]),
    .Z(net22));
 BUF_X1 input23 (.A(rdata[27]),
    .Z(net23));
 BUF_X1 input24 (.A(rdata[28]),
    .Z(net24));
 BUF_X1 input25 (.A(rdata[29]),
    .Z(net25));
 BUF_X1 input26 (.A(rdata[2]),
    .Z(net26));
 BUF_X1 input27 (.A(rdata[30]),
    .Z(net27));
 BUF_X1 input28 (.A(rdata[31]),
    .Z(net28));
 BUF_X1 input29 (.A(rdata[3]),
    .Z(net29));
 BUF_X1 input30 (.A(rdata[4]),
    .Z(net30));
 BUF_X1 input31 (.A(rdata[5]),
    .Z(net31));
 BUF_X1 input32 (.A(rdata[6]),
    .Z(net32));
 BUF_X1 input33 (.A(rdata[7]),
    .Z(net33));
 BUF_X1 input34 (.A(rdata[8]),
    .Z(net34));
 BUF_X1 input35 (.A(rdata[9]),
    .Z(net35));
 BUF_X1 input36 (.A(read_addr[0]),
    .Z(net36));
 BUF_X1 input37 (.A(read_addr[10]),
    .Z(net37));
 BUF_X1 input38 (.A(read_addr[11]),
    .Z(net38));
 BUF_X1 input39 (.A(read_addr[12]),
    .Z(net39));
 BUF_X1 input40 (.A(read_addr[13]),
    .Z(net40));
 BUF_X1 input41 (.A(read_addr[14]),
    .Z(net41));
 BUF_X1 input42 (.A(read_addr[15]),
    .Z(net42));
 BUF_X1 input43 (.A(read_addr[16]),
    .Z(net43));
 BUF_X1 input44 (.A(read_addr[17]),
    .Z(net44));
 BUF_X1 input45 (.A(read_addr[18]),
    .Z(net45));
 BUF_X1 input46 (.A(read_addr[19]),
    .Z(net46));
 BUF_X1 input47 (.A(read_addr[1]),
    .Z(net47));
 BUF_X1 input48 (.A(read_addr[20]),
    .Z(net48));
 BUF_X1 input49 (.A(read_addr[21]),
    .Z(net49));
 BUF_X1 input50 (.A(read_addr[22]),
    .Z(net50));
 BUF_X1 input51 (.A(read_addr[23]),
    .Z(net51));
 BUF_X1 input52 (.A(read_addr[24]),
    .Z(net52));
 BUF_X1 input53 (.A(read_addr[25]),
    .Z(net53));
 BUF_X1 input54 (.A(read_addr[26]),
    .Z(net54));
 BUF_X1 input55 (.A(read_addr[27]),
    .Z(net55));
 BUF_X1 input56 (.A(read_addr[28]),
    .Z(net56));
 BUF_X1 input57 (.A(read_addr[29]),
    .Z(net57));
 BUF_X1 input58 (.A(read_addr[2]),
    .Z(net58));
 BUF_X1 input59 (.A(read_addr[30]),
    .Z(net59));
 BUF_X1 input60 (.A(read_addr[31]),
    .Z(net60));
 BUF_X1 input61 (.A(read_addr[3]),
    .Z(net61));
 BUF_X1 input62 (.A(read_addr[4]),
    .Z(net62));
 BUF_X1 input63 (.A(read_addr[5]),
    .Z(net63));
 BUF_X1 input64 (.A(read_addr[6]),
    .Z(net64));
 BUF_X1 input65 (.A(read_addr[7]),
    .Z(net65));
 BUF_X1 input66 (.A(read_addr[8]),
    .Z(net66));
 BUF_X1 input67 (.A(read_addr[9]),
    .Z(net67));
 CLKBUF_X2 input68 (.A(rvalid),
    .Z(net68));
 BUF_X1 input69 (.A(wready),
    .Z(net69));
 BUF_X1 input70 (.A(write_addr[0]),
    .Z(net70));
 BUF_X1 input71 (.A(write_addr[10]),
    .Z(net71));
 BUF_X1 input72 (.A(write_addr[11]),
    .Z(net72));
 BUF_X1 input73 (.A(write_addr[12]),
    .Z(net73));
 BUF_X1 input74 (.A(write_addr[13]),
    .Z(net74));
 BUF_X1 input75 (.A(write_addr[14]),
    .Z(net75));
 BUF_X1 input76 (.A(write_addr[15]),
    .Z(net76));
 BUF_X1 input77 (.A(write_addr[16]),
    .Z(net77));
 BUF_X1 input78 (.A(write_addr[17]),
    .Z(net78));
 BUF_X1 input79 (.A(write_addr[18]),
    .Z(net79));
 BUF_X1 input80 (.A(write_addr[19]),
    .Z(net80));
 BUF_X1 input81 (.A(write_addr[1]),
    .Z(net81));
 BUF_X1 input82 (.A(write_addr[20]),
    .Z(net82));
 BUF_X1 input83 (.A(write_addr[21]),
    .Z(net83));
 BUF_X1 input84 (.A(write_addr[22]),
    .Z(net84));
 BUF_X1 input85 (.A(write_addr[23]),
    .Z(net85));
 BUF_X1 input86 (.A(write_addr[24]),
    .Z(net86));
 BUF_X1 input87 (.A(write_addr[25]),
    .Z(net87));
 BUF_X1 input88 (.A(write_addr[26]),
    .Z(net88));
 BUF_X1 input89 (.A(write_addr[27]),
    .Z(net89));
 BUF_X1 input90 (.A(write_addr[28]),
    .Z(net90));
 BUF_X1 input91 (.A(write_addr[29]),
    .Z(net91));
 BUF_X1 input92 (.A(write_addr[2]),
    .Z(net92));
 BUF_X1 input93 (.A(write_addr[30]),
    .Z(net93));
 BUF_X1 input94 (.A(write_addr[31]),
    .Z(net94));
 BUF_X1 input95 (.A(write_addr[3]),
    .Z(net95));
 BUF_X1 input96 (.A(write_addr[4]),
    .Z(net96));
 BUF_X1 input97 (.A(write_addr[5]),
    .Z(net97));
 BUF_X1 input98 (.A(write_addr[6]),
    .Z(net98));
 BUF_X1 input99 (.A(write_addr[7]),
    .Z(net99));
 BUF_X1 input100 (.A(write_addr[8]),
    .Z(net100));
 BUF_X1 input101 (.A(write_addr[9]),
    .Z(net101));
 BUF_X1 input102 (.A(write_data[0]),
    .Z(net102));
 BUF_X1 input103 (.A(write_data[10]),
    .Z(net103));
 BUF_X1 input104 (.A(write_data[11]),
    .Z(net104));
 BUF_X1 input105 (.A(write_data[12]),
    .Z(net105));
 BUF_X1 input106 (.A(write_data[13]),
    .Z(net106));
 BUF_X1 input107 (.A(write_data[14]),
    .Z(net107));
 BUF_X1 input108 (.A(write_data[15]),
    .Z(net108));
 BUF_X1 input109 (.A(write_data[16]),
    .Z(net109));
 BUF_X1 input110 (.A(write_data[17]),
    .Z(net110));
 BUF_X1 input111 (.A(write_data[18]),
    .Z(net111));
 BUF_X1 input112 (.A(write_data[19]),
    .Z(net112));
 BUF_X1 input113 (.A(write_data[1]),
    .Z(net113));
 BUF_X1 input114 (.A(write_data[20]),
    .Z(net114));
 BUF_X1 input115 (.A(write_data[21]),
    .Z(net115));
 BUF_X1 input116 (.A(write_data[22]),
    .Z(net116));
 BUF_X1 input117 (.A(write_data[23]),
    .Z(net117));
 BUF_X1 input118 (.A(write_data[24]),
    .Z(net118));
 BUF_X1 input119 (.A(write_data[25]),
    .Z(net119));
 BUF_X1 input120 (.A(write_data[26]),
    .Z(net120));
 BUF_X1 input121 (.A(write_data[27]),
    .Z(net121));
 BUF_X1 input122 (.A(write_data[28]),
    .Z(net122));
 BUF_X1 input123 (.A(write_data[29]),
    .Z(net123));
 BUF_X1 input124 (.A(write_data[2]),
    .Z(net124));
 BUF_X1 input125 (.A(write_data[30]),
    .Z(net125));
 BUF_X1 input126 (.A(write_data[31]),
    .Z(net126));
 BUF_X1 input127 (.A(write_data[3]),
    .Z(net127));
 BUF_X1 input128 (.A(write_data[4]),
    .Z(net128));
 BUF_X1 input129 (.A(write_data[5]),
    .Z(net129));
 BUF_X1 input130 (.A(write_data[6]),
    .Z(net130));
 BUF_X1 input131 (.A(write_data[7]),
    .Z(net131));
 BUF_X1 input132 (.A(write_data[8]),
    .Z(net132));
 BUF_X1 input133 (.A(write_data[9]),
    .Z(net133));
 BUF_X1 input134 (.A(write_strb[0]),
    .Z(net134));
 BUF_X1 input135 (.A(write_strb[1]),
    .Z(net135));
 BUF_X1 input136 (.A(write_strb[2]),
    .Z(net136));
 BUF_X1 input137 (.A(write_strb[3]),
    .Z(net137));
 BUF_X1 output138 (.A(net138),
    .Z(araddr[0]));
 BUF_X1 output139 (.A(net139),
    .Z(araddr[10]));
 BUF_X1 output140 (.A(net140),
    .Z(araddr[11]));
 BUF_X1 output141 (.A(net141),
    .Z(araddr[12]));
 BUF_X1 output142 (.A(net142),
    .Z(araddr[13]));
 BUF_X1 output143 (.A(net143),
    .Z(araddr[14]));
 BUF_X1 output144 (.A(net144),
    .Z(araddr[15]));
 BUF_X1 output145 (.A(net145),
    .Z(araddr[16]));
 BUF_X1 output146 (.A(net146),
    .Z(araddr[17]));
 BUF_X1 output147 (.A(net147),
    .Z(araddr[18]));
 BUF_X1 output148 (.A(net148),
    .Z(araddr[19]));
 BUF_X1 output149 (.A(net149),
    .Z(araddr[1]));
 BUF_X1 output150 (.A(net150),
    .Z(araddr[20]));
 BUF_X1 output151 (.A(net151),
    .Z(araddr[21]));
 BUF_X1 output152 (.A(net152),
    .Z(araddr[22]));
 BUF_X1 output153 (.A(net153),
    .Z(araddr[23]));
 BUF_X1 output154 (.A(net154),
    .Z(araddr[24]));
 BUF_X1 output155 (.A(net155),
    .Z(araddr[25]));
 BUF_X1 output156 (.A(net156),
    .Z(araddr[26]));
 BUF_X1 output157 (.A(net157),
    .Z(araddr[27]));
 BUF_X1 output158 (.A(net158),
    .Z(araddr[28]));
 BUF_X1 output159 (.A(net159),
    .Z(araddr[29]));
 BUF_X1 output160 (.A(net160),
    .Z(araddr[2]));
 BUF_X1 output161 (.A(net161),
    .Z(araddr[30]));
 BUF_X1 output162 (.A(net162),
    .Z(araddr[31]));
 BUF_X1 output163 (.A(net163),
    .Z(araddr[3]));
 BUF_X1 output164 (.A(net164),
    .Z(araddr[4]));
 BUF_X1 output165 (.A(net165),
    .Z(araddr[5]));
 BUF_X1 output166 (.A(net166),
    .Z(araddr[6]));
 BUF_X1 output167 (.A(net167),
    .Z(araddr[7]));
 BUF_X1 output168 (.A(net168),
    .Z(araddr[8]));
 BUF_X1 output169 (.A(net169),
    .Z(araddr[9]));
 BUF_X1 output170 (.A(net170),
    .Z(arvalid));
 BUF_X1 output171 (.A(net171),
    .Z(awaddr[0]));
 BUF_X1 output172 (.A(net172),
    .Z(awaddr[10]));
 BUF_X1 output173 (.A(net173),
    .Z(awaddr[11]));
 BUF_X1 output174 (.A(net174),
    .Z(awaddr[12]));
 BUF_X1 output175 (.A(net175),
    .Z(awaddr[13]));
 BUF_X1 output176 (.A(net176),
    .Z(awaddr[14]));
 BUF_X1 output177 (.A(net177),
    .Z(awaddr[15]));
 BUF_X1 output178 (.A(net178),
    .Z(awaddr[16]));
 BUF_X1 output179 (.A(net179),
    .Z(awaddr[17]));
 BUF_X1 output180 (.A(net180),
    .Z(awaddr[18]));
 BUF_X1 output181 (.A(net181),
    .Z(awaddr[19]));
 BUF_X1 output182 (.A(net182),
    .Z(awaddr[1]));
 BUF_X1 output183 (.A(net183),
    .Z(awaddr[20]));
 BUF_X1 output184 (.A(net184),
    .Z(awaddr[21]));
 BUF_X1 output185 (.A(net185),
    .Z(awaddr[22]));
 BUF_X1 output186 (.A(net186),
    .Z(awaddr[23]));
 BUF_X1 output187 (.A(net187),
    .Z(awaddr[24]));
 BUF_X1 output188 (.A(net188),
    .Z(awaddr[25]));
 BUF_X1 output189 (.A(net189),
    .Z(awaddr[26]));
 BUF_X1 output190 (.A(net190),
    .Z(awaddr[27]));
 BUF_X1 output191 (.A(net191),
    .Z(awaddr[28]));
 BUF_X1 output192 (.A(net192),
    .Z(awaddr[29]));
 BUF_X1 output193 (.A(net193),
    .Z(awaddr[2]));
 BUF_X1 output194 (.A(net194),
    .Z(awaddr[30]));
 BUF_X1 output195 (.A(net195),
    .Z(awaddr[31]));
 BUF_X1 output196 (.A(net196),
    .Z(awaddr[3]));
 BUF_X1 output197 (.A(net197),
    .Z(awaddr[4]));
 BUF_X1 output198 (.A(net198),
    .Z(awaddr[5]));
 BUF_X1 output199 (.A(net199),
    .Z(awaddr[6]));
 BUF_X1 output200 (.A(net200),
    .Z(awaddr[7]));
 BUF_X1 output201 (.A(net201),
    .Z(awaddr[8]));
 BUF_X1 output202 (.A(net202),
    .Z(awaddr[9]));
 BUF_X1 output203 (.A(net203),
    .Z(awvalid));
 BUF_X1 output204 (.A(net204),
    .Z(bready));
 BUF_X1 output205 (.A(net205),
    .Z(read_data[0]));
 BUF_X1 output206 (.A(net206),
    .Z(read_data[10]));
 BUF_X1 output207 (.A(net207),
    .Z(read_data[11]));
 BUF_X1 output208 (.A(net208),
    .Z(read_data[12]));
 BUF_X1 output209 (.A(net209),
    .Z(read_data[13]));
 BUF_X1 output210 (.A(net210),
    .Z(read_data[14]));
 BUF_X1 output211 (.A(net211),
    .Z(read_data[15]));
 BUF_X1 output212 (.A(net212),
    .Z(read_data[16]));
 BUF_X1 output213 (.A(net213),
    .Z(read_data[17]));
 BUF_X1 output214 (.A(net214),
    .Z(read_data[18]));
 BUF_X1 output215 (.A(net215),
    .Z(read_data[19]));
 BUF_X1 output216 (.A(net216),
    .Z(read_data[1]));
 BUF_X1 output217 (.A(net217),
    .Z(read_data[20]));
 BUF_X1 output218 (.A(net218),
    .Z(read_data[21]));
 BUF_X1 output219 (.A(net219),
    .Z(read_data[22]));
 BUF_X1 output220 (.A(net220),
    .Z(read_data[23]));
 BUF_X1 output221 (.A(net221),
    .Z(read_data[24]));
 BUF_X1 output222 (.A(net222),
    .Z(read_data[25]));
 BUF_X1 output223 (.A(net223),
    .Z(read_data[26]));
 BUF_X1 output224 (.A(net224),
    .Z(read_data[27]));
 BUF_X1 output225 (.A(net225),
    .Z(read_data[28]));
 BUF_X1 output226 (.A(net226),
    .Z(read_data[29]));
 BUF_X1 output227 (.A(net227),
    .Z(read_data[2]));
 BUF_X1 output228 (.A(net228),
    .Z(read_data[30]));
 BUF_X1 output229 (.A(net229),
    .Z(read_data[31]));
 BUF_X1 output230 (.A(net230),
    .Z(read_data[3]));
 BUF_X1 output231 (.A(net231),
    .Z(read_data[4]));
 BUF_X1 output232 (.A(net232),
    .Z(read_data[5]));
 BUF_X1 output233 (.A(net233),
    .Z(read_data[6]));
 BUF_X1 output234 (.A(net234),
    .Z(read_data[7]));
 BUF_X1 output235 (.A(net235),
    .Z(read_data[8]));
 BUF_X1 output236 (.A(net236),
    .Z(read_data[9]));
 BUF_X1 output237 (.A(net237),
    .Z(read_done));
 BUF_X1 output238 (.A(net238),
    .Z(rready));
 BUF_X1 output239 (.A(net239),
    .Z(wdata[0]));
 BUF_X1 output240 (.A(net240),
    .Z(wdata[10]));
 BUF_X1 output241 (.A(net241),
    .Z(wdata[11]));
 BUF_X1 output242 (.A(net242),
    .Z(wdata[12]));
 BUF_X1 output243 (.A(net243),
    .Z(wdata[13]));
 BUF_X1 output244 (.A(net244),
    .Z(wdata[14]));
 BUF_X1 output245 (.A(net245),
    .Z(wdata[15]));
 BUF_X1 output246 (.A(net246),
    .Z(wdata[16]));
 BUF_X1 output247 (.A(net247),
    .Z(wdata[17]));
 BUF_X1 output248 (.A(net248),
    .Z(wdata[18]));
 BUF_X1 output249 (.A(net249),
    .Z(wdata[19]));
 BUF_X1 output250 (.A(net250),
    .Z(wdata[1]));
 BUF_X1 output251 (.A(net251),
    .Z(wdata[20]));
 BUF_X1 output252 (.A(net252),
    .Z(wdata[21]));
 BUF_X1 output253 (.A(net253),
    .Z(wdata[22]));
 BUF_X1 output254 (.A(net254),
    .Z(wdata[23]));
 BUF_X1 output255 (.A(net255),
    .Z(wdata[24]));
 BUF_X1 output256 (.A(net256),
    .Z(wdata[25]));
 BUF_X1 output257 (.A(net257),
    .Z(wdata[26]));
 BUF_X1 output258 (.A(net258),
    .Z(wdata[27]));
 BUF_X1 output259 (.A(net259),
    .Z(wdata[28]));
 BUF_X1 output260 (.A(net260),
    .Z(wdata[29]));
 BUF_X1 output261 (.A(net261),
    .Z(wdata[2]));
 BUF_X1 output262 (.A(net262),
    .Z(wdata[30]));
 BUF_X1 output263 (.A(net263),
    .Z(wdata[31]));
 BUF_X1 output264 (.A(net264),
    .Z(wdata[3]));
 BUF_X1 output265 (.A(net265),
    .Z(wdata[4]));
 BUF_X1 output266 (.A(net266),
    .Z(wdata[5]));
 BUF_X1 output267 (.A(net267),
    .Z(wdata[6]));
 BUF_X1 output268 (.A(net268),
    .Z(wdata[7]));
 BUF_X1 output269 (.A(net269),
    .Z(wdata[8]));
 BUF_X1 output270 (.A(net270),
    .Z(wdata[9]));
 BUF_X1 output271 (.A(net271),
    .Z(write_done));
 BUF_X1 output272 (.A(net272),
    .Z(wstrb[0]));
 BUF_X1 output273 (.A(net273),
    .Z(wstrb[1]));
 BUF_X1 output274 (.A(net274),
    .Z(wstrb[2]));
 BUF_X1 output275 (.A(net275),
    .Z(wstrb[3]));
 BUF_X1 output276 (.A(net276),
    .Z(wvalid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 CLKBUF_X1 clkload0 (.A(clknet_4_0_0_clk));
 INV_X2 clkload1 (.A(clknet_4_1_0_clk));
 INV_X4 clkload2 (.A(clknet_4_2_0_clk));
 INV_X2 clkload3 (.A(clknet_4_3_0_clk));
 INV_X2 clkload4 (.A(clknet_4_4_0_clk));
 INV_X4 clkload5 (.A(clknet_4_6_0_clk));
 INV_X2 clkload6 (.A(clknet_4_7_0_clk));
 INV_X2 clkload7 (.A(clknet_4_8_0_clk));
 INV_X4 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_11_0_clk));
 INV_X4 clkload10 (.A(clknet_4_12_0_clk));
 INV_X2 clkload11 (.A(clknet_4_13_0_clk));
 INV_X2 clkload12 (.A(clknet_4_14_0_clk));
 FILLCELL_X2 FILLER_0_1 ();
 FILLCELL_X1 FILLER_0_30 ();
 FILLCELL_X2 FILLER_0_60 ();
 FILLCELL_X1 FILLER_0_65 ();
 FILLCELL_X1 FILLER_0_86 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_113 ();
 FILLCELL_X1 FILLER_0_157 ();
 FILLCELL_X1 FILLER_0_161 ();
 FILLCELL_X2 FILLER_0_195 ();
 FILLCELL_X2 FILLER_0_233 ();
 FILLCELL_X2 FILLER_0_249 ();
 FILLCELL_X1 FILLER_0_251 ();
 FILLCELL_X1 FILLER_1_22 ();
 FILLCELL_X2 FILLER_1_113 ();
 FILLCELL_X1 FILLER_1_126 ();
 FILLCELL_X1 FILLER_1_147 ();
 FILLCELL_X1 FILLER_1_155 ();
 FILLCELL_X1 FILLER_1_163 ();
 FILLCELL_X1 FILLER_1_181 ();
 FILLCELL_X1 FILLER_1_199 ();
 FILLCELL_X1 FILLER_1_204 ();
 FILLCELL_X2 FILLER_1_250 ();
 FILLCELL_X4 FILLER_2_1 ();
 FILLCELL_X2 FILLER_2_80 ();
 FILLCELL_X1 FILLER_2_110 ();
 FILLCELL_X4 FILLER_2_128 ();
 FILLCELL_X1 FILLER_2_132 ();
 FILLCELL_X1 FILLER_2_137 ();
 FILLCELL_X1 FILLER_2_166 ();
 FILLCELL_X1 FILLER_2_191 ();
 FILLCELL_X2 FILLER_2_222 ();
 FILLCELL_X1 FILLER_2_227 ();
 FILLCELL_X2 FILLER_2_231 ();
 FILLCELL_X2 FILLER_2_250 ();
 FILLCELL_X1 FILLER_3_14 ();
 FILLCELL_X1 FILLER_3_25 ();
 FILLCELL_X4 FILLER_3_29 ();
 FILLCELL_X1 FILLER_3_97 ();
 FILLCELL_X8 FILLER_3_104 ();
 FILLCELL_X4 FILLER_3_112 ();
 FILLCELL_X2 FILLER_3_116 ();
 FILLCELL_X8 FILLER_3_125 ();
 FILLCELL_X2 FILLER_3_133 ();
 FILLCELL_X1 FILLER_3_135 ();
 FILLCELL_X4 FILLER_3_153 ();
 FILLCELL_X2 FILLER_3_157 ();
 FILLCELL_X1 FILLER_3_159 ();
 FILLCELL_X2 FILLER_3_173 ();
 FILLCELL_X4 FILLER_3_195 ();
 FILLCELL_X2 FILLER_3_199 ();
 FILLCELL_X1 FILLER_3_201 ();
 FILLCELL_X16 FILLER_3_205 ();
 FILLCELL_X4 FILLER_3_221 ();
 FILLCELL_X1 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_243 ();
 FILLCELL_X2 FILLER_3_247 ();
 FILLCELL_X2 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_20 ();
 FILLCELL_X8 FILLER_4_31 ();
 FILLCELL_X4 FILLER_4_39 ();
 FILLCELL_X2 FILLER_4_43 ();
 FILLCELL_X8 FILLER_4_48 ();
 FILLCELL_X2 FILLER_4_56 ();
 FILLCELL_X1 FILLER_4_58 ();
 FILLCELL_X32 FILLER_4_66 ();
 FILLCELL_X4 FILLER_4_98 ();
 FILLCELL_X1 FILLER_4_102 ();
 FILLCELL_X8 FILLER_4_110 ();
 FILLCELL_X2 FILLER_4_118 ();
 FILLCELL_X32 FILLER_4_124 ();
 FILLCELL_X4 FILLER_4_156 ();
 FILLCELL_X2 FILLER_4_160 ();
 FILLCELL_X4 FILLER_4_172 ();
 FILLCELL_X1 FILLER_4_176 ();
 FILLCELL_X8 FILLER_4_182 ();
 FILLCELL_X8 FILLER_4_211 ();
 FILLCELL_X4 FILLER_4_219 ();
 FILLCELL_X1 FILLER_4_223 ();
 FILLCELL_X4 FILLER_4_227 ();
 FILLCELL_X1 FILLER_4_231 ();
 FILLCELL_X1 FILLER_4_248 ();
 FILLCELL_X1 FILLER_5_7 ();
 FILLCELL_X1 FILLER_5_36 ();
 FILLCELL_X4 FILLER_5_61 ();
 FILLCELL_X2 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_67 ();
 FILLCELL_X2 FILLER_5_92 ();
 FILLCELL_X1 FILLER_5_94 ();
 FILLCELL_X16 FILLER_5_99 ();
 FILLCELL_X8 FILLER_5_136 ();
 FILLCELL_X4 FILLER_5_144 ();
 FILLCELL_X1 FILLER_5_165 ();
 FILLCELL_X8 FILLER_5_185 ();
 FILLCELL_X8 FILLER_5_217 ();
 FILLCELL_X1 FILLER_5_225 ();
 FILLCELL_X2 FILLER_5_247 ();
 FILLCELL_X1 FILLER_6_21 ();
 FILLCELL_X1 FILLER_6_25 ();
 FILLCELL_X4 FILLER_6_33 ();
 FILLCELL_X1 FILLER_6_37 ();
 FILLCELL_X16 FILLER_6_42 ();
 FILLCELL_X4 FILLER_6_66 ();
 FILLCELL_X2 FILLER_6_70 ();
 FILLCELL_X8 FILLER_6_76 ();
 FILLCELL_X1 FILLER_6_84 ();
 FILLCELL_X4 FILLER_6_109 ();
 FILLCELL_X2 FILLER_6_113 ();
 FILLCELL_X16 FILLER_6_126 ();
 FILLCELL_X1 FILLER_6_142 ();
 FILLCELL_X8 FILLER_6_154 ();
 FILLCELL_X4 FILLER_6_162 ();
 FILLCELL_X2 FILLER_6_166 ();
 FILLCELL_X4 FILLER_6_172 ();
 FILLCELL_X2 FILLER_6_176 ();
 FILLCELL_X2 FILLER_6_195 ();
 FILLCELL_X4 FILLER_6_201 ();
 FILLCELL_X2 FILLER_6_205 ();
 FILLCELL_X1 FILLER_6_207 ();
 FILLCELL_X4 FILLER_6_212 ();
 FILLCELL_X2 FILLER_6_216 ();
 FILLCELL_X1 FILLER_6_218 ();
 FILLCELL_X2 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_6 ();
 FILLCELL_X2 FILLER_7_24 ();
 FILLCELL_X2 FILLER_7_33 ();
 FILLCELL_X1 FILLER_7_35 ();
 FILLCELL_X2 FILLER_7_40 ();
 FILLCELL_X1 FILLER_7_42 ();
 FILLCELL_X2 FILLER_7_60 ();
 FILLCELL_X1 FILLER_7_79 ();
 FILLCELL_X4 FILLER_7_87 ();
 FILLCELL_X1 FILLER_7_91 ();
 FILLCELL_X16 FILLER_7_96 ();
 FILLCELL_X2 FILLER_7_112 ();
 FILLCELL_X4 FILLER_7_131 ();
 FILLCELL_X1 FILLER_7_135 ();
 FILLCELL_X1 FILLER_7_160 ();
 FILLCELL_X16 FILLER_7_178 ();
 FILLCELL_X2 FILLER_7_236 ();
 FILLCELL_X1 FILLER_8_4 ();
 FILLCELL_X1 FILLER_8_12 ();
 FILLCELL_X1 FILLER_8_34 ();
 FILLCELL_X4 FILLER_8_52 ();
 FILLCELL_X1 FILLER_8_56 ();
 FILLCELL_X4 FILLER_8_61 ();
 FILLCELL_X16 FILLER_8_107 ();
 FILLCELL_X8 FILLER_8_123 ();
 FILLCELL_X4 FILLER_8_131 ();
 FILLCELL_X2 FILLER_8_135 ();
 FILLCELL_X2 FILLER_8_181 ();
 FILLCELL_X1 FILLER_8_183 ();
 FILLCELL_X8 FILLER_8_189 ();
 FILLCELL_X2 FILLER_8_197 ();
 FILLCELL_X1 FILLER_8_199 ();
 FILLCELL_X8 FILLER_8_204 ();
 FILLCELL_X2 FILLER_8_212 ();
 FILLCELL_X1 FILLER_8_214 ();
 FILLCELL_X4 FILLER_8_245 ();
 FILLCELL_X1 FILLER_9_18 ();
 FILLCELL_X2 FILLER_9_22 ();
 FILLCELL_X1 FILLER_9_28 ();
 FILLCELL_X1 FILLER_9_32 ();
 FILLCELL_X2 FILLER_9_54 ();
 FILLCELL_X1 FILLER_9_56 ();
 FILLCELL_X16 FILLER_9_62 ();
 FILLCELL_X8 FILLER_9_82 ();
 FILLCELL_X4 FILLER_9_95 ();
 FILLCELL_X1 FILLER_9_99 ();
 FILLCELL_X32 FILLER_9_110 ();
 FILLCELL_X8 FILLER_9_142 ();
 FILLCELL_X2 FILLER_9_150 ();
 FILLCELL_X2 FILLER_9_156 ();
 FILLCELL_X1 FILLER_9_158 ();
 FILLCELL_X16 FILLER_9_172 ();
 FILLCELL_X8 FILLER_9_188 ();
 FILLCELL_X2 FILLER_9_196 ();
 FILLCELL_X2 FILLER_9_222 ();
 FILLCELL_X1 FILLER_9_224 ();
 FILLCELL_X2 FILLER_9_231 ();
 FILLCELL_X2 FILLER_9_243 ();
 FILLCELL_X1 FILLER_9_245 ();
 FILLCELL_X1 FILLER_10_42 ();
 FILLCELL_X32 FILLER_10_59 ();
 FILLCELL_X32 FILLER_10_91 ();
 FILLCELL_X16 FILLER_10_123 ();
 FILLCELL_X8 FILLER_10_139 ();
 FILLCELL_X32 FILLER_10_157 ();
 FILLCELL_X16 FILLER_10_189 ();
 FILLCELL_X8 FILLER_10_205 ();
 FILLCELL_X4 FILLER_10_222 ();
 FILLCELL_X1 FILLER_10_226 ();
 FILLCELL_X1 FILLER_10_248 ();
 FILLCELL_X2 FILLER_11_7 ();
 FILLCELL_X8 FILLER_11_12 ();
 FILLCELL_X1 FILLER_11_20 ();
 FILLCELL_X32 FILLER_11_63 ();
 FILLCELL_X32 FILLER_11_95 ();
 FILLCELL_X8 FILLER_11_127 ();
 FILLCELL_X4 FILLER_11_135 ();
 FILLCELL_X2 FILLER_11_139 ();
 FILLCELL_X1 FILLER_11_141 ();
 FILLCELL_X32 FILLER_11_149 ();
 FILLCELL_X16 FILLER_11_181 ();
 FILLCELL_X4 FILLER_11_197 ();
 FILLCELL_X1 FILLER_11_244 ();
 FILLCELL_X1 FILLER_12_7 ();
 FILLCELL_X2 FILLER_12_11 ();
 FILLCELL_X1 FILLER_12_37 ();
 FILLCELL_X32 FILLER_12_54 ();
 FILLCELL_X32 FILLER_12_86 ();
 FILLCELL_X32 FILLER_12_118 ();
 FILLCELL_X32 FILLER_12_150 ();
 FILLCELL_X16 FILLER_12_182 ();
 FILLCELL_X8 FILLER_12_198 ();
 FILLCELL_X4 FILLER_12_206 ();
 FILLCELL_X2 FILLER_12_210 ();
 FILLCELL_X1 FILLER_12_212 ();
 FILLCELL_X2 FILLER_12_216 ();
 FILLCELL_X1 FILLER_12_241 ();
 FILLCELL_X1 FILLER_12_245 ();
 FILLCELL_X2 FILLER_13_4 ();
 FILLCELL_X1 FILLER_13_28 ();
 FILLCELL_X32 FILLER_13_63 ();
 FILLCELL_X32 FILLER_13_95 ();
 FILLCELL_X32 FILLER_13_127 ();
 FILLCELL_X8 FILLER_13_159 ();
 FILLCELL_X4 FILLER_13_167 ();
 FILLCELL_X1 FILLER_13_171 ();
 FILLCELL_X16 FILLER_13_189 ();
 FILLCELL_X8 FILLER_13_205 ();
 FILLCELL_X2 FILLER_13_216 ();
 FILLCELL_X1 FILLER_13_218 ();
 FILLCELL_X2 FILLER_13_226 ();
 FILLCELL_X1 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_5 ();
 FILLCELL_X2 FILLER_14_46 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X8 FILLER_14_113 ();
 FILLCELL_X2 FILLER_14_121 ();
 FILLCELL_X8 FILLER_14_157 ();
 FILLCELL_X2 FILLER_14_165 ();
 FILLCELL_X16 FILLER_14_190 ();
 FILLCELL_X1 FILLER_14_206 ();
 FILLCELL_X2 FILLER_14_218 ();
 FILLCELL_X1 FILLER_14_220 ();
 FILLCELL_X1 FILLER_14_228 ();
 FILLCELL_X1 FILLER_14_233 ();
 FILLCELL_X1 FILLER_14_238 ();
 FILLCELL_X2 FILLER_14_243 ();
 FILLCELL_X1 FILLER_14_248 ();
 FILLCELL_X2 FILLER_15_21 ();
 FILLCELL_X1 FILLER_15_30 ();
 FILLCELL_X2 FILLER_15_35 ();
 FILLCELL_X2 FILLER_15_40 ();
 FILLCELL_X2 FILLER_15_49 ();
 FILLCELL_X1 FILLER_15_51 ();
 FILLCELL_X32 FILLER_15_56 ();
 FILLCELL_X32 FILLER_15_88 ();
 FILLCELL_X8 FILLER_15_120 ();
 FILLCELL_X4 FILLER_15_128 ();
 FILLCELL_X2 FILLER_15_136 ();
 FILLCELL_X2 FILLER_15_142 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X1 FILLER_15_151 ();
 FILLCELL_X1 FILLER_15_154 ();
 FILLCELL_X2 FILLER_15_162 ();
 FILLCELL_X1 FILLER_15_164 ();
 FILLCELL_X1 FILLER_15_179 ();
 FILLCELL_X4 FILLER_15_200 ();
 FILLCELL_X1 FILLER_15_204 ();
 FILLCELL_X2 FILLER_15_225 ();
 FILLCELL_X1 FILLER_15_227 ();
 FILLCELL_X1 FILLER_16_4 ();
 FILLCELL_X16 FILLER_16_22 ();
 FILLCELL_X8 FILLER_16_38 ();
 FILLCELL_X4 FILLER_16_46 ();
 FILLCELL_X2 FILLER_16_50 ();
 FILLCELL_X32 FILLER_16_56 ();
 FILLCELL_X32 FILLER_16_88 ();
 FILLCELL_X16 FILLER_16_120 ();
 FILLCELL_X8 FILLER_16_136 ();
 FILLCELL_X1 FILLER_16_144 ();
 FILLCELL_X1 FILLER_16_171 ();
 FILLCELL_X4 FILLER_16_176 ();
 FILLCELL_X2 FILLER_16_180 ();
 FILLCELL_X16 FILLER_16_189 ();
 FILLCELL_X8 FILLER_16_205 ();
 FILLCELL_X1 FILLER_16_213 ();
 FILLCELL_X2 FILLER_16_225 ();
 FILLCELL_X2 FILLER_16_240 ();
 FILLCELL_X2 FILLER_17_7 ();
 FILLCELL_X1 FILLER_17_9 ();
 FILLCELL_X32 FILLER_17_42 ();
 FILLCELL_X8 FILLER_17_74 ();
 FILLCELL_X2 FILLER_17_82 ();
 FILLCELL_X16 FILLER_17_89 ();
 FILLCELL_X8 FILLER_17_105 ();
 FILLCELL_X4 FILLER_17_113 ();
 FILLCELL_X2 FILLER_17_117 ();
 FILLCELL_X2 FILLER_17_124 ();
 FILLCELL_X2 FILLER_17_140 ();
 FILLCELL_X2 FILLER_17_160 ();
 FILLCELL_X8 FILLER_17_167 ();
 FILLCELL_X8 FILLER_17_186 ();
 FILLCELL_X4 FILLER_17_194 ();
 FILLCELL_X2 FILLER_17_215 ();
 FILLCELL_X1 FILLER_17_217 ();
 FILLCELL_X2 FILLER_17_222 ();
 FILLCELL_X1 FILLER_17_224 ();
 FILLCELL_X4 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_32 ();
 FILLCELL_X4 FILLER_18_50 ();
 FILLCELL_X1 FILLER_18_54 ();
 FILLCELL_X4 FILLER_18_60 ();
 FILLCELL_X2 FILLER_18_64 ();
 FILLCELL_X1 FILLER_18_66 ();
 FILLCELL_X32 FILLER_18_71 ();
 FILLCELL_X8 FILLER_18_103 ();
 FILLCELL_X2 FILLER_18_128 ();
 FILLCELL_X8 FILLER_18_137 ();
 FILLCELL_X1 FILLER_18_145 ();
 FILLCELL_X1 FILLER_18_163 ();
 FILLCELL_X4 FILLER_18_179 ();
 FILLCELL_X1 FILLER_18_183 ();
 FILLCELL_X16 FILLER_18_188 ();
 FILLCELL_X4 FILLER_18_204 ();
 FILLCELL_X4 FILLER_18_225 ();
 FILLCELL_X2 FILLER_18_229 ();
 FILLCELL_X1 FILLER_18_231 ();
 FILLCELL_X16 FILLER_18_236 ();
 FILLCELL_X2 FILLER_19_30 ();
 FILLCELL_X4 FILLER_19_36 ();
 FILLCELL_X2 FILLER_19_40 ();
 FILLCELL_X1 FILLER_19_46 ();
 FILLCELL_X1 FILLER_19_64 ();
 FILLCELL_X8 FILLER_19_70 ();
 FILLCELL_X2 FILLER_19_78 ();
 FILLCELL_X32 FILLER_19_87 ();
 FILLCELL_X16 FILLER_19_119 ();
 FILLCELL_X4 FILLER_19_135 ();
 FILLCELL_X2 FILLER_19_139 ();
 FILLCELL_X8 FILLER_19_143 ();
 FILLCELL_X2 FILLER_19_151 ();
 FILLCELL_X1 FILLER_19_153 ();
 FILLCELL_X2 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_184 ();
 FILLCELL_X2 FILLER_19_188 ();
 FILLCELL_X16 FILLER_19_207 ();
 FILLCELL_X1 FILLER_19_223 ();
 FILLCELL_X2 FILLER_20_22 ();
 FILLCELL_X2 FILLER_20_35 ();
 FILLCELL_X4 FILLER_20_44 ();
 FILLCELL_X2 FILLER_20_48 ();
 FILLCELL_X32 FILLER_20_71 ();
 FILLCELL_X16 FILLER_20_103 ();
 FILLCELL_X8 FILLER_20_119 ();
 FILLCELL_X1 FILLER_20_127 ();
 FILLCELL_X1 FILLER_20_131 ();
 FILLCELL_X4 FILLER_20_135 ();
 FILLCELL_X2 FILLER_20_139 ();
 FILLCELL_X4 FILLER_20_146 ();
 FILLCELL_X4 FILLER_20_159 ();
 FILLCELL_X1 FILLER_20_163 ();
 FILLCELL_X2 FILLER_20_179 ();
 FILLCELL_X1 FILLER_20_181 ();
 FILLCELL_X4 FILLER_20_189 ();
 FILLCELL_X2 FILLER_20_193 ();
 FILLCELL_X1 FILLER_20_195 ();
 FILLCELL_X16 FILLER_20_201 ();
 FILLCELL_X2 FILLER_20_220 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_22 ();
 FILLCELL_X8 FILLER_21_28 ();
 FILLCELL_X2 FILLER_21_36 ();
 FILLCELL_X1 FILLER_21_38 ();
 FILLCELL_X1 FILLER_21_42 ();
 FILLCELL_X32 FILLER_21_67 ();
 FILLCELL_X16 FILLER_21_99 ();
 FILLCELL_X8 FILLER_21_115 ();
 FILLCELL_X1 FILLER_21_140 ();
 FILLCELL_X1 FILLER_21_177 ();
 FILLCELL_X16 FILLER_21_185 ();
 FILLCELL_X8 FILLER_21_201 ();
 FILLCELL_X4 FILLER_21_209 ();
 FILLCELL_X1 FILLER_21_213 ();
 FILLCELL_X4 FILLER_21_217 ();
 FILLCELL_X2 FILLER_21_221 ();
 FILLCELL_X2 FILLER_21_237 ();
 FILLCELL_X1 FILLER_21_239 ();
 FILLCELL_X1 FILLER_21_243 ();
 FILLCELL_X2 FILLER_21_247 ();
 FILLCELL_X2 FILLER_22_7 ();
 FILLCELL_X1 FILLER_22_13 ();
 FILLCELL_X2 FILLER_22_34 ();
 FILLCELL_X32 FILLER_22_53 ();
 FILLCELL_X32 FILLER_22_85 ();
 FILLCELL_X4 FILLER_22_117 ();
 FILLCELL_X1 FILLER_22_121 ();
 FILLCELL_X2 FILLER_22_126 ();
 FILLCELL_X1 FILLER_22_128 ();
 FILLCELL_X1 FILLER_22_133 ();
 FILLCELL_X8 FILLER_22_138 ();
 FILLCELL_X1 FILLER_22_146 ();
 FILLCELL_X8 FILLER_22_151 ();
 FILLCELL_X4 FILLER_22_159 ();
 FILLCELL_X2 FILLER_22_185 ();
 FILLCELL_X16 FILLER_22_190 ();
 FILLCELL_X2 FILLER_22_206 ();
 FILLCELL_X1 FILLER_22_208 ();
 FILLCELL_X1 FILLER_22_214 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_59 ();
 FILLCELL_X1 FILLER_23_61 ();
 FILLCELL_X32 FILLER_23_66 ();
 FILLCELL_X16 FILLER_23_98 ();
 FILLCELL_X2 FILLER_23_114 ();
 FILLCELL_X1 FILLER_23_116 ();
 FILLCELL_X8 FILLER_23_134 ();
 FILLCELL_X2 FILLER_23_159 ();
 FILLCELL_X1 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_198 ();
 FILLCELL_X2 FILLER_23_228 ();
 FILLCELL_X2 FILLER_23_250 ();
 FILLCELL_X1 FILLER_24_4 ();
 FILLCELL_X1 FILLER_24_12 ();
 FILLCELL_X4 FILLER_24_23 ();
 FILLCELL_X1 FILLER_24_27 ();
 FILLCELL_X2 FILLER_24_38 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X8 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_105 ();
 FILLCELL_X8 FILLER_24_116 ();
 FILLCELL_X2 FILLER_24_141 ();
 FILLCELL_X16 FILLER_24_160 ();
 FILLCELL_X8 FILLER_24_176 ();
 FILLCELL_X4 FILLER_24_184 ();
 FILLCELL_X2 FILLER_24_188 ();
 FILLCELL_X1 FILLER_24_190 ();
 FILLCELL_X8 FILLER_24_195 ();
 FILLCELL_X2 FILLER_24_203 ();
 FILLCELL_X2 FILLER_24_217 ();
 FILLCELL_X1 FILLER_24_229 ();
 FILLCELL_X1 FILLER_24_241 ();
 FILLCELL_X1 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_26 ();
 FILLCELL_X1 FILLER_25_28 ();
 FILLCELL_X4 FILLER_25_43 ();
 FILLCELL_X1 FILLER_25_47 ();
 FILLCELL_X2 FILLER_25_52 ();
 FILLCELL_X2 FILLER_25_71 ();
 FILLCELL_X1 FILLER_25_73 ();
 FILLCELL_X2 FILLER_25_81 ();
 FILLCELL_X32 FILLER_25_91 ();
 FILLCELL_X8 FILLER_25_123 ();
 FILLCELL_X4 FILLER_25_135 ();
 FILLCELL_X2 FILLER_25_139 ();
 FILLCELL_X2 FILLER_25_144 ();
 FILLCELL_X4 FILLER_25_151 ();
 FILLCELL_X1 FILLER_25_155 ();
 FILLCELL_X32 FILLER_25_163 ();
 FILLCELL_X4 FILLER_25_219 ();
 FILLCELL_X1 FILLER_25_223 ();
 FILLCELL_X2 FILLER_25_250 ();
 FILLCELL_X1 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_25 ();
 FILLCELL_X4 FILLER_26_52 ();
 FILLCELL_X2 FILLER_26_56 ();
 FILLCELL_X1 FILLER_26_58 ();
 FILLCELL_X4 FILLER_26_66 ();
 FILLCELL_X2 FILLER_26_70 ();
 FILLCELL_X1 FILLER_26_72 ();
 FILLCELL_X2 FILLER_26_90 ();
 FILLCELL_X2 FILLER_26_109 ();
 FILLCELL_X32 FILLER_26_119 ();
 FILLCELL_X2 FILLER_26_151 ();
 FILLCELL_X2 FILLER_26_157 ();
 FILLCELL_X1 FILLER_26_159 ();
 FILLCELL_X4 FILLER_26_168 ();
 FILLCELL_X2 FILLER_26_172 ();
 FILLCELL_X1 FILLER_26_174 ();
 FILLCELL_X1 FILLER_26_179 ();
 FILLCELL_X8 FILLER_26_184 ();
 FILLCELL_X16 FILLER_26_196 ();
 FILLCELL_X8 FILLER_26_212 ();
 FILLCELL_X1 FILLER_26_220 ();
 FILLCELL_X1 FILLER_26_245 ();
 FILLCELL_X8 FILLER_27_26 ();
 FILLCELL_X16 FILLER_27_41 ();
 FILLCELL_X1 FILLER_27_74 ();
 FILLCELL_X1 FILLER_27_79 ();
 FILLCELL_X1 FILLER_27_87 ();
 FILLCELL_X1 FILLER_27_92 ();
 FILLCELL_X8 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_105 ();
 FILLCELL_X2 FILLER_27_109 ();
 FILLCELL_X2 FILLER_27_128 ();
 FILLCELL_X1 FILLER_27_147 ();
 FILLCELL_X2 FILLER_27_165 ();
 FILLCELL_X2 FILLER_27_201 ();
 FILLCELL_X2 FILLER_27_220 ();
 FILLCELL_X1 FILLER_27_226 ();
 FILLCELL_X2 FILLER_27_231 ();
 FILLCELL_X1 FILLER_27_237 ();
 FILLCELL_X8 FILLER_28_32 ();
 FILLCELL_X2 FILLER_28_40 ();
 FILLCELL_X1 FILLER_28_42 ();
 FILLCELL_X4 FILLER_28_54 ();
 FILLCELL_X2 FILLER_28_58 ();
 FILLCELL_X4 FILLER_28_64 ();
 FILLCELL_X2 FILLER_28_68 ();
 FILLCELL_X16 FILLER_28_94 ();
 FILLCELL_X1 FILLER_28_110 ();
 FILLCELL_X16 FILLER_28_118 ();
 FILLCELL_X1 FILLER_28_134 ();
 FILLCELL_X8 FILLER_28_139 ();
 FILLCELL_X2 FILLER_28_147 ();
 FILLCELL_X1 FILLER_28_149 ();
 FILLCELL_X8 FILLER_28_157 ();
 FILLCELL_X4 FILLER_28_165 ();
 FILLCELL_X16 FILLER_28_174 ();
 FILLCELL_X8 FILLER_28_190 ();
 FILLCELL_X2 FILLER_28_198 ();
 FILLCELL_X8 FILLER_28_204 ();
 FILLCELL_X1 FILLER_28_212 ();
 FILLCELL_X1 FILLER_28_251 ();
 FILLCELL_X1 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_5 ();
 FILLCELL_X16 FILLER_29_26 ();
 FILLCELL_X1 FILLER_29_42 ();
 FILLCELL_X16 FILLER_29_81 ();
 FILLCELL_X2 FILLER_29_97 ();
 FILLCELL_X1 FILLER_29_99 ();
 FILLCELL_X16 FILLER_29_121 ();
 FILLCELL_X4 FILLER_29_137 ();
 FILLCELL_X2 FILLER_29_141 ();
 FILLCELL_X4 FILLER_29_174 ();
 FILLCELL_X1 FILLER_29_178 ();
 FILLCELL_X4 FILLER_29_186 ();
 FILLCELL_X2 FILLER_29_190 ();
 FILLCELL_X1 FILLER_29_192 ();
 FILLCELL_X8 FILLER_29_217 ();
 FILLCELL_X1 FILLER_29_251 ();
 FILLCELL_X4 FILLER_30_19 ();
 FILLCELL_X8 FILLER_30_27 ();
 FILLCELL_X4 FILLER_30_35 ();
 FILLCELL_X2 FILLER_30_39 ();
 FILLCELL_X1 FILLER_30_41 ();
 FILLCELL_X4 FILLER_30_45 ();
 FILLCELL_X1 FILLER_30_49 ();
 FILLCELL_X1 FILLER_30_53 ();
 FILLCELL_X2 FILLER_30_60 ();
 FILLCELL_X1 FILLER_30_62 ();
 FILLCELL_X2 FILLER_30_66 ();
 FILLCELL_X1 FILLER_30_68 ();
 FILLCELL_X8 FILLER_30_90 ();
 FILLCELL_X2 FILLER_30_105 ();
 FILLCELL_X1 FILLER_30_107 ();
 FILLCELL_X32 FILLER_30_111 ();
 FILLCELL_X8 FILLER_30_143 ();
 FILLCELL_X2 FILLER_30_151 ();
 FILLCELL_X1 FILLER_30_153 ();
 FILLCELL_X8 FILLER_30_183 ();
 FILLCELL_X4 FILLER_30_191 ();
 FILLCELL_X1 FILLER_30_195 ();
 FILLCELL_X1 FILLER_30_203 ();
 FILLCELL_X8 FILLER_30_221 ();
 FILLCELL_X2 FILLER_30_229 ();
 FILLCELL_X1 FILLER_30_248 ();
 FILLCELL_X16 FILLER_31_1 ();
 FILLCELL_X4 FILLER_31_17 ();
 FILLCELL_X2 FILLER_31_64 ();
 FILLCELL_X1 FILLER_31_72 ();
 FILLCELL_X1 FILLER_31_111 ();
 FILLCELL_X8 FILLER_31_133 ();
 FILLCELL_X2 FILLER_31_141 ();
 FILLCELL_X1 FILLER_31_143 ();
 FILLCELL_X4 FILLER_31_148 ();
 FILLCELL_X16 FILLER_31_213 ();
 FILLCELL_X8 FILLER_31_229 ();
 FILLCELL_X1 FILLER_31_237 ();
 FILLCELL_X2 FILLER_31_241 ();
 FILLCELL_X1 FILLER_32_83 ();
 FILLCELL_X1 FILLER_32_91 ();
 FILLCELL_X1 FILLER_32_112 ();
 FILLCELL_X2 FILLER_32_120 ();
 FILLCELL_X1 FILLER_32_122 ();
 FILLCELL_X2 FILLER_32_196 ();
 FILLCELL_X1 FILLER_32_216 ();
 FILLCELL_X1 FILLER_32_251 ();
 FILLCELL_X1 FILLER_33_18 ();
 FILLCELL_X1 FILLER_33_53 ();
 FILLCELL_X1 FILLER_33_61 ();
 FILLCELL_X2 FILLER_33_238 ();
 FILLCELL_X8 FILLER_33_243 ();
 FILLCELL_X1 FILLER_33_251 ();
endmodule
