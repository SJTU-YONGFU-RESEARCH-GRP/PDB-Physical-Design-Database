module parameterized_uart_rx (clk,
    data_valid,
    frame_error,
    parity_error,
    rst_n,
    rx,
    data_out);
 input clk;
 output data_valid;
 output frame_error;
 output parity_error;
 input rst_n;
 input rx;
 output [7:0] data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire \bit_index[0] ;
 wire \bit_index[1] ;
 wire \bit_index[2] ;
 wire \clk_counter[0] ;
 wire \clk_counter[10] ;
 wire \clk_counter[11] ;
 wire \clk_counter[12] ;
 wire \clk_counter[13] ;
 wire \clk_counter[14] ;
 wire \clk_counter[15] ;
 wire \clk_counter[16] ;
 wire \clk_counter[17] ;
 wire \clk_counter[18] ;
 wire \clk_counter[19] ;
 wire \clk_counter[1] ;
 wire \clk_counter[20] ;
 wire \clk_counter[21] ;
 wire \clk_counter[22] ;
 wire \clk_counter[23] ;
 wire \clk_counter[24] ;
 wire \clk_counter[25] ;
 wire \clk_counter[26] ;
 wire \clk_counter[27] ;
 wire \clk_counter[28] ;
 wire \clk_counter[29] ;
 wire \clk_counter[2] ;
 wire \clk_counter[30] ;
 wire \clk_counter[31] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \clk_counter[6] ;
 wire \clk_counter[7] ;
 wire \clk_counter[8] ;
 wire \clk_counter[9] ;
 wire \rx_data[0] ;
 wire \rx_data[1] ;
 wire \rx_data[2] ;
 wire \rx_data[3] ;
 wire \rx_data[4] ;
 wire \rx_data[5] ;
 wire \rx_data[6] ;
 wire \rx_data[7] ;
 wire rx_meta;
 wire rx_sync;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net15;

 gf180mcu_fd_sc_mcu9t5v0__or2_2 _343_ (.A1(\clk_counter[17] ),
    .A2(\clk_counter[16] ),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _344_ (.A1(\clk_counter[13] ),
    .A2(\clk_counter[12] ),
    .A3(\clk_counter[15] ),
    .A4(\clk_counter[14] ),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _345_ (.A1(\clk_counter[8] ),
    .A2(\clk_counter[11] ),
    .A3(\clk_counter[10] ),
    .A4(\clk_counter[19] ),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _346_ (.A1(\clk_counter[7] ),
    .A2(\clk_counter[6] ),
    .A3(\clk_counter[9] ),
    .A4(\clk_counter[30] ),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _347_ (.A1(_057_),
    .A2(_058_),
    .A3(_059_),
    .A4(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _348_ (.A1(\clk_counter[24] ),
    .A2(\clk_counter[29] ),
    .A3(\clk_counter[28] ),
    .A4(\clk_counter[31] ),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _349_ (.A1(\clk_counter[18] ),
    .A2(\clk_counter[25] ),
    .A3(\clk_counter[27] ),
    .A4(\clk_counter[26] ),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _350_ (.A1(\clk_counter[21] ),
    .A2(\clk_counter[20] ),
    .A3(\clk_counter[23] ),
    .A4(\clk_counter[22] ),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _351_ (.A1(_062_),
    .A2(_063_),
    .A3(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _352_ (.I(\clk_counter[3] ),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _353_ (.I(\clk_counter[2] ),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _354_ (.A1(\clk_counter[5] ),
    .A2(\clk_counter[4] ),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _355_ (.A1(_066_),
    .A2(_067_),
    .A3(_327_),
    .A4(_068_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _356_ (.A1(_061_),
    .A2(_065_),
    .A3(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _357_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _358_ (.A1(\state[2] ),
    .A2(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _359_ (.A1(_070_),
    .A2(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _360_ (.I(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _361_ (.I(_074_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _362_ (.I(\clk_counter[0] ),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _363_ (.I(\bit_index[0] ),
    .ZN(_333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _364_ (.I(\clk_counter[1] ),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _365_ (.I(\bit_index[1] ),
    .ZN(_334_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _366_ (.I(\state[1] ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _367_ (.A1(_075_),
    .A2(\state[0] ),
    .A3(\state[2] ),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _368_ (.A1(_341_),
    .A2(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _369_ (.A1(\bit_index[0] ),
    .A2(_077_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _370_ (.A1(_057_),
    .A2(_058_),
    .A3(_059_),
    .A4(_060_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _371_ (.A1(_062_),
    .A2(_063_),
    .A3(_064_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _372_ (.A1(_079_),
    .A2(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _373_ (.I(\state[0] ),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _374_ (.I(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _375_ (.A1(_066_),
    .A2(_067_),
    .A3(_327_),
    .A4(_068_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _376_ (.I(\state[1] ),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _377_ (.I(rx_sync),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _378_ (.A1(_085_),
    .A2(_086_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _379_ (.A1(\clk_counter[4] ),
    .A2(_329_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _380_ (.A1(_066_),
    .A2(\clk_counter[2] ),
    .A3(\clk_counter[5] ),
    .A4(_088_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _381_ (.A1(_083_),
    .A2(_084_),
    .B1(_087_),
    .B2(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _382_ (.I(\state[2] ),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _383_ (.I(_091_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _384_ (.A1(_092_),
    .A2(_071_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _385_ (.A1(\state[2] ),
    .A2(_081_),
    .A3(_090_),
    .B(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _386_ (.I0(\bit_index[0] ),
    .I1(_078_),
    .S(_094_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _387_ (.I(_336_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _388_ (.A1(_095_),
    .A2(_077_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _389_ (.I0(\bit_index[1] ),
    .I1(_096_),
    .S(_094_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _390_ (.A1(_085_),
    .A2(_083_),
    .A3(_092_),
    .A4(_342_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _391_ (.I0(\bit_index[2] ),
    .I1(_097_),
    .S(_094_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _392_ (.A1(_085_),
    .A2(\state[2] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _393_ (.A1(_066_),
    .A2(\clk_counter[2] ),
    .A3(\clk_counter[5] ),
    .A4(_088_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _394_ (.A1(_075_),
    .A2(_082_),
    .A3(_091_),
    .A4(rx_sync),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _395_ (.A1(_061_),
    .A2(_065_),
    .A3(_099_),
    .A4(_100_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _396_ (.A1(_098_),
    .A2(_101_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _397_ (.I(\clk_counter[5] ),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _398_ (.A1(_103_),
    .A2(_325_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _399_ (.I(\clk_counter[4] ),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _400_ (.A1(\clk_counter[3] ),
    .A2(\clk_counter[2] ),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _401_ (.A1(_105_),
    .A2(\state[2] ),
    .A3(_106_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _402_ (.A1(_075_),
    .A2(_082_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _403_ (.A1(_092_),
    .A2(_089_),
    .B1(_104_),
    .B2(_107_),
    .C(_108_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _404_ (.A1(_085_),
    .A2(_092_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _405_ (.A1(_072_),
    .A2(_110_),
    .B(_084_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _406_ (.A1(_085_),
    .A2(\state[2] ),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _407_ (.A1(_079_),
    .A2(_080_),
    .B1(_071_),
    .B2(_092_),
    .C(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _408_ (.A1(_109_),
    .A2(_111_),
    .A3(_113_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _409_ (.I0(_102_),
    .I1(_114_),
    .S(_323_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _410_ (.I(\clk_counter[10] ),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _411_ (.A1(_098_),
    .A2(_101_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _412_ (.A1(_109_),
    .A2(_111_),
    .A3(_113_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _413_ (.A1(\clk_counter[3] ),
    .A2(\clk_counter[2] ),
    .A3(_331_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _414_ (.A1(\clk_counter[7] ),
    .A2(\clk_counter[6] ),
    .A3(_068_),
    .A4(_118_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _415_ (.A1(\clk_counter[9] ),
    .A2(\clk_counter[8] ),
    .A3(_119_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _416_ (.A1(\clk_counter[10] ),
    .A2(_120_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _417_ (.A1(_115_),
    .A2(_116_),
    .B1(_117_),
    .B2(_121_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _418_ (.I(\clk_counter[11] ),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _419_ (.I(_116_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _420_ (.I(_109_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _421_ (.I(_111_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _422_ (.I(_113_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _423_ (.A1(\clk_counter[3] ),
    .A2(\clk_counter[2] ),
    .A3(\clk_counter[0] ),
    .A4(\clk_counter[1] ),
    .Z(_127_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _424_ (.A1(\clk_counter[5] ),
    .A2(\clk_counter[4] ),
    .A3(\clk_counter[6] ),
    .Z(_128_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _425_ (.A1(\clk_counter[9] ),
    .A2(\clk_counter[8] ),
    .A3(\clk_counter[10] ),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _426_ (.A1(\clk_counter[7] ),
    .A2(_127_),
    .A3(_128_),
    .A4(_129_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _427_ (.A1(\clk_counter[11] ),
    .A2(_130_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _428_ (.A1(\clk_counter[11] ),
    .A2(_130_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _429_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_131_),
    .B2(_132_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _430_ (.A1(_122_),
    .A2(_123_),
    .B(_133_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _431_ (.I(\clk_counter[12] ),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _432_ (.A1(\clk_counter[9] ),
    .A2(\clk_counter[8] ),
    .A3(\clk_counter[11] ),
    .A4(\clk_counter[10] ),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _433_ (.A1(_134_),
    .A2(_119_),
    .A3(_135_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _434_ (.A1(_119_),
    .A2(_135_),
    .B(_134_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _435_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_136_),
    .B2(_137_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _436_ (.A1(_134_),
    .A2(_123_),
    .B(_138_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _437_ (.I(\clk_counter[13] ),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _438_ (.A1(\clk_counter[5] ),
    .A2(\clk_counter[4] ),
    .A3(\clk_counter[7] ),
    .A4(\clk_counter[6] ),
    .Z(_140_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _439_ (.A1(\clk_counter[12] ),
    .A2(_127_),
    .A3(_135_),
    .A4(_140_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _440_ (.A1(\clk_counter[13] ),
    .A2(_141_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _441_ (.A1(\clk_counter[13] ),
    .A2(_141_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _442_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_142_),
    .B2(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _443_ (.A1(_139_),
    .A2(_123_),
    .B(_144_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _444_ (.I(\clk_counter[14] ),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _445_ (.A1(\clk_counter[13] ),
    .A2(\clk_counter[12] ),
    .A3(_119_),
    .A4(_135_),
    .Z(_146_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _446_ (.A1(\clk_counter[14] ),
    .A2(_146_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _447_ (.A1(_145_),
    .A2(_116_),
    .B1(_117_),
    .B2(_147_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _448_ (.I(\clk_counter[15] ),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _449_ (.A1(\clk_counter[13] ),
    .A2(\clk_counter[12] ),
    .A3(\clk_counter[14] ),
    .Z(_149_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _450_ (.A1(_127_),
    .A2(_135_),
    .A3(_140_),
    .A4(_149_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _451_ (.I(_150_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _452_ (.A1(_148_),
    .A2(_151_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _453_ (.A1(_148_),
    .A2(_151_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _454_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_152_),
    .B2(_153_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _455_ (.A1(_148_),
    .A2(_123_),
    .B(_154_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _456_ (.I(\clk_counter[16] ),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _457_ (.A1(_118_),
    .A2(_135_),
    .A3(_140_),
    .A4(_149_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _458_ (.I(_156_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _459_ (.A1(\clk_counter[15] ),
    .A2(_155_),
    .A3(_157_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _460_ (.A1(\clk_counter[15] ),
    .A2(_157_),
    .B(_155_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _461_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_158_),
    .B2(_159_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _462_ (.A1(_155_),
    .A2(_123_),
    .B(_160_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _463_ (.I(\clk_counter[17] ),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _464_ (.A1(\clk_counter[15] ),
    .A2(\clk_counter[16] ),
    .Z(_162_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _465_ (.A1(_161_),
    .A2(_150_),
    .A3(_162_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _466_ (.A1(_151_),
    .A2(_162_),
    .B(_161_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _467_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_163_),
    .B2(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _468_ (.A1(_161_),
    .A2(_123_),
    .B(_165_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _469_ (.I(\clk_counter[18] ),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _470_ (.A1(_118_),
    .A2(_135_),
    .A3(_140_),
    .A4(_149_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _471_ (.A1(\clk_counter[15] ),
    .A2(\clk_counter[17] ),
    .A3(\clk_counter[16] ),
    .Z(_168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _472_ (.A1(_167_),
    .A2(_168_),
    .B(_166_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _473_ (.A1(_166_),
    .A2(_167_),
    .A3(_168_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _474_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B1(_169_),
    .B2(_170_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _475_ (.A1(_166_),
    .A2(_123_),
    .B(_171_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _476_ (.I(\clk_counter[19] ),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _477_ (.I(_109_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _478_ (.I(_111_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _479_ (.I(_113_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _480_ (.A1(\clk_counter[18] ),
    .A2(_168_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _481_ (.A1(_151_),
    .A2(_176_),
    .B(_172_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _482_ (.A1(_172_),
    .A2(_150_),
    .A3(_176_),
    .Z(_178_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _483_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_177_),
    .B2(_178_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _484_ (.A1(_172_),
    .A2(_123_),
    .B(_179_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _485_ (.I(_326_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _486_ (.A1(_324_),
    .A2(_116_),
    .B1(_117_),
    .B2(_180_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _487_ (.I(\clk_counter[20] ),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _488_ (.A1(\clk_counter[19] ),
    .A2(\clk_counter[18] ),
    .A3(_156_),
    .A4(_168_),
    .Z(_182_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _489_ (.A1(\clk_counter[20] ),
    .A2(_182_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _490_ (.A1(_181_),
    .A2(_116_),
    .B1(_117_),
    .B2(_183_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _491_ (.I(\clk_counter[21] ),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _492_ (.A1(\clk_counter[19] ),
    .A2(\clk_counter[18] ),
    .A3(\clk_counter[20] ),
    .Z(_185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _493_ (.A1(_168_),
    .A2(_185_),
    .Z(_186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _494_ (.A1(_151_),
    .A2(_186_),
    .B(_184_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _495_ (.A1(_184_),
    .A2(_150_),
    .A3(_186_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _496_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_187_),
    .B2(_188_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _497_ (.A1(_184_),
    .A2(_123_),
    .B(_189_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _498_ (.I(\clk_counter[22] ),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _499_ (.A1(\clk_counter[21] ),
    .A2(_168_),
    .A3(_185_),
    .Z(_191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _500_ (.A1(_157_),
    .A2(_191_),
    .B(_190_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _501_ (.A1(_190_),
    .A2(_157_),
    .A3(_191_),
    .Z(_193_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _502_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_192_),
    .B2(_193_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _503_ (.A1(_190_),
    .A2(_123_),
    .B(_194_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _504_ (.I(\clk_counter[23] ),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _505_ (.I(_116_),
    .Z(_196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _506_ (.A1(\clk_counter[21] ),
    .A2(\clk_counter[22] ),
    .Z(_197_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _507_ (.A1(_168_),
    .A2(_185_),
    .A3(_197_),
    .Z(_198_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _508_ (.I(_198_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _509_ (.A1(_195_),
    .A2(_150_),
    .A3(_199_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _510_ (.A1(_151_),
    .A2(_199_),
    .B(_195_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _511_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_200_),
    .B2(_201_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _512_ (.A1(_195_),
    .A2(_196_),
    .B(_202_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _513_ (.I(\clk_counter[24] ),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _514_ (.I(_109_),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _515_ (.I(_111_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _516_ (.I(_113_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _517_ (.A1(\clk_counter[23] ),
    .A2(_157_),
    .A3(_199_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _518_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_207_),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _519_ (.A1(\clk_counter[23] ),
    .A2(_203_),
    .A3(_156_),
    .A4(_198_),
    .Z(_209_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _520_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_209_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _521_ (.A1(_061_),
    .A2(_065_),
    .A3(_099_),
    .A4(_100_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _522_ (.A1(_112_),
    .A2(_211_),
    .B(\clk_counter[24] ),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _523_ (.A1(_203_),
    .A2(_208_),
    .B(_210_),
    .C(_212_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _524_ (.I(\clk_counter[25] ),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _525_ (.A1(\clk_counter[23] ),
    .A2(\clk_counter[24] ),
    .Z(_214_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _526_ (.A1(_168_),
    .A2(_185_),
    .A3(_197_),
    .A4(_214_),
    .Z(_215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _527_ (.A1(_151_),
    .A2(_215_),
    .B(_213_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _528_ (.A1(_213_),
    .A2(_150_),
    .A3(_215_),
    .Z(_217_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _529_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_216_),
    .B2(_217_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _530_ (.A1(_213_),
    .A2(_196_),
    .B(_218_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _531_ (.I(\clk_counter[26] ),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _532_ (.A1(\clk_counter[23] ),
    .A2(\clk_counter[22] ),
    .A3(\clk_counter[25] ),
    .A4(\clk_counter[24] ),
    .Z(_220_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _533_ (.A1(\clk_counter[21] ),
    .A2(_168_),
    .A3(_185_),
    .A4(_220_),
    .Z(_221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _534_ (.A1(_157_),
    .A2(_221_),
    .B(_219_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _535_ (.A1(_219_),
    .A2(_157_),
    .A3(_221_),
    .Z(_223_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _536_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_222_),
    .B2(_223_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _537_ (.A1(_219_),
    .A2(_196_),
    .B(_224_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _538_ (.I(\clk_counter[27] ),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _539_ (.A1(\clk_counter[23] ),
    .A2(\clk_counter[25] ),
    .A3(\clk_counter[24] ),
    .A4(\clk_counter[26] ),
    .Z(_226_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _540_ (.A1(_150_),
    .A2(_199_),
    .A3(_226_),
    .Z(_227_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _541_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _542_ (.A1(\clk_counter[27] ),
    .A2(_098_),
    .A3(_101_),
    .Z(_229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _543_ (.A1(_151_),
    .A2(_199_),
    .A3(_226_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _544_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_230_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _545_ (.A1(_225_),
    .A2(_228_),
    .B1(_229_),
    .B2(_231_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _546_ (.I(\clk_counter[28] ),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _547_ (.A1(\clk_counter[27] ),
    .A2(_156_),
    .A3(_198_),
    .A4(_226_),
    .Z(_233_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _548_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_233_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _549_ (.A1(\clk_counter[28] ),
    .A2(_098_),
    .A3(_101_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _550_ (.A1(\clk_counter[27] ),
    .A2(_157_),
    .A3(_199_),
    .A4(_226_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _551_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_236_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _552_ (.A1(_232_),
    .A2(_234_),
    .B1(_235_),
    .B2(_237_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _553_ (.I(\clk_counter[29] ),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _554_ (.A1(\clk_counter[27] ),
    .A2(\clk_counter[28] ),
    .A3(_226_),
    .Z(_239_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _555_ (.A1(_150_),
    .A2(_199_),
    .A3(_239_),
    .Z(_240_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _556_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_240_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _557_ (.A1(\clk_counter[29] ),
    .A2(_098_),
    .A3(_101_),
    .Z(_242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _558_ (.A1(_151_),
    .A2(_199_),
    .A3(_239_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _559_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_243_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _560_ (.A1(_238_),
    .A2(_241_),
    .B1(_242_),
    .B2(_244_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _561_ (.A1(_067_),
    .A2(_331_),
    .Z(_245_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _562_ (.A1(_067_),
    .A2(_331_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _563_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_245_),
    .B2(_246_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _564_ (.A1(_067_),
    .A2(_196_),
    .B(_247_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _565_ (.I(\clk_counter[30] ),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _566_ (.A1(\clk_counter[27] ),
    .A2(\clk_counter[29] ),
    .A3(\clk_counter[28] ),
    .A4(_226_),
    .Z(_249_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _567_ (.A1(_157_),
    .A2(_198_),
    .A3(_249_),
    .Z(_250_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _568_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _569_ (.A1(\clk_counter[30] ),
    .A2(_098_),
    .A3(_101_),
    .Z(_252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _570_ (.A1(_157_),
    .A2(_199_),
    .A3(_249_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _571_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B(_253_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _572_ (.A1(_248_),
    .A2(_251_),
    .B1(_252_),
    .B2(_254_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _573_ (.I(\clk_counter[31] ),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _574_ (.A1(\clk_counter[30] ),
    .A2(_150_),
    .A3(_198_),
    .A4(_249_),
    .Z(_256_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _575_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .B(_256_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _576_ (.A1(\clk_counter[31] ),
    .A2(_098_),
    .A3(_101_),
    .Z(_258_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _577_ (.A1(\clk_counter[30] ),
    .A2(_151_),
    .A3(_199_),
    .A4(_249_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _578_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B(_259_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _579_ (.A1(_255_),
    .A2(_257_),
    .B1(_258_),
    .B2(_260_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _580_ (.A1(_067_),
    .A2(_323_),
    .A3(_324_),
    .Z(_261_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _581_ (.A1(\clk_counter[3] ),
    .A2(_261_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _582_ (.A1(\clk_counter[3] ),
    .A2(_261_),
    .Z(_263_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _583_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_262_),
    .B2(_263_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _584_ (.A1(_066_),
    .A2(_196_),
    .B(_264_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _585_ (.A1(_105_),
    .A2(_118_),
    .Z(_265_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _586_ (.A1(_105_),
    .A2(_118_),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _587_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_265_),
    .B2(_266_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _588_ (.A1(_105_),
    .A2(_196_),
    .B(_267_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _589_ (.A1(\clk_counter[4] ),
    .A2(_127_),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _590_ (.A1(\clk_counter[5] ),
    .A2(_268_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _591_ (.A1(\clk_counter[5] ),
    .A2(_268_),
    .Z(_270_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _592_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .B1(_269_),
    .B2(_270_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _593_ (.A1(_103_),
    .A2(_196_),
    .B(_271_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _594_ (.I(\clk_counter[6] ),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _595_ (.A1(_068_),
    .A2(_118_),
    .ZN(_273_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _596_ (.A1(\clk_counter[6] ),
    .A2(_273_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _597_ (.A1(\clk_counter[6] ),
    .A2(_273_),
    .Z(_275_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _598_ (.A1(_109_),
    .A2(_111_),
    .A3(_113_),
    .B1(_274_),
    .B2(_275_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _599_ (.A1(_272_),
    .A2(_196_),
    .B(_276_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _600_ (.I(\clk_counter[7] ),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _601_ (.A1(_127_),
    .A2(_128_),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _602_ (.A1(\clk_counter[7] ),
    .A2(_278_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _603_ (.A1(\clk_counter[7] ),
    .A2(_278_),
    .Z(_280_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _604_ (.A1(_109_),
    .A2(_111_),
    .A3(_113_),
    .B1(_279_),
    .B2(_280_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _605_ (.A1(_277_),
    .A2(_196_),
    .B(_281_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _606_ (.I(\clk_counter[8] ),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _607_ (.A1(_282_),
    .A2(_119_),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _608_ (.A1(_282_),
    .A2(_119_),
    .Z(_284_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _609_ (.A1(_109_),
    .A2(_111_),
    .A3(_113_),
    .B1(_283_),
    .B2(_284_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _610_ (.A1(_282_),
    .A2(_196_),
    .B(_285_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _611_ (.I(\clk_counter[9] ),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _612_ (.A1(_277_),
    .A2(_282_),
    .A3(_278_),
    .B(\clk_counter[9] ),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _613_ (.A1(_277_),
    .A2(\clk_counter[9] ),
    .A3(_282_),
    .A4(_278_),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _614_ (.A1(_124_),
    .A2(_125_),
    .A3(_126_),
    .B(_288_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _615_ (.A1(_286_),
    .A2(_116_),
    .B1(_117_),
    .B2(_287_),
    .C(_289_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _616_ (.I0(\rx_data[0] ),
    .I1(net4),
    .S(_074_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _617_ (.I0(\rx_data[1] ),
    .I1(net5),
    .S(_074_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _618_ (.I0(\rx_data[2] ),
    .I1(net6),
    .S(_074_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _619_ (.I0(\rx_data[3] ),
    .I1(net7),
    .S(_074_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _620_ (.I0(\rx_data[4] ),
    .I1(net8),
    .S(_074_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _621_ (.I0(\rx_data[5] ),
    .I1(net9),
    .S(_074_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _622_ (.I0(\rx_data[6] ),
    .I1(net10),
    .S(_074_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _623_ (.I0(\rx_data[7] ),
    .I1(net11),
    .S(_074_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _624_ (.A1(_085_),
    .A2(_082_),
    .A3(_086_),
    .A4(_070_),
    .Z(_290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _625_ (.I(net13),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _626_ (.A1(_092_),
    .A2(_071_),
    .B1(_290_),
    .B2(_291_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _627_ (.A1(_082_),
    .A2(_092_),
    .A3(_086_),
    .Z(_292_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _628_ (.A1(_079_),
    .A2(_080_),
    .A3(_084_),
    .A4(_292_),
    .Z(_293_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _629_ (.A1(net14),
    .A2(_293_),
    .B(_085_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _630_ (.A1(_082_),
    .A2(\state[2] ),
    .B(net14),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _631_ (.A1(_294_),
    .A2(_295_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _632_ (.A1(_061_),
    .A2(_065_),
    .A3(_069_),
    .A4(_076_),
    .Z(_296_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _633_ (.A1(\bit_index[2] ),
    .A2(_335_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _634_ (.A1(\bit_index[0] ),
    .A2(\bit_index[1] ),
    .A3(\bit_index[2] ),
    .A4(_336_),
    .Z(_298_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _635_ (.A1(_296_),
    .A2(_297_),
    .A3(_298_),
    .Z(_299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _636_ (.I0(_086_),
    .I1(\rx_data[0] ),
    .S(_299_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _637_ (.A1(\bit_index[2] ),
    .A2(_335_),
    .Z(_300_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _638_ (.A1(_296_),
    .A2(_300_),
    .Z(_301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _639_ (.A1(_086_),
    .A2(\bit_index[0] ),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _640_ (.A1(_095_),
    .A2(_302_),
    .Z(_303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _641_ (.A1(_337_),
    .A2(_297_),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _642_ (.A1(_296_),
    .A2(_304_),
    .B(\rx_data[1] ),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _643_ (.A1(_301_),
    .A2(_303_),
    .B(_305_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _644_ (.A1(\bit_index[1] ),
    .A2(\bit_index[2] ),
    .B(_333_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _645_ (.A1(_095_),
    .A2(_296_),
    .A3(_300_),
    .A4(_306_),
    .Z(_307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _646_ (.I0(_086_),
    .I1(\rx_data[2] ),
    .S(_307_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _647_ (.A1(_339_),
    .A2(_297_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _648_ (.A1(_296_),
    .A2(_308_),
    .B(\rx_data[3] ),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _649_ (.A1(_336_),
    .A2(_301_),
    .A3(_302_),
    .B(_309_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _650_ (.A1(_336_),
    .A2(_296_),
    .A3(_300_),
    .A4(_306_),
    .Z(_310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _651_ (.I0(_086_),
    .I1(\rx_data[4] ),
    .S(_310_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _652_ (.A1(_296_),
    .A2(_297_),
    .Z(_311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _653_ (.A1(_337_),
    .A2(_300_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _654_ (.A1(_296_),
    .A2(_312_),
    .B(\rx_data[5] ),
    .ZN(_313_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _655_ (.A1(_311_),
    .A2(_303_),
    .B(_313_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _656_ (.A1(_095_),
    .A2(_296_),
    .A3(_297_),
    .A4(_306_),
    .Z(_314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _657_ (.I0(_086_),
    .I1(\rx_data[6] ),
    .S(_314_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _658_ (.A1(_339_),
    .A2(_300_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _659_ (.A1(_296_),
    .A2(_315_),
    .B(\rx_data[7] ),
    .ZN(_316_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _660_ (.A1(_336_),
    .A2(_311_),
    .A3(_302_),
    .B(_316_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _661_ (.A1(_092_),
    .A2(_086_),
    .B(_085_),
    .C(_082_),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _662_ (.I0(_082_),
    .I1(_317_),
    .S(_117_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _663_ (.I0(_077_),
    .I1(\state[2] ),
    .S(_070_),
    .Z(_318_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _664_ (.A1(\state[2] ),
    .A2(_086_),
    .A3(_108_),
    .Z(_319_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _665_ (.A1(_075_),
    .A2(_318_),
    .B1(_319_),
    .B2(_114_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _666_ (.A1(_082_),
    .A2(_079_),
    .A3(_080_),
    .Z(_320_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _667_ (.A1(_105_),
    .A2(_106_),
    .A3(_104_),
    .A4(_320_),
    .Z(_321_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _668_ (.A1(_082_),
    .A2(_341_),
    .B(_092_),
    .C(_085_),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _669_ (.A1(_085_),
    .A2(_092_),
    .A3(_321_),
    .B1(_322_),
    .B2(_070_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _670_ (.A(_323_),
    .B(_324_),
    .CO(_325_),
    .S(_326_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _671_ (.A(_323_),
    .B(\clk_counter[1] ),
    .CO(_327_),
    .S(_328_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _672_ (.A(\clk_counter[0] ),
    .B(_324_),
    .CO(_329_),
    .S(_330_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _673_ (.A(\clk_counter[0] ),
    .B(\clk_counter[1] ),
    .CO(_331_),
    .S(_332_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _674_ (.A(_333_),
    .B(_334_),
    .CO(_335_),
    .S(_336_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _675_ (.A(\bit_index[0] ),
    .B(_334_),
    .CO(_337_),
    .S(_338_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _676_ (.A(\bit_index[0] ),
    .B(\bit_index[1] ),
    .CO(_339_),
    .S(_340_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _677_ (.A(\bit_index[2] ),
    .B(_339_),
    .CO(_341_),
    .S(_342_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_index[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\bit_index[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_index[1]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\bit_index[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_index[2]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\bit_index[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[0]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\clk_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[10]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[11]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[12]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[13]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[14]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[15]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[16]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[17]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[18]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[19]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[1]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\clk_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[20]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[21]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\clk_counter[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[22]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[23]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[24]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\clk_counter[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[25]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[26]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[27]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[28]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[29]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[2]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[30]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\clk_counter[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[31]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\clk_counter[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[3]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[4]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[5]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[6]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[7]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\clk_counter[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[8]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[9]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\clk_counter[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[0]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[1]$_DFFE_PN0P_  (.D(_037_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[2]$_DFFE_PN0P_  (.D(_038_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[3]$_DFFE_PN0P_  (.D(_039_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[4]$_DFFE_PN0P_  (.D(_040_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[5]$_DFFE_PN0P_  (.D(_041_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[6]$_DFFE_PN0P_  (.D(_042_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_out[7]$_DFFE_PN0P_  (.D(_043_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_valid$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \frame_error$_DFFE_PN0P_  (.D(_044_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \parity_error$_DFFE_PN0P_  (.D(_045_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_046_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\rx_data[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_047_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\rx_data[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_048_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\rx_data[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_049_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\rx_data[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_050_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\rx_data[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_051_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\rx_data[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_052_),
    .RN(net1),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\rx_data[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_053_),
    .RN(net1),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\rx_data[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \rx_meta$_DFF_PN1_  (.D(net3),
    .SETN(net2),
    .CLK(clknet_3_5__leaf_clk),
    .Q(rx_meta));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \rx_sync$_DFF_PN1_  (.D(rx_meta),
    .SETN(net2),
    .CLK(clknet_3_5__leaf_clk),
    .Q(rx_sync));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[0]$_DFFE_PN0P_  (.D(_054_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFFE_PN0P_  (.D(_055_),
    .RN(net1),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[2]$_DFFE_PN0P_  (.D(_056_),
    .RN(net1),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_83 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_84 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_90 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_124 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input1 (.I(net15),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(rx),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net4),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net5),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net7),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net8),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net9),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net10),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net11),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net12),
    .Z(data_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(frame_error));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(parity_error));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_4__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_5__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_6__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_3_7__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload0 (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload1 (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload2 (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload3 (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload4 (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload5 (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload6 (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_378 ();
endmodule
