module elastic_buffer (rd_almost_empty,
    rd_clk,
    rd_empty,
    rd_en,
    rd_rst_n,
    wr_almost_full,
    wr_clk,
    wr_en,
    wr_full,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output rd_almost_empty;
 input rd_clk;
 output rd_empty;
 input rd_en;
 input rd_rst_n;
 output wr_almost_full;
 input wr_clk;
 input wr_en;
 output wr_full;
 input wr_rst_n;
 output [3:0] rd_count;
 output [7:0] rd_data;
 output [3:0] wr_count;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin_sync[3] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin_sync[3] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;

 XOR2_X2 _348_ (.A(_332_),
    .B(_322_),
    .Z(net10));
 XNOR2_X2 _349_ (.A(\wr_ptr_bin_sync[3] ),
    .B(\rd_ptr_bin[3] ),
    .ZN(_091_));
 INV_X1 _350_ (.A(_333_),
    .ZN(_092_));
 INV_X1 _351_ (.A(_334_),
    .ZN(_093_));
 OAI21_X1 _352_ (.A(_092_),
    .B1(_093_),
    .B2(_344_),
    .ZN(_094_));
 AOI21_X2 _353_ (.A(_331_),
    .B1(_094_),
    .B2(_332_),
    .ZN(_095_));
 XNOR2_X2 _354_ (.A(_091_),
    .B(_095_),
    .ZN(net11));
 INV_X1 _355_ (.A(_345_),
    .ZN(net8));
 XNOR2_X2 _356_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(\rd_ptr_bin_sync[3] ),
    .ZN(_338_));
 XNOR2_X2 _357_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(_338_),
    .ZN(_326_));
 INV_X1 _358_ (.A(_326_),
    .ZN(_335_));
 INV_X2 _359_ (.A(_347_),
    .ZN(net22));
 XNOR2_X2 _360_ (.A(_340_),
    .B(_327_),
    .ZN(net24));
 XOR2_X2 _361_ (.A(\rd_ptr_bin_sync[3] ),
    .B(\wr_ptr_bin[3] ),
    .Z(_096_));
 INV_X1 _362_ (.A(_336_),
    .ZN(_097_));
 INV_X1 _363_ (.A(_337_),
    .ZN(_098_));
 OAI21_X1 _364_ (.A(_097_),
    .B1(_325_),
    .B2(_098_),
    .ZN(_099_));
 AOI21_X2 _365_ (.A(_339_),
    .B1(_099_),
    .B2(_340_),
    .ZN(_100_));
 XNOR2_X2 _366_ (.A(_096_),
    .B(_100_),
    .ZN(_101_));
 INV_X1 _367_ (.A(_101_),
    .ZN(net25));
 XNOR2_X2 _368_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(\rd_ptr_gray[0] ),
    .ZN(_102_));
 XNOR2_X2 _369_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(\rd_ptr_gray[2] ),
    .ZN(_103_));
 XNOR2_X2 _370_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(\rd_ptr_gray[1] ),
    .ZN(_104_));
 NAND4_X4 _371_ (.A1(_091_),
    .A2(_102_),
    .A3(_103_),
    .A4(_104_),
    .ZN(_105_));
 INV_X1 _372_ (.A(_105_),
    .ZN(net20));
 XNOR2_X2 _373_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(\wr_ptr_gray[0] ),
    .ZN(_106_));
 XNOR2_X2 _374_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(\wr_ptr_gray[2] ),
    .ZN(_107_));
 XNOR2_X2 _375_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(\wr_ptr_gray[1] ),
    .ZN(_108_));
 NAND4_X4 _376_ (.A1(_096_),
    .A2(_106_),
    .A3(_107_),
    .A4(_108_),
    .ZN(_109_));
 INV_X1 _377_ (.A(_109_),
    .ZN(net26));
 XOR2_X2 _378_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(\wr_ptr_bin_sync[3] ),
    .Z(_330_));
 XOR2_X2 _379_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(_330_),
    .Z(_320_));
 XOR2_X2 _380_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(_326_),
    .Z(_346_));
 INV_X1 _381_ (.A(_344_),
    .ZN(_319_));
 XNOR2_X1 _382_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(_320_),
    .ZN(_343_));
 BUF_X2 _383_ (.A(wr_data[0]),
    .Z(_110_));
 CLKBUF_X3 _384_ (.A(\wr_ptr_bin[2] ),
    .Z(_111_));
 BUF_X4 _385_ (.A(\wr_ptr_bin[1] ),
    .Z(_112_));
 CLKBUF_X3 _386_ (.A(\wr_ptr_bin[0] ),
    .Z(_113_));
 NAND2_X2 _387_ (.A1(net5),
    .A2(_109_),
    .ZN(_114_));
 BUF_X8 _388_ (.A(_114_),
    .Z(_115_));
 NOR4_X4 _389_ (.A1(_111_),
    .A2(_112_),
    .A3(_113_),
    .A4(_115_),
    .ZN(_116_));
 MUX2_X1 _390_ (.A(\mem[0][0] ),
    .B(_110_),
    .S(_116_),
    .Z(_005_));
 CLKBUF_X2 _391_ (.A(wr_data[1]),
    .Z(_117_));
 MUX2_X1 _392_ (.A(\mem[0][1] ),
    .B(_117_),
    .S(_116_),
    .Z(_006_));
 CLKBUF_X2 _393_ (.A(wr_data[2]),
    .Z(_118_));
 MUX2_X1 _394_ (.A(\mem[0][2] ),
    .B(_118_),
    .S(_116_),
    .Z(_007_));
 CLKBUF_X2 _395_ (.A(wr_data[3]),
    .Z(_119_));
 MUX2_X1 _396_ (.A(\mem[0][3] ),
    .B(_119_),
    .S(_116_),
    .Z(_008_));
 CLKBUF_X2 _397_ (.A(wr_data[4]),
    .Z(_120_));
 MUX2_X1 _398_ (.A(\mem[0][4] ),
    .B(_120_),
    .S(_116_),
    .Z(_009_));
 CLKBUF_X2 _399_ (.A(wr_data[5]),
    .Z(_121_));
 MUX2_X1 _400_ (.A(\mem[0][5] ),
    .B(_121_),
    .S(_116_),
    .Z(_010_));
 CLKBUF_X2 _401_ (.A(wr_data[6]),
    .Z(_122_));
 MUX2_X1 _402_ (.A(\mem[0][6] ),
    .B(_122_),
    .S(_116_),
    .Z(_011_));
 CLKBUF_X2 _403_ (.A(wr_data[7]),
    .Z(_123_));
 MUX2_X1 _404_ (.A(\mem[0][7] ),
    .B(_123_),
    .S(_116_),
    .Z(_012_));
 NOR4_X4 _405_ (.A1(_111_),
    .A2(_112_),
    .A3(_003_),
    .A4(_115_),
    .ZN(_124_));
 MUX2_X1 _406_ (.A(\mem[1][0] ),
    .B(_110_),
    .S(_124_),
    .Z(_013_));
 MUX2_X1 _407_ (.A(\mem[1][1] ),
    .B(_117_),
    .S(_124_),
    .Z(_014_));
 MUX2_X1 _408_ (.A(\mem[1][2] ),
    .B(_118_),
    .S(_124_),
    .Z(_015_));
 MUX2_X1 _409_ (.A(\mem[1][3] ),
    .B(_119_),
    .S(_124_),
    .Z(_016_));
 MUX2_X1 _410_ (.A(\mem[1][4] ),
    .B(_120_),
    .S(_124_),
    .Z(_017_));
 MUX2_X1 _411_ (.A(\mem[1][5] ),
    .B(_121_),
    .S(_124_),
    .Z(_018_));
 MUX2_X1 _412_ (.A(\mem[1][6] ),
    .B(_122_),
    .S(_124_),
    .Z(_019_));
 MUX2_X1 _413_ (.A(\mem[1][7] ),
    .B(_123_),
    .S(_124_),
    .Z(_020_));
 INV_X1 _414_ (.A(_112_),
    .ZN(_125_));
 OR4_X1 _415_ (.A1(_111_),
    .A2(_125_),
    .A3(_113_),
    .A4(_114_),
    .ZN(_126_));
 BUF_X4 _416_ (.A(_126_),
    .Z(_127_));
 MUX2_X1 _417_ (.A(_110_),
    .B(\mem[2][0] ),
    .S(_127_),
    .Z(_021_));
 MUX2_X1 _418_ (.A(_117_),
    .B(\mem[2][1] ),
    .S(_127_),
    .Z(_022_));
 MUX2_X1 _419_ (.A(_118_),
    .B(\mem[2][2] ),
    .S(_127_),
    .Z(_023_));
 MUX2_X1 _420_ (.A(_119_),
    .B(\mem[2][3] ),
    .S(_127_),
    .Z(_024_));
 MUX2_X1 _421_ (.A(_120_),
    .B(\mem[2][4] ),
    .S(_127_),
    .Z(_025_));
 MUX2_X1 _422_ (.A(_121_),
    .B(\mem[2][5] ),
    .S(_127_),
    .Z(_026_));
 MUX2_X1 _423_ (.A(_122_),
    .B(\mem[2][6] ),
    .S(_127_),
    .Z(_027_));
 MUX2_X1 _424_ (.A(_123_),
    .B(\mem[2][7] ),
    .S(_127_),
    .Z(_028_));
 OR4_X1 _425_ (.A1(_111_),
    .A2(_125_),
    .A3(_003_),
    .A4(_114_),
    .ZN(_128_));
 CLKBUF_X3 _426_ (.A(_128_),
    .Z(_129_));
 MUX2_X1 _427_ (.A(_110_),
    .B(\mem[3][0] ),
    .S(_129_),
    .Z(_029_));
 MUX2_X1 _428_ (.A(_117_),
    .B(\mem[3][1] ),
    .S(_129_),
    .Z(_030_));
 MUX2_X1 _429_ (.A(_118_),
    .B(\mem[3][2] ),
    .S(_129_),
    .Z(_031_));
 MUX2_X1 _430_ (.A(_119_),
    .B(\mem[3][3] ),
    .S(_129_),
    .Z(_032_));
 MUX2_X1 _431_ (.A(_120_),
    .B(\mem[3][4] ),
    .S(_129_),
    .Z(_033_));
 MUX2_X1 _432_ (.A(_121_),
    .B(\mem[3][5] ),
    .S(_129_),
    .Z(_034_));
 MUX2_X1 _433_ (.A(_122_),
    .B(\mem[3][6] ),
    .S(_129_),
    .Z(_035_));
 MUX2_X1 _434_ (.A(_123_),
    .B(\mem[3][7] ),
    .S(_129_),
    .Z(_036_));
 INV_X1 _435_ (.A(_111_),
    .ZN(_130_));
 NOR4_X4 _436_ (.A1(_130_),
    .A2(_112_),
    .A3(_113_),
    .A4(_115_),
    .ZN(_131_));
 MUX2_X1 _437_ (.A(\mem[4][0] ),
    .B(_110_),
    .S(_131_),
    .Z(_037_));
 MUX2_X1 _438_ (.A(\mem[4][1] ),
    .B(_117_),
    .S(_131_),
    .Z(_038_));
 MUX2_X1 _439_ (.A(\mem[4][2] ),
    .B(_118_),
    .S(_131_),
    .Z(_039_));
 MUX2_X1 _440_ (.A(\mem[4][3] ),
    .B(_119_),
    .S(_131_),
    .Z(_040_));
 MUX2_X1 _441_ (.A(\mem[4][4] ),
    .B(_120_),
    .S(_131_),
    .Z(_041_));
 MUX2_X1 _442_ (.A(\mem[4][5] ),
    .B(_121_),
    .S(_131_),
    .Z(_042_));
 MUX2_X1 _443_ (.A(\mem[4][6] ),
    .B(_122_),
    .S(_131_),
    .Z(_043_));
 MUX2_X1 _444_ (.A(\mem[4][7] ),
    .B(_123_),
    .S(_131_),
    .Z(_044_));
 OR4_X1 _445_ (.A1(_130_),
    .A2(_112_),
    .A3(_003_),
    .A4(_114_),
    .ZN(_132_));
 CLKBUF_X3 _446_ (.A(_132_),
    .Z(_133_));
 MUX2_X1 _447_ (.A(_110_),
    .B(\mem[5][0] ),
    .S(_133_),
    .Z(_045_));
 MUX2_X1 _448_ (.A(_117_),
    .B(\mem[5][1] ),
    .S(_133_),
    .Z(_046_));
 MUX2_X1 _449_ (.A(_118_),
    .B(\mem[5][2] ),
    .S(_133_),
    .Z(_047_));
 MUX2_X1 _450_ (.A(_119_),
    .B(\mem[5][3] ),
    .S(_133_),
    .Z(_048_));
 MUX2_X1 _451_ (.A(_120_),
    .B(\mem[5][4] ),
    .S(_133_),
    .Z(_049_));
 MUX2_X1 _452_ (.A(_121_),
    .B(\mem[5][5] ),
    .S(_133_),
    .Z(_050_));
 MUX2_X1 _453_ (.A(_122_),
    .B(\mem[5][6] ),
    .S(_133_),
    .Z(_051_));
 MUX2_X1 _454_ (.A(_123_),
    .B(\mem[5][7] ),
    .S(_133_),
    .Z(_052_));
 OR4_X1 _455_ (.A1(_130_),
    .A2(_125_),
    .A3(_113_),
    .A4(_114_),
    .ZN(_134_));
 BUF_X4 _456_ (.A(_134_),
    .Z(_135_));
 MUX2_X1 _457_ (.A(_110_),
    .B(\mem[6][0] ),
    .S(_135_),
    .Z(_053_));
 MUX2_X1 _458_ (.A(_117_),
    .B(\mem[6][1] ),
    .S(_135_),
    .Z(_054_));
 MUX2_X1 _459_ (.A(_118_),
    .B(\mem[6][2] ),
    .S(_135_),
    .Z(_055_));
 MUX2_X1 _460_ (.A(_119_),
    .B(\mem[6][3] ),
    .S(_135_),
    .Z(_056_));
 MUX2_X1 _461_ (.A(_120_),
    .B(\mem[6][4] ),
    .S(_135_),
    .Z(_057_));
 MUX2_X1 _462_ (.A(_121_),
    .B(\mem[6][5] ),
    .S(_135_),
    .Z(_058_));
 MUX2_X1 _463_ (.A(_122_),
    .B(\mem[6][6] ),
    .S(_135_),
    .Z(_059_));
 MUX2_X1 _464_ (.A(_123_),
    .B(\mem[6][7] ),
    .S(_135_),
    .Z(_060_));
 NAND3_X1 _465_ (.A1(_111_),
    .A2(_112_),
    .A3(_113_),
    .ZN(_136_));
 OR2_X1 _466_ (.A1(_115_),
    .A2(_136_),
    .ZN(_137_));
 BUF_X4 _467_ (.A(_137_),
    .Z(_138_));
 MUX2_X1 _468_ (.A(_110_),
    .B(\mem[7][0] ),
    .S(_138_),
    .Z(_061_));
 MUX2_X1 _469_ (.A(_117_),
    .B(\mem[7][1] ),
    .S(_138_),
    .Z(_062_));
 MUX2_X1 _470_ (.A(_118_),
    .B(\mem[7][2] ),
    .S(_138_),
    .Z(_063_));
 MUX2_X1 _471_ (.A(_119_),
    .B(\mem[7][3] ),
    .S(_138_),
    .Z(_064_));
 MUX2_X1 _472_ (.A(_120_),
    .B(\mem[7][4] ),
    .S(_138_),
    .Z(_065_));
 MUX2_X1 _473_ (.A(_121_),
    .B(\mem[7][5] ),
    .S(_138_),
    .Z(_066_));
 MUX2_X1 _474_ (.A(_122_),
    .B(\mem[7][6] ),
    .S(_138_),
    .Z(_067_));
 MUX2_X1 _475_ (.A(_123_),
    .B(\mem[7][7] ),
    .S(_138_),
    .Z(_068_));
 CLKBUF_X3 _476_ (.A(\rd_ptr_bin[2] ),
    .Z(_139_));
 BUF_X4 _477_ (.A(_139_),
    .Z(_140_));
 MUX2_X1 _478_ (.A(\mem[3][0] ),
    .B(\mem[7][0] ),
    .S(_140_),
    .Z(_141_));
 CLKBUF_X3 _479_ (.A(\rd_ptr_bin[0] ),
    .Z(_142_));
 CLKBUF_X3 _480_ (.A(\rd_ptr_bin[1] ),
    .Z(_143_));
 NAND2_X4 _481_ (.A1(_142_),
    .A2(_143_),
    .ZN(_144_));
 BUF_X4 _482_ (.A(_139_),
    .Z(_145_));
 MUX2_X1 _483_ (.A(\mem[1][0] ),
    .B(\mem[5][0] ),
    .S(_145_),
    .Z(_146_));
 INV_X2 _484_ (.A(_143_),
    .ZN(_147_));
 NAND2_X4 _485_ (.A1(_142_),
    .A2(_147_),
    .ZN(_148_));
 OAI22_X1 _486_ (.A1(_141_),
    .A2(_144_),
    .B1(_146_),
    .B2(_148_),
    .ZN(_149_));
 MUX2_X1 _487_ (.A(\mem[2][0] ),
    .B(\mem[6][0] ),
    .S(_140_),
    .Z(_150_));
 INV_X2 _488_ (.A(_142_),
    .ZN(_151_));
 NAND2_X4 _489_ (.A1(_151_),
    .A2(_143_),
    .ZN(_152_));
 BUF_X4 _490_ (.A(_139_),
    .Z(_153_));
 MUX2_X1 _491_ (.A(\mem[0][0] ),
    .B(\mem[4][0] ),
    .S(_153_),
    .Z(_154_));
 NAND2_X4 _492_ (.A1(_151_),
    .A2(_147_),
    .ZN(_155_));
 OAI22_X1 _493_ (.A1(_150_),
    .A2(_152_),
    .B1(_154_),
    .B2(_155_),
    .ZN(_156_));
 NOR2_X1 _494_ (.A1(_149_),
    .A2(_156_),
    .ZN(_157_));
 NAND2_X2 _495_ (.A1(net2),
    .A2(_105_),
    .ZN(_158_));
 BUF_X4 _496_ (.A(_158_),
    .Z(_159_));
 MUX2_X1 _497_ (.A(_157_),
    .B(net12),
    .S(_159_),
    .Z(_069_));
 MUX2_X1 _498_ (.A(\mem[3][1] ),
    .B(\mem[7][1] ),
    .S(_140_),
    .Z(_160_));
 MUX2_X1 _499_ (.A(\mem[1][1] ),
    .B(\mem[5][1] ),
    .S(_145_),
    .Z(_161_));
 OAI22_X1 _500_ (.A1(_144_),
    .A2(_160_),
    .B1(_161_),
    .B2(_148_),
    .ZN(_162_));
 MUX2_X1 _501_ (.A(\mem[2][1] ),
    .B(\mem[6][1] ),
    .S(_145_),
    .Z(_163_));
 MUX2_X1 _502_ (.A(\mem[0][1] ),
    .B(\mem[4][1] ),
    .S(_153_),
    .Z(_164_));
 OAI22_X2 _503_ (.A1(_152_),
    .A2(_163_),
    .B1(_164_),
    .B2(_155_),
    .ZN(_165_));
 NOR2_X1 _504_ (.A1(_162_),
    .A2(_165_),
    .ZN(_166_));
 MUX2_X1 _505_ (.A(_166_),
    .B(net13),
    .S(_159_),
    .Z(_070_));
 MUX2_X1 _506_ (.A(\mem[3][2] ),
    .B(\mem[7][2] ),
    .S(_140_),
    .Z(_167_));
 MUX2_X1 _507_ (.A(\mem[1][2] ),
    .B(\mem[5][2] ),
    .S(_145_),
    .Z(_168_));
 OAI22_X1 _508_ (.A1(_144_),
    .A2(_167_),
    .B1(_168_),
    .B2(_148_),
    .ZN(_169_));
 MUX2_X1 _509_ (.A(\mem[2][2] ),
    .B(\mem[6][2] ),
    .S(_145_),
    .Z(_170_));
 MUX2_X1 _510_ (.A(\mem[0][2] ),
    .B(\mem[4][2] ),
    .S(_153_),
    .Z(_171_));
 OAI22_X1 _511_ (.A1(_152_),
    .A2(_170_),
    .B1(_171_),
    .B2(_155_),
    .ZN(_172_));
 NOR2_X1 _512_ (.A1(_169_),
    .A2(_172_),
    .ZN(_173_));
 MUX2_X1 _513_ (.A(_173_),
    .B(net14),
    .S(_159_),
    .Z(_071_));
 MUX2_X1 _514_ (.A(\mem[3][3] ),
    .B(\mem[7][3] ),
    .S(_140_),
    .Z(_174_));
 MUX2_X1 _515_ (.A(\mem[1][3] ),
    .B(\mem[5][3] ),
    .S(_145_),
    .Z(_175_));
 OAI22_X1 _516_ (.A1(_144_),
    .A2(_174_),
    .B1(_175_),
    .B2(_148_),
    .ZN(_176_));
 MUX2_X1 _517_ (.A(\mem[2][3] ),
    .B(\mem[6][3] ),
    .S(_153_),
    .Z(_177_));
 MUX2_X1 _518_ (.A(\mem[0][3] ),
    .B(\mem[4][3] ),
    .S(_153_),
    .Z(_178_));
 OAI22_X1 _519_ (.A1(_152_),
    .A2(_177_),
    .B1(_178_),
    .B2(_155_),
    .ZN(_179_));
 NOR2_X1 _520_ (.A1(_176_),
    .A2(_179_),
    .ZN(_180_));
 MUX2_X1 _521_ (.A(_180_),
    .B(net15),
    .S(_159_),
    .Z(_072_));
 MUX2_X1 _522_ (.A(\mem[3][4] ),
    .B(\mem[7][4] ),
    .S(_140_),
    .Z(_181_));
 MUX2_X1 _523_ (.A(\mem[1][4] ),
    .B(\mem[5][4] ),
    .S(_145_),
    .Z(_182_));
 OAI22_X1 _524_ (.A1(_144_),
    .A2(_181_),
    .B1(_182_),
    .B2(_148_),
    .ZN(_183_));
 MUX2_X1 _525_ (.A(\mem[2][4] ),
    .B(\mem[6][4] ),
    .S(_153_),
    .Z(_184_));
 MUX2_X1 _526_ (.A(\mem[0][4] ),
    .B(\mem[4][4] ),
    .S(_153_),
    .Z(_185_));
 OAI22_X1 _527_ (.A1(_152_),
    .A2(_184_),
    .B1(_185_),
    .B2(_155_),
    .ZN(_186_));
 NOR2_X1 _528_ (.A1(_183_),
    .A2(_186_),
    .ZN(_187_));
 MUX2_X1 _529_ (.A(_187_),
    .B(net16),
    .S(_159_),
    .Z(_073_));
 MUX2_X1 _530_ (.A(\mem[3][5] ),
    .B(\mem[7][5] ),
    .S(_140_),
    .Z(_188_));
 MUX2_X1 _531_ (.A(\mem[1][5] ),
    .B(\mem[5][5] ),
    .S(_145_),
    .Z(_189_));
 OAI22_X1 _532_ (.A1(_144_),
    .A2(_188_),
    .B1(_189_),
    .B2(_148_),
    .ZN(_190_));
 MUX2_X1 _533_ (.A(\mem[2][5] ),
    .B(\mem[6][5] ),
    .S(_153_),
    .Z(_191_));
 MUX2_X1 _534_ (.A(\mem[0][5] ),
    .B(\mem[4][5] ),
    .S(_139_),
    .Z(_192_));
 OAI22_X1 _535_ (.A1(_152_),
    .A2(_191_),
    .B1(_192_),
    .B2(_155_),
    .ZN(_193_));
 NOR2_X1 _536_ (.A1(_190_),
    .A2(_193_),
    .ZN(_194_));
 MUX2_X1 _537_ (.A(_194_),
    .B(net17),
    .S(_159_),
    .Z(_074_));
 MUX2_X1 _538_ (.A(\mem[3][6] ),
    .B(\mem[7][6] ),
    .S(_140_),
    .Z(_195_));
 MUX2_X1 _539_ (.A(\mem[1][6] ),
    .B(\mem[5][6] ),
    .S(_145_),
    .Z(_196_));
 OAI22_X1 _540_ (.A1(_144_),
    .A2(_195_),
    .B1(_196_),
    .B2(_148_),
    .ZN(_197_));
 MUX2_X1 _541_ (.A(\mem[2][6] ),
    .B(\mem[6][6] ),
    .S(_153_),
    .Z(_198_));
 MUX2_X1 _542_ (.A(\mem[0][6] ),
    .B(\mem[4][6] ),
    .S(_139_),
    .Z(_199_));
 OAI22_X1 _543_ (.A1(_152_),
    .A2(_198_),
    .B1(_199_),
    .B2(_155_),
    .ZN(_200_));
 NOR2_X1 _544_ (.A1(_197_),
    .A2(_200_),
    .ZN(_201_));
 MUX2_X1 _545_ (.A(_201_),
    .B(net18),
    .S(_159_),
    .Z(_075_));
 MUX2_X1 _546_ (.A(\mem[3][7] ),
    .B(\mem[7][7] ),
    .S(_140_),
    .Z(_202_));
 MUX2_X1 _547_ (.A(\mem[1][7] ),
    .B(\mem[5][7] ),
    .S(_145_),
    .Z(_203_));
 OAI22_X1 _548_ (.A1(_144_),
    .A2(_202_),
    .B1(_203_),
    .B2(_148_),
    .ZN(_204_));
 MUX2_X1 _549_ (.A(\mem[2][7] ),
    .B(\mem[6][7] ),
    .S(_153_),
    .Z(_205_));
 MUX2_X1 _550_ (.A(\mem[0][7] ),
    .B(\mem[4][7] ),
    .S(_139_),
    .Z(_206_));
 OAI22_X1 _551_ (.A1(_152_),
    .A2(_205_),
    .B1(_206_),
    .B2(_155_),
    .ZN(_207_));
 NOR2_X1 _552_ (.A1(_204_),
    .A2(_207_),
    .ZN(_208_));
 MUX2_X1 _553_ (.A(_208_),
    .B(net19),
    .S(_159_),
    .Z(_076_));
 MUX2_X1 _554_ (.A(_001_),
    .B(_142_),
    .S(_159_),
    .Z(_077_));
 MUX2_X1 _555_ (.A(_002_),
    .B(_143_),
    .S(_159_),
    .Z(_078_));
 XNOR2_X2 _556_ (.A(_341_),
    .B(_329_),
    .ZN(_209_));
 MUX2_X1 _557_ (.A(_209_),
    .B(_140_),
    .S(_158_),
    .Z(_079_));
 XNOR2_X1 _558_ (.A(_142_),
    .B(_002_),
    .ZN(_210_));
 MUX2_X1 _559_ (.A(_210_),
    .B(\rd_ptr_gray[0] ),
    .S(_158_),
    .Z(_080_));
 XOR2_X1 _560_ (.A(_002_),
    .B(_209_),
    .Z(_211_));
 MUX2_X1 _561_ (.A(_211_),
    .B(\rd_ptr_gray[1] ),
    .S(_158_),
    .Z(_081_));
 NAND3_X1 _562_ (.A1(_142_),
    .A2(_143_),
    .A3(_139_),
    .ZN(_212_));
 XOR2_X1 _563_ (.A(\rd_ptr_bin[3] ),
    .B(_212_),
    .Z(_213_));
 XNOR2_X1 _564_ (.A(_209_),
    .B(_213_),
    .ZN(_214_));
 MUX2_X1 _565_ (.A(_214_),
    .B(\rd_ptr_gray[2] ),
    .S(_158_),
    .Z(_082_));
 NOR2_X1 _566_ (.A1(_158_),
    .A2(_212_),
    .ZN(_215_));
 XOR2_X1 _567_ (.A(\rd_ptr_bin[3] ),
    .B(_215_),
    .Z(_083_));
 MUX2_X1 _568_ (.A(_003_),
    .B(_113_),
    .S(_115_),
    .Z(_084_));
 MUX2_X1 _569_ (.A(_004_),
    .B(_112_),
    .S(_115_),
    .Z(_085_));
 XNOR2_X2 _570_ (.A(_342_),
    .B(_000_),
    .ZN(_216_));
 MUX2_X1 _571_ (.A(_216_),
    .B(_111_),
    .S(_115_),
    .Z(_086_));
 XNOR2_X1 _572_ (.A(_113_),
    .B(_004_),
    .ZN(_217_));
 MUX2_X1 _573_ (.A(_217_),
    .B(\wr_ptr_gray[0] ),
    .S(_115_),
    .Z(_087_));
 XOR2_X1 _574_ (.A(_004_),
    .B(_216_),
    .Z(_218_));
 MUX2_X1 _575_ (.A(_218_),
    .B(\wr_ptr_gray[1] ),
    .S(_115_),
    .Z(_088_));
 XOR2_X1 _576_ (.A(\wr_ptr_bin[3] ),
    .B(_216_),
    .Z(_219_));
 XNOR2_X1 _577_ (.A(_136_),
    .B(_219_),
    .ZN(_220_));
 MUX2_X1 _578_ (.A(_220_),
    .B(\wr_ptr_gray[2] ),
    .S(_115_),
    .Z(_089_));
 XNOR2_X1 _579_ (.A(\wr_ptr_bin[3] ),
    .B(_138_),
    .ZN(_090_));
 NOR2_X1 _580_ (.A1(_323_),
    .A2(_345_),
    .ZN(_221_));
 NOR3_X1 _581_ (.A1(net10),
    .A2(net11),
    .A3(_221_),
    .ZN(net7));
 INV_X1 _582_ (.A(_323_),
    .ZN(net9));
 INV_X2 _583_ (.A(_328_),
    .ZN(net23));
 NAND2_X1 _584_ (.A1(net23),
    .A2(net24),
    .ZN(_222_));
 NAND2_X1 _585_ (.A1(_101_),
    .A2(_222_),
    .ZN(net21));
 FA_X1 _586_ (.A(_319_),
    .B(_320_),
    .CI(_321_),
    .CO(_322_),
    .S(_323_));
 FA_X1 _587_ (.A(_324_),
    .B(_325_),
    .CI(_326_),
    .CO(_327_),
    .S(_328_));
 HA_X1 _588_ (.A(_329_),
    .B(_330_),
    .CO(_331_),
    .S(_332_));
 HA_X1 _589_ (.A(_320_),
    .B(_321_),
    .CO(_333_),
    .S(_334_));
 HA_X1 _590_ (.A(\wr_ptr_bin[1] ),
    .B(_335_),
    .CO(_336_),
    .S(_337_));
 HA_X1 _591_ (.A(\wr_ptr_bin[2] ),
    .B(_338_),
    .CO(_339_),
    .S(_340_));
 HA_X1 _592_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .CO(_341_),
    .S(_002_));
 HA_X1 _593_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .CO(_342_),
    .S(_004_));
 HA_X1 _594_ (.A(\rd_ptr_bin[0] ),
    .B(_343_),
    .CO(_344_),
    .S(_345_));
 HA_X1 _595_ (.A(_346_),
    .B(_003_),
    .CO(_325_),
    .S(_347_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_005_),
    .CK(net4),
    .Q(\mem[0][0] ),
    .QN(_302_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_006_),
    .CK(net4),
    .Q(\mem[0][1] ),
    .QN(_301_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_007_),
    .CK(net4),
    .Q(\mem[0][2] ),
    .QN(_300_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_008_),
    .CK(net4),
    .Q(\mem[0][3] ),
    .QN(_299_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_009_),
    .CK(net4),
    .Q(\mem[0][4] ),
    .QN(_298_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_010_),
    .CK(net4),
    .Q(\mem[0][5] ),
    .QN(_297_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_011_),
    .CK(net4),
    .Q(\mem[0][6] ),
    .QN(_296_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_012_),
    .CK(net4),
    .Q(\mem[0][7] ),
    .QN(_295_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_013_),
    .CK(net4),
    .Q(\mem[1][0] ),
    .QN(_294_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_014_),
    .CK(net4),
    .Q(\mem[1][1] ),
    .QN(_293_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_015_),
    .CK(net4),
    .Q(\mem[1][2] ),
    .QN(_292_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_016_),
    .CK(net4),
    .Q(\mem[1][3] ),
    .QN(_291_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_017_),
    .CK(net4),
    .Q(\mem[1][4] ),
    .QN(_290_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_018_),
    .CK(net4),
    .Q(\mem[1][5] ),
    .QN(_289_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_019_),
    .CK(net4),
    .Q(\mem[1][6] ),
    .QN(_288_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_020_),
    .CK(net4),
    .Q(\mem[1][7] ),
    .QN(_287_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_021_),
    .CK(net4),
    .Q(\mem[2][0] ),
    .QN(_286_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_022_),
    .CK(net4),
    .Q(\mem[2][1] ),
    .QN(_285_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_023_),
    .CK(net4),
    .Q(\mem[2][2] ),
    .QN(_284_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_024_),
    .CK(net4),
    .Q(\mem[2][3] ),
    .QN(_283_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_025_),
    .CK(net4),
    .Q(\mem[2][4] ),
    .QN(_282_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_026_),
    .CK(net4),
    .Q(\mem[2][5] ),
    .QN(_281_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_027_),
    .CK(net4),
    .Q(\mem[2][6] ),
    .QN(_280_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_028_),
    .CK(net4),
    .Q(\mem[2][7] ),
    .QN(_279_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_029_),
    .CK(net4),
    .Q(\mem[3][0] ),
    .QN(_278_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_030_),
    .CK(net4),
    .Q(\mem[3][1] ),
    .QN(_277_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_031_),
    .CK(net4),
    .Q(\mem[3][2] ),
    .QN(_276_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_032_),
    .CK(net4),
    .Q(\mem[3][3] ),
    .QN(_275_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_033_),
    .CK(net4),
    .Q(\mem[3][4] ),
    .QN(_274_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_034_),
    .CK(net4),
    .Q(\mem[3][5] ),
    .QN(_273_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_035_),
    .CK(net4),
    .Q(\mem[3][6] ),
    .QN(_272_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_036_),
    .CK(net4),
    .Q(\mem[3][7] ),
    .QN(_271_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_037_),
    .CK(net4),
    .Q(\mem[4][0] ),
    .QN(_270_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_038_),
    .CK(net4),
    .Q(\mem[4][1] ),
    .QN(_269_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_039_),
    .CK(net4),
    .Q(\mem[4][2] ),
    .QN(_268_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_040_),
    .CK(net4),
    .Q(\mem[4][3] ),
    .QN(_267_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_041_),
    .CK(net4),
    .Q(\mem[4][4] ),
    .QN(_266_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_042_),
    .CK(net4),
    .Q(\mem[4][5] ),
    .QN(_265_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_043_),
    .CK(net4),
    .Q(\mem[4][6] ),
    .QN(_264_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_044_),
    .CK(net4),
    .Q(\mem[4][7] ),
    .QN(_263_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_045_),
    .CK(net4),
    .Q(\mem[5][0] ),
    .QN(_262_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_046_),
    .CK(net4),
    .Q(\mem[5][1] ),
    .QN(_261_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_047_),
    .CK(net4),
    .Q(\mem[5][2] ),
    .QN(_260_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_048_),
    .CK(net4),
    .Q(\mem[5][3] ),
    .QN(_259_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_049_),
    .CK(net4),
    .Q(\mem[5][4] ),
    .QN(_258_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_050_),
    .CK(net4),
    .Q(\mem[5][5] ),
    .QN(_257_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_051_),
    .CK(net4),
    .Q(\mem[5][6] ),
    .QN(_256_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_052_),
    .CK(net4),
    .Q(\mem[5][7] ),
    .QN(_255_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_053_),
    .CK(net4),
    .Q(\mem[6][0] ),
    .QN(_254_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_054_),
    .CK(net4),
    .Q(\mem[6][1] ),
    .QN(_253_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_055_),
    .CK(net4),
    .Q(\mem[6][2] ),
    .QN(_252_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_056_),
    .CK(net4),
    .Q(\mem[6][3] ),
    .QN(_251_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_057_),
    .CK(net4),
    .Q(\mem[6][4] ),
    .QN(_250_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_058_),
    .CK(net4),
    .Q(\mem[6][5] ),
    .QN(_249_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_059_),
    .CK(net4),
    .Q(\mem[6][6] ),
    .QN(_248_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_060_),
    .CK(net4),
    .Q(\mem[6][7] ),
    .QN(_247_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_061_),
    .CK(net4),
    .Q(\mem[7][0] ),
    .QN(_246_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_062_),
    .CK(net4),
    .Q(\mem[7][1] ),
    .QN(_245_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_063_),
    .CK(net4),
    .Q(\mem[7][2] ),
    .QN(_244_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_064_),
    .CK(net4),
    .Q(\mem[7][3] ),
    .QN(_243_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_065_),
    .CK(net4),
    .Q(\mem[7][4] ),
    .QN(_242_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_066_),
    .CK(net4),
    .Q(\mem[7][5] ),
    .QN(_241_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_067_),
    .CK(net4),
    .Q(\mem[7][6] ),
    .QN(_240_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_068_),
    .CK(net4),
    .Q(\mem[7][7] ),
    .QN(_239_));
 DFFR_X2 \rd_data_reg[0]$_DFFE_PN0P_  (.D(_069_),
    .RN(net3),
    .CK(net1),
    .Q(net12),
    .QN(_238_));
 DFFR_X2 \rd_data_reg[1]$_DFFE_PN0P_  (.D(_070_),
    .RN(net3),
    .CK(net1),
    .Q(net13),
    .QN(_237_));
 DFFR_X2 \rd_data_reg[2]$_DFFE_PN0P_  (.D(_071_),
    .RN(net3),
    .CK(net1),
    .Q(net14),
    .QN(_236_));
 DFFR_X2 \rd_data_reg[3]$_DFFE_PN0P_  (.D(_072_),
    .RN(net3),
    .CK(net1),
    .Q(net15),
    .QN(_235_));
 DFFR_X2 \rd_data_reg[4]$_DFFE_PN0P_  (.D(_073_),
    .RN(net3),
    .CK(net1),
    .Q(net16),
    .QN(_234_));
 DFFR_X2 \rd_data_reg[5]$_DFFE_PN0P_  (.D(_074_),
    .RN(net3),
    .CK(net1),
    .Q(net17),
    .QN(_233_));
 DFFR_X2 \rd_data_reg[6]$_DFFE_PN0P_  (.D(_075_),
    .RN(net3),
    .CK(net1),
    .Q(net18),
    .QN(_232_));
 DFFR_X2 \rd_data_reg[7]$_DFFE_PN0P_  (.D(_076_),
    .RN(net3),
    .CK(net1),
    .Q(net19),
    .QN(_231_));
 DFFR_X1 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_077_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[0] ),
    .QN(_001_));
 DFFR_X1 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_078_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[1] ),
    .QN(_321_));
 DFFR_X1 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_079_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[2] ),
    .QN(_329_));
 DFFR_X2 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_080_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[0] ),
    .QN(_230_));
 DFFR_X1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_081_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[1] ),
    .QN(_229_));
 DFFR_X1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_082_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[2] ),
    .QN(_228_));
 DFFR_X2 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_083_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[3] ),
    .QN(_303_));
 DFFR_X1 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[0] ),
    .QN(_304_));
 DFFR_X1 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[1] ),
    .QN(_305_));
 DFFR_X1 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[2] ),
    .QN(_306_));
 DFFR_X1 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_bin[3] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync1[3] ),
    .QN(_307_));
 DFFR_X2 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[0] ),
    .QN(_308_));
 DFFR_X2 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[1] ),
    .QN(_309_));
 DFFR_X2 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_gray_sync2[2] ),
    .QN(_310_));
 DFFR_X2 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .RN(net6),
    .CK(net4),
    .Q(\rd_ptr_bin_sync[3] ),
    .QN(_227_));
 DFFR_X2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_084_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[0] ),
    .QN(_003_));
 DFFR_X2 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_085_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[1] ),
    .QN(_324_));
 DFFR_X1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_086_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[2] ),
    .QN(_000_));
 DFFR_X1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_087_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[0] ),
    .QN(_226_));
 DFFR_X2 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_088_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[1] ),
    .QN(_225_));
 DFFR_X1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_089_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_gray[2] ),
    .QN(_224_));
 DFFR_X2 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_090_),
    .RN(net6),
    .CK(net4),
    .Q(\wr_ptr_bin[3] ),
    .QN(_311_));
 DFFR_X1 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[0] ),
    .QN(_312_));
 DFFR_X1 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[1] ),
    .QN(_313_));
 DFFR_X1 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[2] ),
    .QN(_314_));
 DFFR_X1 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_bin[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[3] ),
    .QN(_315_));
 DFFR_X1 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[0] ),
    .QN(_316_));
 DFFR_X2 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[1] ),
    .QN(_317_));
 DFFR_X2 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[2] ),
    .QN(_318_));
 DFFR_X1 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_bin_sync[3] ),
    .QN(_223_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Left_573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_1000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_1003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1006 ();
 BUF_X8 input1 (.A(rd_clk),
    .Z(net1));
 CLKBUF_X3 input2 (.A(rd_en),
    .Z(net2));
 BUF_X8 input3 (.A(rd_rst_n),
    .Z(net3));
 BUF_X16 input4 (.A(wr_clk),
    .Z(net4));
 BUF_X2 input5 (.A(wr_en),
    .Z(net5));
 BUF_X8 input6 (.A(wr_rst_n),
    .Z(net6));
 BUF_X1 output7 (.A(net7),
    .Z(rd_almost_empty));
 BUF_X1 output8 (.A(net8),
    .Z(rd_count[0]));
 BUF_X1 output9 (.A(net9),
    .Z(rd_count[1]));
 BUF_X1 output10 (.A(net10),
    .Z(rd_count[2]));
 BUF_X1 output11 (.A(net11),
    .Z(rd_count[3]));
 BUF_X1 output12 (.A(net12),
    .Z(rd_data[0]));
 BUF_X1 output13 (.A(net13),
    .Z(rd_data[1]));
 BUF_X1 output14 (.A(net14),
    .Z(rd_data[2]));
 BUF_X1 output15 (.A(net15),
    .Z(rd_data[3]));
 BUF_X1 output16 (.A(net16),
    .Z(rd_data[4]));
 BUF_X1 output17 (.A(net17),
    .Z(rd_data[5]));
 BUF_X1 output18 (.A(net18),
    .Z(rd_data[6]));
 BUF_X1 output19 (.A(net19),
    .Z(rd_data[7]));
 BUF_X1 output20 (.A(net20),
    .Z(rd_empty));
 BUF_X1 output21 (.A(net21),
    .Z(wr_almost_full));
 BUF_X1 output22 (.A(net22),
    .Z(wr_count[0]));
 BUF_X1 output23 (.A(net23),
    .Z(wr_count[1]));
 BUF_X1 output24 (.A(net24),
    .Z(wr_count[2]));
 BUF_X1 output25 (.A(net25),
    .Z(wr_count[3]));
 BUF_X1 output26 (.A(net26),
    .Z(wr_full));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X32 FILLER_0_856 ();
 FILLCELL_X32 FILLER_0_888 ();
 FILLCELL_X32 FILLER_0_920 ();
 FILLCELL_X32 FILLER_0_952 ();
 FILLCELL_X32 FILLER_0_984 ();
 FILLCELL_X32 FILLER_0_1016 ();
 FILLCELL_X32 FILLER_0_1048 ();
 FILLCELL_X32 FILLER_0_1080 ();
 FILLCELL_X32 FILLER_0_1112 ();
 FILLCELL_X32 FILLER_0_1144 ();
 FILLCELL_X32 FILLER_0_1176 ();
 FILLCELL_X32 FILLER_0_1208 ();
 FILLCELL_X16 FILLER_0_1240 ();
 FILLCELL_X4 FILLER_0_1256 ();
 FILLCELL_X2 FILLER_0_1260 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X32 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_0_1679 ();
 FILLCELL_X32 FILLER_0_1711 ();
 FILLCELL_X32 FILLER_0_1743 ();
 FILLCELL_X32 FILLER_0_1775 ();
 FILLCELL_X32 FILLER_0_1807 ();
 FILLCELL_X32 FILLER_0_1839 ();
 FILLCELL_X16 FILLER_0_1871 ();
 FILLCELL_X4 FILLER_0_1887 ();
 FILLCELL_X2 FILLER_0_1891 ();
 FILLCELL_X32 FILLER_0_1894 ();
 FILLCELL_X32 FILLER_0_1926 ();
 FILLCELL_X32 FILLER_0_1958 ();
 FILLCELL_X32 FILLER_0_1990 ();
 FILLCELL_X32 FILLER_0_2022 ();
 FILLCELL_X32 FILLER_0_2054 ();
 FILLCELL_X16 FILLER_0_2086 ();
 FILLCELL_X8 FILLER_0_2102 ();
 FILLCELL_X4 FILLER_0_2110 ();
 FILLCELL_X1 FILLER_0_2114 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X32 FILLER_1_801 ();
 FILLCELL_X32 FILLER_1_833 ();
 FILLCELL_X32 FILLER_1_865 ();
 FILLCELL_X32 FILLER_1_897 ();
 FILLCELL_X32 FILLER_1_929 ();
 FILLCELL_X32 FILLER_1_961 ();
 FILLCELL_X32 FILLER_1_993 ();
 FILLCELL_X32 FILLER_1_1025 ();
 FILLCELL_X32 FILLER_1_1057 ();
 FILLCELL_X32 FILLER_1_1089 ();
 FILLCELL_X32 FILLER_1_1121 ();
 FILLCELL_X32 FILLER_1_1153 ();
 FILLCELL_X32 FILLER_1_1185 ();
 FILLCELL_X32 FILLER_1_1217 ();
 FILLCELL_X8 FILLER_1_1249 ();
 FILLCELL_X4 FILLER_1_1257 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X32 FILLER_1_1648 ();
 FILLCELL_X32 FILLER_1_1680 ();
 FILLCELL_X32 FILLER_1_1712 ();
 FILLCELL_X32 FILLER_1_1744 ();
 FILLCELL_X32 FILLER_1_1776 ();
 FILLCELL_X32 FILLER_1_1808 ();
 FILLCELL_X32 FILLER_1_1840 ();
 FILLCELL_X32 FILLER_1_1872 ();
 FILLCELL_X32 FILLER_1_1904 ();
 FILLCELL_X32 FILLER_1_1936 ();
 FILLCELL_X32 FILLER_1_1968 ();
 FILLCELL_X32 FILLER_1_2000 ();
 FILLCELL_X32 FILLER_1_2032 ();
 FILLCELL_X32 FILLER_1_2064 ();
 FILLCELL_X16 FILLER_1_2096 ();
 FILLCELL_X2 FILLER_1_2112 ();
 FILLCELL_X1 FILLER_1_2114 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X32 FILLER_2_952 ();
 FILLCELL_X32 FILLER_2_984 ();
 FILLCELL_X32 FILLER_2_1016 ();
 FILLCELL_X32 FILLER_2_1048 ();
 FILLCELL_X32 FILLER_2_1080 ();
 FILLCELL_X32 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1144 ();
 FILLCELL_X32 FILLER_2_1176 ();
 FILLCELL_X32 FILLER_2_1208 ();
 FILLCELL_X32 FILLER_2_1240 ();
 FILLCELL_X32 FILLER_2_1272 ();
 FILLCELL_X32 FILLER_2_1304 ();
 FILLCELL_X32 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1368 ();
 FILLCELL_X32 FILLER_2_1400 ();
 FILLCELL_X32 FILLER_2_1432 ();
 FILLCELL_X32 FILLER_2_1464 ();
 FILLCELL_X32 FILLER_2_1496 ();
 FILLCELL_X32 FILLER_2_1528 ();
 FILLCELL_X32 FILLER_2_1560 ();
 FILLCELL_X32 FILLER_2_1592 ();
 FILLCELL_X32 FILLER_2_1624 ();
 FILLCELL_X32 FILLER_2_1656 ();
 FILLCELL_X32 FILLER_2_1688 ();
 FILLCELL_X32 FILLER_2_1720 ();
 FILLCELL_X32 FILLER_2_1752 ();
 FILLCELL_X32 FILLER_2_1784 ();
 FILLCELL_X32 FILLER_2_1816 ();
 FILLCELL_X32 FILLER_2_1848 ();
 FILLCELL_X8 FILLER_2_1880 ();
 FILLCELL_X4 FILLER_2_1888 ();
 FILLCELL_X2 FILLER_2_1892 ();
 FILLCELL_X32 FILLER_2_1895 ();
 FILLCELL_X32 FILLER_2_1927 ();
 FILLCELL_X32 FILLER_2_1959 ();
 FILLCELL_X32 FILLER_2_1991 ();
 FILLCELL_X32 FILLER_2_2023 ();
 FILLCELL_X32 FILLER_2_2055 ();
 FILLCELL_X16 FILLER_2_2087 ();
 FILLCELL_X8 FILLER_2_2103 ();
 FILLCELL_X4 FILLER_2_2111 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X32 FILLER_3_1648 ();
 FILLCELL_X32 FILLER_3_1680 ();
 FILLCELL_X32 FILLER_3_1712 ();
 FILLCELL_X32 FILLER_3_1744 ();
 FILLCELL_X32 FILLER_3_1776 ();
 FILLCELL_X32 FILLER_3_1808 ();
 FILLCELL_X32 FILLER_3_1840 ();
 FILLCELL_X32 FILLER_3_1872 ();
 FILLCELL_X32 FILLER_3_1904 ();
 FILLCELL_X32 FILLER_3_1936 ();
 FILLCELL_X32 FILLER_3_1968 ();
 FILLCELL_X32 FILLER_3_2000 ();
 FILLCELL_X32 FILLER_3_2032 ();
 FILLCELL_X32 FILLER_3_2064 ();
 FILLCELL_X16 FILLER_3_2096 ();
 FILLCELL_X2 FILLER_3_2112 ();
 FILLCELL_X1 FILLER_3_2114 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X32 FILLER_4_1304 ();
 FILLCELL_X32 FILLER_4_1336 ();
 FILLCELL_X32 FILLER_4_1368 ();
 FILLCELL_X32 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1432 ();
 FILLCELL_X32 FILLER_4_1464 ();
 FILLCELL_X32 FILLER_4_1496 ();
 FILLCELL_X32 FILLER_4_1528 ();
 FILLCELL_X32 FILLER_4_1560 ();
 FILLCELL_X32 FILLER_4_1592 ();
 FILLCELL_X32 FILLER_4_1624 ();
 FILLCELL_X32 FILLER_4_1656 ();
 FILLCELL_X32 FILLER_4_1688 ();
 FILLCELL_X32 FILLER_4_1720 ();
 FILLCELL_X32 FILLER_4_1752 ();
 FILLCELL_X32 FILLER_4_1784 ();
 FILLCELL_X32 FILLER_4_1816 ();
 FILLCELL_X32 FILLER_4_1848 ();
 FILLCELL_X8 FILLER_4_1880 ();
 FILLCELL_X4 FILLER_4_1888 ();
 FILLCELL_X2 FILLER_4_1892 ();
 FILLCELL_X32 FILLER_4_1895 ();
 FILLCELL_X32 FILLER_4_1927 ();
 FILLCELL_X32 FILLER_4_1959 ();
 FILLCELL_X32 FILLER_4_1991 ();
 FILLCELL_X32 FILLER_4_2023 ();
 FILLCELL_X32 FILLER_4_2055 ();
 FILLCELL_X16 FILLER_4_2087 ();
 FILLCELL_X8 FILLER_4_2103 ();
 FILLCELL_X4 FILLER_4_2111 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X32 FILLER_5_1648 ();
 FILLCELL_X32 FILLER_5_1680 ();
 FILLCELL_X32 FILLER_5_1712 ();
 FILLCELL_X32 FILLER_5_1744 ();
 FILLCELL_X32 FILLER_5_1776 ();
 FILLCELL_X32 FILLER_5_1808 ();
 FILLCELL_X32 FILLER_5_1840 ();
 FILLCELL_X32 FILLER_5_1872 ();
 FILLCELL_X32 FILLER_5_1904 ();
 FILLCELL_X32 FILLER_5_1936 ();
 FILLCELL_X32 FILLER_5_1968 ();
 FILLCELL_X32 FILLER_5_2000 ();
 FILLCELL_X32 FILLER_5_2032 ();
 FILLCELL_X32 FILLER_5_2064 ();
 FILLCELL_X16 FILLER_5_2096 ();
 FILLCELL_X2 FILLER_5_2112 ();
 FILLCELL_X1 FILLER_5_2114 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X32 FILLER_6_1304 ();
 FILLCELL_X32 FILLER_6_1336 ();
 FILLCELL_X32 FILLER_6_1368 ();
 FILLCELL_X32 FILLER_6_1400 ();
 FILLCELL_X32 FILLER_6_1432 ();
 FILLCELL_X32 FILLER_6_1464 ();
 FILLCELL_X32 FILLER_6_1496 ();
 FILLCELL_X32 FILLER_6_1528 ();
 FILLCELL_X32 FILLER_6_1560 ();
 FILLCELL_X32 FILLER_6_1592 ();
 FILLCELL_X32 FILLER_6_1624 ();
 FILLCELL_X32 FILLER_6_1656 ();
 FILLCELL_X32 FILLER_6_1688 ();
 FILLCELL_X32 FILLER_6_1720 ();
 FILLCELL_X32 FILLER_6_1752 ();
 FILLCELL_X32 FILLER_6_1784 ();
 FILLCELL_X32 FILLER_6_1816 ();
 FILLCELL_X32 FILLER_6_1848 ();
 FILLCELL_X8 FILLER_6_1880 ();
 FILLCELL_X4 FILLER_6_1888 ();
 FILLCELL_X2 FILLER_6_1892 ();
 FILLCELL_X32 FILLER_6_1895 ();
 FILLCELL_X32 FILLER_6_1927 ();
 FILLCELL_X32 FILLER_6_1959 ();
 FILLCELL_X32 FILLER_6_1991 ();
 FILLCELL_X32 FILLER_6_2023 ();
 FILLCELL_X32 FILLER_6_2055 ();
 FILLCELL_X16 FILLER_6_2087 ();
 FILLCELL_X8 FILLER_6_2103 ();
 FILLCELL_X4 FILLER_6_2111 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X32 FILLER_7_1648 ();
 FILLCELL_X32 FILLER_7_1680 ();
 FILLCELL_X32 FILLER_7_1712 ();
 FILLCELL_X32 FILLER_7_1744 ();
 FILLCELL_X32 FILLER_7_1776 ();
 FILLCELL_X32 FILLER_7_1808 ();
 FILLCELL_X32 FILLER_7_1840 ();
 FILLCELL_X32 FILLER_7_1872 ();
 FILLCELL_X32 FILLER_7_1904 ();
 FILLCELL_X32 FILLER_7_1936 ();
 FILLCELL_X32 FILLER_7_1968 ();
 FILLCELL_X32 FILLER_7_2000 ();
 FILLCELL_X32 FILLER_7_2032 ();
 FILLCELL_X32 FILLER_7_2064 ();
 FILLCELL_X16 FILLER_7_2096 ();
 FILLCELL_X2 FILLER_7_2112 ();
 FILLCELL_X1 FILLER_7_2114 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X32 FILLER_8_1304 ();
 FILLCELL_X32 FILLER_8_1336 ();
 FILLCELL_X32 FILLER_8_1368 ();
 FILLCELL_X32 FILLER_8_1400 ();
 FILLCELL_X32 FILLER_8_1432 ();
 FILLCELL_X32 FILLER_8_1464 ();
 FILLCELL_X32 FILLER_8_1496 ();
 FILLCELL_X32 FILLER_8_1528 ();
 FILLCELL_X32 FILLER_8_1560 ();
 FILLCELL_X32 FILLER_8_1592 ();
 FILLCELL_X32 FILLER_8_1624 ();
 FILLCELL_X32 FILLER_8_1656 ();
 FILLCELL_X32 FILLER_8_1688 ();
 FILLCELL_X32 FILLER_8_1720 ();
 FILLCELL_X32 FILLER_8_1752 ();
 FILLCELL_X32 FILLER_8_1784 ();
 FILLCELL_X32 FILLER_8_1816 ();
 FILLCELL_X32 FILLER_8_1848 ();
 FILLCELL_X8 FILLER_8_1880 ();
 FILLCELL_X4 FILLER_8_1888 ();
 FILLCELL_X2 FILLER_8_1892 ();
 FILLCELL_X32 FILLER_8_1895 ();
 FILLCELL_X32 FILLER_8_1927 ();
 FILLCELL_X32 FILLER_8_1959 ();
 FILLCELL_X32 FILLER_8_1991 ();
 FILLCELL_X32 FILLER_8_2023 ();
 FILLCELL_X32 FILLER_8_2055 ();
 FILLCELL_X16 FILLER_8_2087 ();
 FILLCELL_X8 FILLER_8_2103 ();
 FILLCELL_X4 FILLER_8_2111 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X32 FILLER_9_1648 ();
 FILLCELL_X32 FILLER_9_1680 ();
 FILLCELL_X32 FILLER_9_1712 ();
 FILLCELL_X32 FILLER_9_1744 ();
 FILLCELL_X32 FILLER_9_1776 ();
 FILLCELL_X32 FILLER_9_1808 ();
 FILLCELL_X32 FILLER_9_1840 ();
 FILLCELL_X32 FILLER_9_1872 ();
 FILLCELL_X32 FILLER_9_1904 ();
 FILLCELL_X32 FILLER_9_1936 ();
 FILLCELL_X32 FILLER_9_1968 ();
 FILLCELL_X32 FILLER_9_2000 ();
 FILLCELL_X32 FILLER_9_2032 ();
 FILLCELL_X32 FILLER_9_2064 ();
 FILLCELL_X16 FILLER_9_2096 ();
 FILLCELL_X2 FILLER_9_2112 ();
 FILLCELL_X1 FILLER_9_2114 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X32 FILLER_10_1304 ();
 FILLCELL_X32 FILLER_10_1336 ();
 FILLCELL_X32 FILLER_10_1368 ();
 FILLCELL_X32 FILLER_10_1400 ();
 FILLCELL_X32 FILLER_10_1432 ();
 FILLCELL_X32 FILLER_10_1464 ();
 FILLCELL_X32 FILLER_10_1496 ();
 FILLCELL_X32 FILLER_10_1528 ();
 FILLCELL_X32 FILLER_10_1560 ();
 FILLCELL_X32 FILLER_10_1592 ();
 FILLCELL_X32 FILLER_10_1624 ();
 FILLCELL_X32 FILLER_10_1656 ();
 FILLCELL_X32 FILLER_10_1688 ();
 FILLCELL_X32 FILLER_10_1720 ();
 FILLCELL_X32 FILLER_10_1752 ();
 FILLCELL_X32 FILLER_10_1784 ();
 FILLCELL_X32 FILLER_10_1816 ();
 FILLCELL_X32 FILLER_10_1848 ();
 FILLCELL_X8 FILLER_10_1880 ();
 FILLCELL_X4 FILLER_10_1888 ();
 FILLCELL_X2 FILLER_10_1892 ();
 FILLCELL_X32 FILLER_10_1895 ();
 FILLCELL_X32 FILLER_10_1927 ();
 FILLCELL_X32 FILLER_10_1959 ();
 FILLCELL_X32 FILLER_10_1991 ();
 FILLCELL_X32 FILLER_10_2023 ();
 FILLCELL_X32 FILLER_10_2055 ();
 FILLCELL_X16 FILLER_10_2087 ();
 FILLCELL_X8 FILLER_10_2103 ();
 FILLCELL_X4 FILLER_10_2111 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X32 FILLER_11_1648 ();
 FILLCELL_X32 FILLER_11_1680 ();
 FILLCELL_X32 FILLER_11_1712 ();
 FILLCELL_X32 FILLER_11_1744 ();
 FILLCELL_X32 FILLER_11_1776 ();
 FILLCELL_X32 FILLER_11_1808 ();
 FILLCELL_X32 FILLER_11_1840 ();
 FILLCELL_X32 FILLER_11_1872 ();
 FILLCELL_X32 FILLER_11_1904 ();
 FILLCELL_X32 FILLER_11_1936 ();
 FILLCELL_X32 FILLER_11_1968 ();
 FILLCELL_X32 FILLER_11_2000 ();
 FILLCELL_X32 FILLER_11_2032 ();
 FILLCELL_X32 FILLER_11_2064 ();
 FILLCELL_X16 FILLER_11_2096 ();
 FILLCELL_X2 FILLER_11_2112 ();
 FILLCELL_X1 FILLER_11_2114 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X32 FILLER_12_1592 ();
 FILLCELL_X32 FILLER_12_1624 ();
 FILLCELL_X32 FILLER_12_1656 ();
 FILLCELL_X32 FILLER_12_1688 ();
 FILLCELL_X32 FILLER_12_1720 ();
 FILLCELL_X32 FILLER_12_1752 ();
 FILLCELL_X32 FILLER_12_1784 ();
 FILLCELL_X32 FILLER_12_1816 ();
 FILLCELL_X32 FILLER_12_1848 ();
 FILLCELL_X8 FILLER_12_1880 ();
 FILLCELL_X4 FILLER_12_1888 ();
 FILLCELL_X2 FILLER_12_1892 ();
 FILLCELL_X32 FILLER_12_1895 ();
 FILLCELL_X32 FILLER_12_1927 ();
 FILLCELL_X32 FILLER_12_1959 ();
 FILLCELL_X32 FILLER_12_1991 ();
 FILLCELL_X32 FILLER_12_2023 ();
 FILLCELL_X32 FILLER_12_2055 ();
 FILLCELL_X16 FILLER_12_2087 ();
 FILLCELL_X8 FILLER_12_2103 ();
 FILLCELL_X4 FILLER_12_2111 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X32 FILLER_13_1648 ();
 FILLCELL_X32 FILLER_13_1680 ();
 FILLCELL_X32 FILLER_13_1712 ();
 FILLCELL_X32 FILLER_13_1744 ();
 FILLCELL_X32 FILLER_13_1776 ();
 FILLCELL_X32 FILLER_13_1808 ();
 FILLCELL_X32 FILLER_13_1840 ();
 FILLCELL_X32 FILLER_13_1872 ();
 FILLCELL_X32 FILLER_13_1904 ();
 FILLCELL_X32 FILLER_13_1936 ();
 FILLCELL_X32 FILLER_13_1968 ();
 FILLCELL_X32 FILLER_13_2000 ();
 FILLCELL_X32 FILLER_13_2032 ();
 FILLCELL_X32 FILLER_13_2064 ();
 FILLCELL_X16 FILLER_13_2096 ();
 FILLCELL_X2 FILLER_13_2112 ();
 FILLCELL_X1 FILLER_13_2114 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X32 FILLER_14_1688 ();
 FILLCELL_X32 FILLER_14_1720 ();
 FILLCELL_X32 FILLER_14_1752 ();
 FILLCELL_X32 FILLER_14_1784 ();
 FILLCELL_X32 FILLER_14_1816 ();
 FILLCELL_X32 FILLER_14_1848 ();
 FILLCELL_X8 FILLER_14_1880 ();
 FILLCELL_X4 FILLER_14_1888 ();
 FILLCELL_X2 FILLER_14_1892 ();
 FILLCELL_X32 FILLER_14_1895 ();
 FILLCELL_X32 FILLER_14_1927 ();
 FILLCELL_X32 FILLER_14_1959 ();
 FILLCELL_X32 FILLER_14_1991 ();
 FILLCELL_X32 FILLER_14_2023 ();
 FILLCELL_X32 FILLER_14_2055 ();
 FILLCELL_X16 FILLER_14_2087 ();
 FILLCELL_X8 FILLER_14_2103 ();
 FILLCELL_X4 FILLER_14_2111 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X32 FILLER_15_1584 ();
 FILLCELL_X32 FILLER_15_1616 ();
 FILLCELL_X32 FILLER_15_1648 ();
 FILLCELL_X32 FILLER_15_1680 ();
 FILLCELL_X32 FILLER_15_1712 ();
 FILLCELL_X32 FILLER_15_1744 ();
 FILLCELL_X32 FILLER_15_1776 ();
 FILLCELL_X32 FILLER_15_1808 ();
 FILLCELL_X32 FILLER_15_1840 ();
 FILLCELL_X32 FILLER_15_1872 ();
 FILLCELL_X32 FILLER_15_1904 ();
 FILLCELL_X32 FILLER_15_1936 ();
 FILLCELL_X32 FILLER_15_1968 ();
 FILLCELL_X32 FILLER_15_2000 ();
 FILLCELL_X32 FILLER_15_2032 ();
 FILLCELL_X32 FILLER_15_2064 ();
 FILLCELL_X16 FILLER_15_2096 ();
 FILLCELL_X2 FILLER_15_2112 ();
 FILLCELL_X1 FILLER_15_2114 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X32 FILLER_16_1592 ();
 FILLCELL_X32 FILLER_16_1624 ();
 FILLCELL_X32 FILLER_16_1656 ();
 FILLCELL_X32 FILLER_16_1688 ();
 FILLCELL_X32 FILLER_16_1720 ();
 FILLCELL_X32 FILLER_16_1752 ();
 FILLCELL_X32 FILLER_16_1784 ();
 FILLCELL_X32 FILLER_16_1816 ();
 FILLCELL_X32 FILLER_16_1848 ();
 FILLCELL_X8 FILLER_16_1880 ();
 FILLCELL_X4 FILLER_16_1888 ();
 FILLCELL_X2 FILLER_16_1892 ();
 FILLCELL_X32 FILLER_16_1895 ();
 FILLCELL_X32 FILLER_16_1927 ();
 FILLCELL_X32 FILLER_16_1959 ();
 FILLCELL_X32 FILLER_16_1991 ();
 FILLCELL_X32 FILLER_16_2023 ();
 FILLCELL_X32 FILLER_16_2055 ();
 FILLCELL_X16 FILLER_16_2087 ();
 FILLCELL_X8 FILLER_16_2103 ();
 FILLCELL_X4 FILLER_16_2111 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X32 FILLER_17_1584 ();
 FILLCELL_X32 FILLER_17_1616 ();
 FILLCELL_X32 FILLER_17_1648 ();
 FILLCELL_X32 FILLER_17_1680 ();
 FILLCELL_X32 FILLER_17_1712 ();
 FILLCELL_X32 FILLER_17_1744 ();
 FILLCELL_X32 FILLER_17_1776 ();
 FILLCELL_X32 FILLER_17_1808 ();
 FILLCELL_X32 FILLER_17_1840 ();
 FILLCELL_X32 FILLER_17_1872 ();
 FILLCELL_X32 FILLER_17_1904 ();
 FILLCELL_X32 FILLER_17_1936 ();
 FILLCELL_X32 FILLER_17_1968 ();
 FILLCELL_X32 FILLER_17_2000 ();
 FILLCELL_X32 FILLER_17_2032 ();
 FILLCELL_X32 FILLER_17_2064 ();
 FILLCELL_X16 FILLER_17_2096 ();
 FILLCELL_X2 FILLER_17_2112 ();
 FILLCELL_X1 FILLER_17_2114 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X32 FILLER_18_1752 ();
 FILLCELL_X32 FILLER_18_1784 ();
 FILLCELL_X32 FILLER_18_1816 ();
 FILLCELL_X32 FILLER_18_1848 ();
 FILLCELL_X8 FILLER_18_1880 ();
 FILLCELL_X4 FILLER_18_1888 ();
 FILLCELL_X2 FILLER_18_1892 ();
 FILLCELL_X32 FILLER_18_1895 ();
 FILLCELL_X32 FILLER_18_1927 ();
 FILLCELL_X32 FILLER_18_1959 ();
 FILLCELL_X32 FILLER_18_1991 ();
 FILLCELL_X32 FILLER_18_2023 ();
 FILLCELL_X32 FILLER_18_2055 ();
 FILLCELL_X16 FILLER_18_2087 ();
 FILLCELL_X8 FILLER_18_2103 ();
 FILLCELL_X4 FILLER_18_2111 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X32 FILLER_19_1584 ();
 FILLCELL_X32 FILLER_19_1616 ();
 FILLCELL_X32 FILLER_19_1648 ();
 FILLCELL_X32 FILLER_19_1680 ();
 FILLCELL_X32 FILLER_19_1712 ();
 FILLCELL_X32 FILLER_19_1744 ();
 FILLCELL_X32 FILLER_19_1776 ();
 FILLCELL_X32 FILLER_19_1808 ();
 FILLCELL_X32 FILLER_19_1840 ();
 FILLCELL_X32 FILLER_19_1872 ();
 FILLCELL_X32 FILLER_19_1904 ();
 FILLCELL_X32 FILLER_19_1936 ();
 FILLCELL_X32 FILLER_19_1968 ();
 FILLCELL_X32 FILLER_19_2000 ();
 FILLCELL_X32 FILLER_19_2032 ();
 FILLCELL_X32 FILLER_19_2064 ();
 FILLCELL_X16 FILLER_19_2096 ();
 FILLCELL_X2 FILLER_19_2112 ();
 FILLCELL_X1 FILLER_19_2114 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X32 FILLER_20_1592 ();
 FILLCELL_X32 FILLER_20_1624 ();
 FILLCELL_X32 FILLER_20_1656 ();
 FILLCELL_X32 FILLER_20_1688 ();
 FILLCELL_X32 FILLER_20_1720 ();
 FILLCELL_X32 FILLER_20_1752 ();
 FILLCELL_X32 FILLER_20_1784 ();
 FILLCELL_X32 FILLER_20_1816 ();
 FILLCELL_X32 FILLER_20_1848 ();
 FILLCELL_X8 FILLER_20_1880 ();
 FILLCELL_X4 FILLER_20_1888 ();
 FILLCELL_X2 FILLER_20_1892 ();
 FILLCELL_X32 FILLER_20_1895 ();
 FILLCELL_X32 FILLER_20_1927 ();
 FILLCELL_X32 FILLER_20_1959 ();
 FILLCELL_X32 FILLER_20_1991 ();
 FILLCELL_X32 FILLER_20_2023 ();
 FILLCELL_X32 FILLER_20_2055 ();
 FILLCELL_X16 FILLER_20_2087 ();
 FILLCELL_X8 FILLER_20_2103 ();
 FILLCELL_X4 FILLER_20_2111 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X32 FILLER_21_1744 ();
 FILLCELL_X32 FILLER_21_1776 ();
 FILLCELL_X32 FILLER_21_1808 ();
 FILLCELL_X32 FILLER_21_1840 ();
 FILLCELL_X32 FILLER_21_1872 ();
 FILLCELL_X32 FILLER_21_1904 ();
 FILLCELL_X32 FILLER_21_1936 ();
 FILLCELL_X32 FILLER_21_1968 ();
 FILLCELL_X32 FILLER_21_2000 ();
 FILLCELL_X32 FILLER_21_2032 ();
 FILLCELL_X32 FILLER_21_2064 ();
 FILLCELL_X16 FILLER_21_2096 ();
 FILLCELL_X2 FILLER_21_2112 ();
 FILLCELL_X1 FILLER_21_2114 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X32 FILLER_22_1752 ();
 FILLCELL_X32 FILLER_22_1784 ();
 FILLCELL_X32 FILLER_22_1816 ();
 FILLCELL_X32 FILLER_22_1848 ();
 FILLCELL_X8 FILLER_22_1880 ();
 FILLCELL_X4 FILLER_22_1888 ();
 FILLCELL_X2 FILLER_22_1892 ();
 FILLCELL_X32 FILLER_22_1895 ();
 FILLCELL_X32 FILLER_22_1927 ();
 FILLCELL_X32 FILLER_22_1959 ();
 FILLCELL_X32 FILLER_22_1991 ();
 FILLCELL_X32 FILLER_22_2023 ();
 FILLCELL_X32 FILLER_22_2055 ();
 FILLCELL_X16 FILLER_22_2087 ();
 FILLCELL_X8 FILLER_22_2103 ();
 FILLCELL_X4 FILLER_22_2111 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X32 FILLER_23_1584 ();
 FILLCELL_X32 FILLER_23_1616 ();
 FILLCELL_X32 FILLER_23_1648 ();
 FILLCELL_X32 FILLER_23_1680 ();
 FILLCELL_X32 FILLER_23_1712 ();
 FILLCELL_X32 FILLER_23_1744 ();
 FILLCELL_X32 FILLER_23_1776 ();
 FILLCELL_X32 FILLER_23_1808 ();
 FILLCELL_X32 FILLER_23_1840 ();
 FILLCELL_X32 FILLER_23_1872 ();
 FILLCELL_X32 FILLER_23_1904 ();
 FILLCELL_X32 FILLER_23_1936 ();
 FILLCELL_X32 FILLER_23_1968 ();
 FILLCELL_X32 FILLER_23_2000 ();
 FILLCELL_X32 FILLER_23_2032 ();
 FILLCELL_X32 FILLER_23_2064 ();
 FILLCELL_X16 FILLER_23_2096 ();
 FILLCELL_X2 FILLER_23_2112 ();
 FILLCELL_X1 FILLER_23_2114 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X32 FILLER_24_1592 ();
 FILLCELL_X32 FILLER_24_1624 ();
 FILLCELL_X32 FILLER_24_1656 ();
 FILLCELL_X32 FILLER_24_1688 ();
 FILLCELL_X32 FILLER_24_1720 ();
 FILLCELL_X32 FILLER_24_1752 ();
 FILLCELL_X32 FILLER_24_1784 ();
 FILLCELL_X32 FILLER_24_1816 ();
 FILLCELL_X32 FILLER_24_1848 ();
 FILLCELL_X8 FILLER_24_1880 ();
 FILLCELL_X4 FILLER_24_1888 ();
 FILLCELL_X2 FILLER_24_1892 ();
 FILLCELL_X32 FILLER_24_1895 ();
 FILLCELL_X32 FILLER_24_1927 ();
 FILLCELL_X32 FILLER_24_1959 ();
 FILLCELL_X32 FILLER_24_1991 ();
 FILLCELL_X32 FILLER_24_2023 ();
 FILLCELL_X32 FILLER_24_2055 ();
 FILLCELL_X16 FILLER_24_2087 ();
 FILLCELL_X8 FILLER_24_2103 ();
 FILLCELL_X4 FILLER_24_2111 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X32 FILLER_25_1584 ();
 FILLCELL_X32 FILLER_25_1616 ();
 FILLCELL_X32 FILLER_25_1648 ();
 FILLCELL_X32 FILLER_25_1680 ();
 FILLCELL_X32 FILLER_25_1712 ();
 FILLCELL_X32 FILLER_25_1744 ();
 FILLCELL_X32 FILLER_25_1776 ();
 FILLCELL_X32 FILLER_25_1808 ();
 FILLCELL_X32 FILLER_25_1840 ();
 FILLCELL_X32 FILLER_25_1872 ();
 FILLCELL_X32 FILLER_25_1904 ();
 FILLCELL_X32 FILLER_25_1936 ();
 FILLCELL_X32 FILLER_25_1968 ();
 FILLCELL_X32 FILLER_25_2000 ();
 FILLCELL_X32 FILLER_25_2032 ();
 FILLCELL_X32 FILLER_25_2064 ();
 FILLCELL_X16 FILLER_25_2096 ();
 FILLCELL_X2 FILLER_25_2112 ();
 FILLCELL_X1 FILLER_25_2114 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X32 FILLER_26_1592 ();
 FILLCELL_X32 FILLER_26_1624 ();
 FILLCELL_X32 FILLER_26_1656 ();
 FILLCELL_X32 FILLER_26_1688 ();
 FILLCELL_X32 FILLER_26_1720 ();
 FILLCELL_X32 FILLER_26_1752 ();
 FILLCELL_X32 FILLER_26_1784 ();
 FILLCELL_X32 FILLER_26_1816 ();
 FILLCELL_X32 FILLER_26_1848 ();
 FILLCELL_X8 FILLER_26_1880 ();
 FILLCELL_X4 FILLER_26_1888 ();
 FILLCELL_X2 FILLER_26_1892 ();
 FILLCELL_X32 FILLER_26_1895 ();
 FILLCELL_X32 FILLER_26_1927 ();
 FILLCELL_X32 FILLER_26_1959 ();
 FILLCELL_X32 FILLER_26_1991 ();
 FILLCELL_X32 FILLER_26_2023 ();
 FILLCELL_X32 FILLER_26_2055 ();
 FILLCELL_X16 FILLER_26_2087 ();
 FILLCELL_X8 FILLER_26_2103 ();
 FILLCELL_X4 FILLER_26_2111 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X32 FILLER_27_1584 ();
 FILLCELL_X32 FILLER_27_1616 ();
 FILLCELL_X32 FILLER_27_1648 ();
 FILLCELL_X32 FILLER_27_1680 ();
 FILLCELL_X32 FILLER_27_1712 ();
 FILLCELL_X32 FILLER_27_1744 ();
 FILLCELL_X32 FILLER_27_1776 ();
 FILLCELL_X32 FILLER_27_1808 ();
 FILLCELL_X32 FILLER_27_1840 ();
 FILLCELL_X32 FILLER_27_1872 ();
 FILLCELL_X32 FILLER_27_1904 ();
 FILLCELL_X32 FILLER_27_1936 ();
 FILLCELL_X32 FILLER_27_1968 ();
 FILLCELL_X32 FILLER_27_2000 ();
 FILLCELL_X32 FILLER_27_2032 ();
 FILLCELL_X32 FILLER_27_2064 ();
 FILLCELL_X16 FILLER_27_2096 ();
 FILLCELL_X2 FILLER_27_2112 ();
 FILLCELL_X1 FILLER_27_2114 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X32 FILLER_28_1592 ();
 FILLCELL_X32 FILLER_28_1624 ();
 FILLCELL_X32 FILLER_28_1656 ();
 FILLCELL_X32 FILLER_28_1688 ();
 FILLCELL_X32 FILLER_28_1720 ();
 FILLCELL_X32 FILLER_28_1752 ();
 FILLCELL_X32 FILLER_28_1784 ();
 FILLCELL_X32 FILLER_28_1816 ();
 FILLCELL_X32 FILLER_28_1848 ();
 FILLCELL_X8 FILLER_28_1880 ();
 FILLCELL_X4 FILLER_28_1888 ();
 FILLCELL_X2 FILLER_28_1892 ();
 FILLCELL_X32 FILLER_28_1895 ();
 FILLCELL_X32 FILLER_28_1927 ();
 FILLCELL_X32 FILLER_28_1959 ();
 FILLCELL_X32 FILLER_28_1991 ();
 FILLCELL_X32 FILLER_28_2023 ();
 FILLCELL_X32 FILLER_28_2055 ();
 FILLCELL_X16 FILLER_28_2087 ();
 FILLCELL_X8 FILLER_28_2103 ();
 FILLCELL_X4 FILLER_28_2111 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X32 FILLER_29_1584 ();
 FILLCELL_X32 FILLER_29_1616 ();
 FILLCELL_X32 FILLER_29_1648 ();
 FILLCELL_X32 FILLER_29_1680 ();
 FILLCELL_X32 FILLER_29_1712 ();
 FILLCELL_X32 FILLER_29_1744 ();
 FILLCELL_X32 FILLER_29_1776 ();
 FILLCELL_X32 FILLER_29_1808 ();
 FILLCELL_X32 FILLER_29_1840 ();
 FILLCELL_X32 FILLER_29_1872 ();
 FILLCELL_X32 FILLER_29_1904 ();
 FILLCELL_X32 FILLER_29_1936 ();
 FILLCELL_X32 FILLER_29_1968 ();
 FILLCELL_X32 FILLER_29_2000 ();
 FILLCELL_X32 FILLER_29_2032 ();
 FILLCELL_X32 FILLER_29_2064 ();
 FILLCELL_X16 FILLER_29_2096 ();
 FILLCELL_X2 FILLER_29_2112 ();
 FILLCELL_X1 FILLER_29_2114 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X32 FILLER_30_1592 ();
 FILLCELL_X32 FILLER_30_1624 ();
 FILLCELL_X32 FILLER_30_1656 ();
 FILLCELL_X32 FILLER_30_1688 ();
 FILLCELL_X32 FILLER_30_1720 ();
 FILLCELL_X32 FILLER_30_1752 ();
 FILLCELL_X32 FILLER_30_1784 ();
 FILLCELL_X32 FILLER_30_1816 ();
 FILLCELL_X32 FILLER_30_1848 ();
 FILLCELL_X8 FILLER_30_1880 ();
 FILLCELL_X4 FILLER_30_1888 ();
 FILLCELL_X2 FILLER_30_1892 ();
 FILLCELL_X32 FILLER_30_1895 ();
 FILLCELL_X32 FILLER_30_1927 ();
 FILLCELL_X32 FILLER_30_1959 ();
 FILLCELL_X32 FILLER_30_1991 ();
 FILLCELL_X32 FILLER_30_2023 ();
 FILLCELL_X32 FILLER_30_2055 ();
 FILLCELL_X16 FILLER_30_2087 ();
 FILLCELL_X8 FILLER_30_2103 ();
 FILLCELL_X4 FILLER_30_2111 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X32 FILLER_31_1584 ();
 FILLCELL_X32 FILLER_31_1616 ();
 FILLCELL_X32 FILLER_31_1648 ();
 FILLCELL_X32 FILLER_31_1680 ();
 FILLCELL_X32 FILLER_31_1712 ();
 FILLCELL_X32 FILLER_31_1744 ();
 FILLCELL_X32 FILLER_31_1776 ();
 FILLCELL_X32 FILLER_31_1808 ();
 FILLCELL_X32 FILLER_31_1840 ();
 FILLCELL_X32 FILLER_31_1872 ();
 FILLCELL_X32 FILLER_31_1904 ();
 FILLCELL_X32 FILLER_31_1936 ();
 FILLCELL_X32 FILLER_31_1968 ();
 FILLCELL_X32 FILLER_31_2000 ();
 FILLCELL_X32 FILLER_31_2032 ();
 FILLCELL_X32 FILLER_31_2064 ();
 FILLCELL_X16 FILLER_31_2096 ();
 FILLCELL_X2 FILLER_31_2112 ();
 FILLCELL_X1 FILLER_31_2114 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X32 FILLER_32_1592 ();
 FILLCELL_X32 FILLER_32_1624 ();
 FILLCELL_X32 FILLER_32_1656 ();
 FILLCELL_X32 FILLER_32_1688 ();
 FILLCELL_X32 FILLER_32_1720 ();
 FILLCELL_X32 FILLER_32_1752 ();
 FILLCELL_X32 FILLER_32_1784 ();
 FILLCELL_X32 FILLER_32_1816 ();
 FILLCELL_X32 FILLER_32_1848 ();
 FILLCELL_X8 FILLER_32_1880 ();
 FILLCELL_X4 FILLER_32_1888 ();
 FILLCELL_X2 FILLER_32_1892 ();
 FILLCELL_X32 FILLER_32_1895 ();
 FILLCELL_X32 FILLER_32_1927 ();
 FILLCELL_X32 FILLER_32_1959 ();
 FILLCELL_X32 FILLER_32_1991 ();
 FILLCELL_X32 FILLER_32_2023 ();
 FILLCELL_X32 FILLER_32_2055 ();
 FILLCELL_X16 FILLER_32_2087 ();
 FILLCELL_X8 FILLER_32_2103 ();
 FILLCELL_X4 FILLER_32_2111 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X32 FILLER_33_1584 ();
 FILLCELL_X32 FILLER_33_1616 ();
 FILLCELL_X32 FILLER_33_1648 ();
 FILLCELL_X32 FILLER_33_1680 ();
 FILLCELL_X32 FILLER_33_1712 ();
 FILLCELL_X32 FILLER_33_1744 ();
 FILLCELL_X32 FILLER_33_1776 ();
 FILLCELL_X32 FILLER_33_1808 ();
 FILLCELL_X32 FILLER_33_1840 ();
 FILLCELL_X32 FILLER_33_1872 ();
 FILLCELL_X32 FILLER_33_1904 ();
 FILLCELL_X32 FILLER_33_1936 ();
 FILLCELL_X32 FILLER_33_1968 ();
 FILLCELL_X32 FILLER_33_2000 ();
 FILLCELL_X32 FILLER_33_2032 ();
 FILLCELL_X32 FILLER_33_2064 ();
 FILLCELL_X16 FILLER_33_2096 ();
 FILLCELL_X2 FILLER_33_2112 ();
 FILLCELL_X1 FILLER_33_2114 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X32 FILLER_34_1592 ();
 FILLCELL_X32 FILLER_34_1624 ();
 FILLCELL_X32 FILLER_34_1656 ();
 FILLCELL_X32 FILLER_34_1688 ();
 FILLCELL_X32 FILLER_34_1720 ();
 FILLCELL_X32 FILLER_34_1752 ();
 FILLCELL_X32 FILLER_34_1784 ();
 FILLCELL_X32 FILLER_34_1816 ();
 FILLCELL_X32 FILLER_34_1848 ();
 FILLCELL_X8 FILLER_34_1880 ();
 FILLCELL_X4 FILLER_34_1888 ();
 FILLCELL_X2 FILLER_34_1892 ();
 FILLCELL_X32 FILLER_34_1895 ();
 FILLCELL_X32 FILLER_34_1927 ();
 FILLCELL_X32 FILLER_34_1959 ();
 FILLCELL_X32 FILLER_34_1991 ();
 FILLCELL_X32 FILLER_34_2023 ();
 FILLCELL_X32 FILLER_34_2055 ();
 FILLCELL_X16 FILLER_34_2087 ();
 FILLCELL_X8 FILLER_34_2103 ();
 FILLCELL_X4 FILLER_34_2111 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X32 FILLER_35_1584 ();
 FILLCELL_X32 FILLER_35_1616 ();
 FILLCELL_X32 FILLER_35_1648 ();
 FILLCELL_X32 FILLER_35_1680 ();
 FILLCELL_X32 FILLER_35_1712 ();
 FILLCELL_X32 FILLER_35_1744 ();
 FILLCELL_X32 FILLER_35_1776 ();
 FILLCELL_X32 FILLER_35_1808 ();
 FILLCELL_X32 FILLER_35_1840 ();
 FILLCELL_X32 FILLER_35_1872 ();
 FILLCELL_X32 FILLER_35_1904 ();
 FILLCELL_X32 FILLER_35_1936 ();
 FILLCELL_X32 FILLER_35_1968 ();
 FILLCELL_X32 FILLER_35_2000 ();
 FILLCELL_X32 FILLER_35_2032 ();
 FILLCELL_X32 FILLER_35_2064 ();
 FILLCELL_X16 FILLER_35_2096 ();
 FILLCELL_X2 FILLER_35_2112 ();
 FILLCELL_X1 FILLER_35_2114 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X32 FILLER_36_1592 ();
 FILLCELL_X32 FILLER_36_1624 ();
 FILLCELL_X32 FILLER_36_1656 ();
 FILLCELL_X32 FILLER_36_1688 ();
 FILLCELL_X32 FILLER_36_1720 ();
 FILLCELL_X32 FILLER_36_1752 ();
 FILLCELL_X32 FILLER_36_1784 ();
 FILLCELL_X32 FILLER_36_1816 ();
 FILLCELL_X32 FILLER_36_1848 ();
 FILLCELL_X8 FILLER_36_1880 ();
 FILLCELL_X4 FILLER_36_1888 ();
 FILLCELL_X2 FILLER_36_1892 ();
 FILLCELL_X32 FILLER_36_1895 ();
 FILLCELL_X32 FILLER_36_1927 ();
 FILLCELL_X32 FILLER_36_1959 ();
 FILLCELL_X32 FILLER_36_1991 ();
 FILLCELL_X32 FILLER_36_2023 ();
 FILLCELL_X32 FILLER_36_2055 ();
 FILLCELL_X16 FILLER_36_2087 ();
 FILLCELL_X8 FILLER_36_2103 ();
 FILLCELL_X4 FILLER_36_2111 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X32 FILLER_37_1584 ();
 FILLCELL_X32 FILLER_37_1616 ();
 FILLCELL_X32 FILLER_37_1648 ();
 FILLCELL_X32 FILLER_37_1680 ();
 FILLCELL_X32 FILLER_37_1712 ();
 FILLCELL_X32 FILLER_37_1744 ();
 FILLCELL_X32 FILLER_37_1776 ();
 FILLCELL_X32 FILLER_37_1808 ();
 FILLCELL_X32 FILLER_37_1840 ();
 FILLCELL_X32 FILLER_37_1872 ();
 FILLCELL_X32 FILLER_37_1904 ();
 FILLCELL_X32 FILLER_37_1936 ();
 FILLCELL_X32 FILLER_37_1968 ();
 FILLCELL_X32 FILLER_37_2000 ();
 FILLCELL_X32 FILLER_37_2032 ();
 FILLCELL_X32 FILLER_37_2064 ();
 FILLCELL_X16 FILLER_37_2096 ();
 FILLCELL_X2 FILLER_37_2112 ();
 FILLCELL_X1 FILLER_37_2114 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X32 FILLER_38_1592 ();
 FILLCELL_X32 FILLER_38_1624 ();
 FILLCELL_X32 FILLER_38_1656 ();
 FILLCELL_X32 FILLER_38_1688 ();
 FILLCELL_X32 FILLER_38_1720 ();
 FILLCELL_X32 FILLER_38_1752 ();
 FILLCELL_X32 FILLER_38_1784 ();
 FILLCELL_X32 FILLER_38_1816 ();
 FILLCELL_X32 FILLER_38_1848 ();
 FILLCELL_X8 FILLER_38_1880 ();
 FILLCELL_X4 FILLER_38_1888 ();
 FILLCELL_X2 FILLER_38_1892 ();
 FILLCELL_X32 FILLER_38_1895 ();
 FILLCELL_X32 FILLER_38_1927 ();
 FILLCELL_X32 FILLER_38_1959 ();
 FILLCELL_X32 FILLER_38_1991 ();
 FILLCELL_X32 FILLER_38_2023 ();
 FILLCELL_X32 FILLER_38_2055 ();
 FILLCELL_X16 FILLER_38_2087 ();
 FILLCELL_X8 FILLER_38_2103 ();
 FILLCELL_X4 FILLER_38_2111 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X32 FILLER_39_1584 ();
 FILLCELL_X32 FILLER_39_1616 ();
 FILLCELL_X32 FILLER_39_1648 ();
 FILLCELL_X32 FILLER_39_1680 ();
 FILLCELL_X32 FILLER_39_1712 ();
 FILLCELL_X32 FILLER_39_1744 ();
 FILLCELL_X32 FILLER_39_1776 ();
 FILLCELL_X32 FILLER_39_1808 ();
 FILLCELL_X32 FILLER_39_1840 ();
 FILLCELL_X32 FILLER_39_1872 ();
 FILLCELL_X32 FILLER_39_1904 ();
 FILLCELL_X32 FILLER_39_1936 ();
 FILLCELL_X32 FILLER_39_1968 ();
 FILLCELL_X32 FILLER_39_2000 ();
 FILLCELL_X32 FILLER_39_2032 ();
 FILLCELL_X32 FILLER_39_2064 ();
 FILLCELL_X16 FILLER_39_2096 ();
 FILLCELL_X2 FILLER_39_2112 ();
 FILLCELL_X1 FILLER_39_2114 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X32 FILLER_40_1592 ();
 FILLCELL_X32 FILLER_40_1624 ();
 FILLCELL_X32 FILLER_40_1656 ();
 FILLCELL_X32 FILLER_40_1688 ();
 FILLCELL_X32 FILLER_40_1720 ();
 FILLCELL_X32 FILLER_40_1752 ();
 FILLCELL_X32 FILLER_40_1784 ();
 FILLCELL_X32 FILLER_40_1816 ();
 FILLCELL_X32 FILLER_40_1848 ();
 FILLCELL_X8 FILLER_40_1880 ();
 FILLCELL_X4 FILLER_40_1888 ();
 FILLCELL_X2 FILLER_40_1892 ();
 FILLCELL_X32 FILLER_40_1895 ();
 FILLCELL_X32 FILLER_40_1927 ();
 FILLCELL_X32 FILLER_40_1959 ();
 FILLCELL_X32 FILLER_40_1991 ();
 FILLCELL_X32 FILLER_40_2023 ();
 FILLCELL_X32 FILLER_40_2055 ();
 FILLCELL_X16 FILLER_40_2087 ();
 FILLCELL_X8 FILLER_40_2103 ();
 FILLCELL_X4 FILLER_40_2111 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X32 FILLER_41_1584 ();
 FILLCELL_X32 FILLER_41_1616 ();
 FILLCELL_X32 FILLER_41_1648 ();
 FILLCELL_X32 FILLER_41_1680 ();
 FILLCELL_X32 FILLER_41_1712 ();
 FILLCELL_X32 FILLER_41_1744 ();
 FILLCELL_X32 FILLER_41_1776 ();
 FILLCELL_X32 FILLER_41_1808 ();
 FILLCELL_X32 FILLER_41_1840 ();
 FILLCELL_X32 FILLER_41_1872 ();
 FILLCELL_X32 FILLER_41_1904 ();
 FILLCELL_X32 FILLER_41_1936 ();
 FILLCELL_X32 FILLER_41_1968 ();
 FILLCELL_X32 FILLER_41_2000 ();
 FILLCELL_X32 FILLER_41_2032 ();
 FILLCELL_X32 FILLER_41_2064 ();
 FILLCELL_X16 FILLER_41_2096 ();
 FILLCELL_X2 FILLER_41_2112 ();
 FILLCELL_X1 FILLER_41_2114 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X32 FILLER_42_1592 ();
 FILLCELL_X32 FILLER_42_1624 ();
 FILLCELL_X32 FILLER_42_1656 ();
 FILLCELL_X32 FILLER_42_1688 ();
 FILLCELL_X32 FILLER_42_1720 ();
 FILLCELL_X32 FILLER_42_1752 ();
 FILLCELL_X32 FILLER_42_1784 ();
 FILLCELL_X32 FILLER_42_1816 ();
 FILLCELL_X32 FILLER_42_1848 ();
 FILLCELL_X8 FILLER_42_1880 ();
 FILLCELL_X4 FILLER_42_1888 ();
 FILLCELL_X2 FILLER_42_1892 ();
 FILLCELL_X32 FILLER_42_1895 ();
 FILLCELL_X32 FILLER_42_1927 ();
 FILLCELL_X32 FILLER_42_1959 ();
 FILLCELL_X32 FILLER_42_1991 ();
 FILLCELL_X32 FILLER_42_2023 ();
 FILLCELL_X32 FILLER_42_2055 ();
 FILLCELL_X16 FILLER_42_2087 ();
 FILLCELL_X8 FILLER_42_2103 ();
 FILLCELL_X4 FILLER_42_2111 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X32 FILLER_43_1584 ();
 FILLCELL_X32 FILLER_43_1616 ();
 FILLCELL_X32 FILLER_43_1648 ();
 FILLCELL_X32 FILLER_43_1680 ();
 FILLCELL_X32 FILLER_43_1712 ();
 FILLCELL_X32 FILLER_43_1744 ();
 FILLCELL_X32 FILLER_43_1776 ();
 FILLCELL_X32 FILLER_43_1808 ();
 FILLCELL_X32 FILLER_43_1840 ();
 FILLCELL_X32 FILLER_43_1872 ();
 FILLCELL_X32 FILLER_43_1904 ();
 FILLCELL_X32 FILLER_43_1936 ();
 FILLCELL_X32 FILLER_43_1968 ();
 FILLCELL_X32 FILLER_43_2000 ();
 FILLCELL_X32 FILLER_43_2032 ();
 FILLCELL_X32 FILLER_43_2064 ();
 FILLCELL_X16 FILLER_43_2096 ();
 FILLCELL_X2 FILLER_43_2112 ();
 FILLCELL_X1 FILLER_43_2114 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X32 FILLER_44_1592 ();
 FILLCELL_X32 FILLER_44_1624 ();
 FILLCELL_X32 FILLER_44_1656 ();
 FILLCELL_X32 FILLER_44_1688 ();
 FILLCELL_X32 FILLER_44_1720 ();
 FILLCELL_X32 FILLER_44_1752 ();
 FILLCELL_X32 FILLER_44_1784 ();
 FILLCELL_X32 FILLER_44_1816 ();
 FILLCELL_X32 FILLER_44_1848 ();
 FILLCELL_X8 FILLER_44_1880 ();
 FILLCELL_X4 FILLER_44_1888 ();
 FILLCELL_X2 FILLER_44_1892 ();
 FILLCELL_X32 FILLER_44_1895 ();
 FILLCELL_X32 FILLER_44_1927 ();
 FILLCELL_X32 FILLER_44_1959 ();
 FILLCELL_X32 FILLER_44_1991 ();
 FILLCELL_X32 FILLER_44_2023 ();
 FILLCELL_X32 FILLER_44_2055 ();
 FILLCELL_X16 FILLER_44_2087 ();
 FILLCELL_X8 FILLER_44_2103 ();
 FILLCELL_X4 FILLER_44_2111 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X32 FILLER_45_1584 ();
 FILLCELL_X32 FILLER_45_1616 ();
 FILLCELL_X32 FILLER_45_1648 ();
 FILLCELL_X32 FILLER_45_1680 ();
 FILLCELL_X32 FILLER_45_1712 ();
 FILLCELL_X32 FILLER_45_1744 ();
 FILLCELL_X32 FILLER_45_1776 ();
 FILLCELL_X32 FILLER_45_1808 ();
 FILLCELL_X32 FILLER_45_1840 ();
 FILLCELL_X32 FILLER_45_1872 ();
 FILLCELL_X32 FILLER_45_1904 ();
 FILLCELL_X32 FILLER_45_1936 ();
 FILLCELL_X32 FILLER_45_1968 ();
 FILLCELL_X32 FILLER_45_2000 ();
 FILLCELL_X32 FILLER_45_2032 ();
 FILLCELL_X32 FILLER_45_2064 ();
 FILLCELL_X16 FILLER_45_2096 ();
 FILLCELL_X2 FILLER_45_2112 ();
 FILLCELL_X1 FILLER_45_2114 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X32 FILLER_46_1592 ();
 FILLCELL_X32 FILLER_46_1624 ();
 FILLCELL_X32 FILLER_46_1656 ();
 FILLCELL_X32 FILLER_46_1688 ();
 FILLCELL_X32 FILLER_46_1720 ();
 FILLCELL_X32 FILLER_46_1752 ();
 FILLCELL_X32 FILLER_46_1784 ();
 FILLCELL_X32 FILLER_46_1816 ();
 FILLCELL_X32 FILLER_46_1848 ();
 FILLCELL_X8 FILLER_46_1880 ();
 FILLCELL_X4 FILLER_46_1888 ();
 FILLCELL_X2 FILLER_46_1892 ();
 FILLCELL_X32 FILLER_46_1895 ();
 FILLCELL_X32 FILLER_46_1927 ();
 FILLCELL_X32 FILLER_46_1959 ();
 FILLCELL_X32 FILLER_46_1991 ();
 FILLCELL_X32 FILLER_46_2023 ();
 FILLCELL_X32 FILLER_46_2055 ();
 FILLCELL_X16 FILLER_46_2087 ();
 FILLCELL_X8 FILLER_46_2103 ();
 FILLCELL_X4 FILLER_46_2111 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X32 FILLER_47_1584 ();
 FILLCELL_X32 FILLER_47_1616 ();
 FILLCELL_X32 FILLER_47_1648 ();
 FILLCELL_X32 FILLER_47_1680 ();
 FILLCELL_X32 FILLER_47_1712 ();
 FILLCELL_X32 FILLER_47_1744 ();
 FILLCELL_X32 FILLER_47_1776 ();
 FILLCELL_X32 FILLER_47_1808 ();
 FILLCELL_X32 FILLER_47_1840 ();
 FILLCELL_X32 FILLER_47_1872 ();
 FILLCELL_X32 FILLER_47_1904 ();
 FILLCELL_X32 FILLER_47_1936 ();
 FILLCELL_X32 FILLER_47_1968 ();
 FILLCELL_X32 FILLER_47_2000 ();
 FILLCELL_X32 FILLER_47_2032 ();
 FILLCELL_X32 FILLER_47_2064 ();
 FILLCELL_X16 FILLER_47_2096 ();
 FILLCELL_X2 FILLER_47_2112 ();
 FILLCELL_X1 FILLER_47_2114 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X32 FILLER_48_1592 ();
 FILLCELL_X32 FILLER_48_1624 ();
 FILLCELL_X32 FILLER_48_1656 ();
 FILLCELL_X32 FILLER_48_1688 ();
 FILLCELL_X32 FILLER_48_1720 ();
 FILLCELL_X32 FILLER_48_1752 ();
 FILLCELL_X32 FILLER_48_1784 ();
 FILLCELL_X32 FILLER_48_1816 ();
 FILLCELL_X32 FILLER_48_1848 ();
 FILLCELL_X8 FILLER_48_1880 ();
 FILLCELL_X4 FILLER_48_1888 ();
 FILLCELL_X2 FILLER_48_1892 ();
 FILLCELL_X32 FILLER_48_1895 ();
 FILLCELL_X32 FILLER_48_1927 ();
 FILLCELL_X32 FILLER_48_1959 ();
 FILLCELL_X32 FILLER_48_1991 ();
 FILLCELL_X32 FILLER_48_2023 ();
 FILLCELL_X32 FILLER_48_2055 ();
 FILLCELL_X16 FILLER_48_2087 ();
 FILLCELL_X8 FILLER_48_2103 ();
 FILLCELL_X4 FILLER_48_2111 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X32 FILLER_49_1584 ();
 FILLCELL_X32 FILLER_49_1616 ();
 FILLCELL_X32 FILLER_49_1648 ();
 FILLCELL_X32 FILLER_49_1680 ();
 FILLCELL_X32 FILLER_49_1712 ();
 FILLCELL_X32 FILLER_49_1744 ();
 FILLCELL_X32 FILLER_49_1776 ();
 FILLCELL_X32 FILLER_49_1808 ();
 FILLCELL_X32 FILLER_49_1840 ();
 FILLCELL_X32 FILLER_49_1872 ();
 FILLCELL_X32 FILLER_49_1904 ();
 FILLCELL_X32 FILLER_49_1936 ();
 FILLCELL_X32 FILLER_49_1968 ();
 FILLCELL_X32 FILLER_49_2000 ();
 FILLCELL_X32 FILLER_49_2032 ();
 FILLCELL_X32 FILLER_49_2064 ();
 FILLCELL_X16 FILLER_49_2096 ();
 FILLCELL_X2 FILLER_49_2112 ();
 FILLCELL_X1 FILLER_49_2114 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X32 FILLER_50_1592 ();
 FILLCELL_X32 FILLER_50_1624 ();
 FILLCELL_X32 FILLER_50_1656 ();
 FILLCELL_X32 FILLER_50_1688 ();
 FILLCELL_X32 FILLER_50_1720 ();
 FILLCELL_X32 FILLER_50_1752 ();
 FILLCELL_X32 FILLER_50_1784 ();
 FILLCELL_X32 FILLER_50_1816 ();
 FILLCELL_X32 FILLER_50_1848 ();
 FILLCELL_X8 FILLER_50_1880 ();
 FILLCELL_X4 FILLER_50_1888 ();
 FILLCELL_X2 FILLER_50_1892 ();
 FILLCELL_X32 FILLER_50_1895 ();
 FILLCELL_X32 FILLER_50_1927 ();
 FILLCELL_X32 FILLER_50_1959 ();
 FILLCELL_X32 FILLER_50_1991 ();
 FILLCELL_X32 FILLER_50_2023 ();
 FILLCELL_X32 FILLER_50_2055 ();
 FILLCELL_X16 FILLER_50_2087 ();
 FILLCELL_X8 FILLER_50_2103 ();
 FILLCELL_X4 FILLER_50_2111 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X32 FILLER_51_1584 ();
 FILLCELL_X32 FILLER_51_1616 ();
 FILLCELL_X32 FILLER_51_1648 ();
 FILLCELL_X32 FILLER_51_1680 ();
 FILLCELL_X32 FILLER_51_1712 ();
 FILLCELL_X32 FILLER_51_1744 ();
 FILLCELL_X32 FILLER_51_1776 ();
 FILLCELL_X32 FILLER_51_1808 ();
 FILLCELL_X32 FILLER_51_1840 ();
 FILLCELL_X32 FILLER_51_1872 ();
 FILLCELL_X32 FILLER_51_1904 ();
 FILLCELL_X32 FILLER_51_1936 ();
 FILLCELL_X32 FILLER_51_1968 ();
 FILLCELL_X32 FILLER_51_2000 ();
 FILLCELL_X32 FILLER_51_2032 ();
 FILLCELL_X32 FILLER_51_2064 ();
 FILLCELL_X16 FILLER_51_2096 ();
 FILLCELL_X2 FILLER_51_2112 ();
 FILLCELL_X1 FILLER_51_2114 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X32 FILLER_52_1592 ();
 FILLCELL_X32 FILLER_52_1624 ();
 FILLCELL_X32 FILLER_52_1656 ();
 FILLCELL_X32 FILLER_52_1688 ();
 FILLCELL_X32 FILLER_52_1720 ();
 FILLCELL_X32 FILLER_52_1752 ();
 FILLCELL_X32 FILLER_52_1784 ();
 FILLCELL_X32 FILLER_52_1816 ();
 FILLCELL_X32 FILLER_52_1848 ();
 FILLCELL_X8 FILLER_52_1880 ();
 FILLCELL_X4 FILLER_52_1888 ();
 FILLCELL_X2 FILLER_52_1892 ();
 FILLCELL_X32 FILLER_52_1895 ();
 FILLCELL_X32 FILLER_52_1927 ();
 FILLCELL_X32 FILLER_52_1959 ();
 FILLCELL_X32 FILLER_52_1991 ();
 FILLCELL_X32 FILLER_52_2023 ();
 FILLCELL_X32 FILLER_52_2055 ();
 FILLCELL_X16 FILLER_52_2087 ();
 FILLCELL_X8 FILLER_52_2103 ();
 FILLCELL_X4 FILLER_52_2111 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X32 FILLER_53_1584 ();
 FILLCELL_X32 FILLER_53_1616 ();
 FILLCELL_X32 FILLER_53_1648 ();
 FILLCELL_X32 FILLER_53_1680 ();
 FILLCELL_X32 FILLER_53_1712 ();
 FILLCELL_X32 FILLER_53_1744 ();
 FILLCELL_X32 FILLER_53_1776 ();
 FILLCELL_X32 FILLER_53_1808 ();
 FILLCELL_X32 FILLER_53_1840 ();
 FILLCELL_X32 FILLER_53_1872 ();
 FILLCELL_X32 FILLER_53_1904 ();
 FILLCELL_X32 FILLER_53_1936 ();
 FILLCELL_X32 FILLER_53_1968 ();
 FILLCELL_X32 FILLER_53_2000 ();
 FILLCELL_X32 FILLER_53_2032 ();
 FILLCELL_X32 FILLER_53_2064 ();
 FILLCELL_X16 FILLER_53_2096 ();
 FILLCELL_X2 FILLER_53_2112 ();
 FILLCELL_X1 FILLER_53_2114 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X32 FILLER_54_1592 ();
 FILLCELL_X32 FILLER_54_1624 ();
 FILLCELL_X32 FILLER_54_1656 ();
 FILLCELL_X32 FILLER_54_1688 ();
 FILLCELL_X32 FILLER_54_1720 ();
 FILLCELL_X32 FILLER_54_1752 ();
 FILLCELL_X32 FILLER_54_1784 ();
 FILLCELL_X32 FILLER_54_1816 ();
 FILLCELL_X32 FILLER_54_1848 ();
 FILLCELL_X8 FILLER_54_1880 ();
 FILLCELL_X4 FILLER_54_1888 ();
 FILLCELL_X2 FILLER_54_1892 ();
 FILLCELL_X32 FILLER_54_1895 ();
 FILLCELL_X32 FILLER_54_1927 ();
 FILLCELL_X32 FILLER_54_1959 ();
 FILLCELL_X32 FILLER_54_1991 ();
 FILLCELL_X32 FILLER_54_2023 ();
 FILLCELL_X32 FILLER_54_2055 ();
 FILLCELL_X16 FILLER_54_2087 ();
 FILLCELL_X8 FILLER_54_2103 ();
 FILLCELL_X4 FILLER_54_2111 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X32 FILLER_55_1584 ();
 FILLCELL_X32 FILLER_55_1616 ();
 FILLCELL_X32 FILLER_55_1648 ();
 FILLCELL_X32 FILLER_55_1680 ();
 FILLCELL_X32 FILLER_55_1712 ();
 FILLCELL_X32 FILLER_55_1744 ();
 FILLCELL_X32 FILLER_55_1776 ();
 FILLCELL_X32 FILLER_55_1808 ();
 FILLCELL_X32 FILLER_55_1840 ();
 FILLCELL_X32 FILLER_55_1872 ();
 FILLCELL_X32 FILLER_55_1904 ();
 FILLCELL_X32 FILLER_55_1936 ();
 FILLCELL_X32 FILLER_55_1968 ();
 FILLCELL_X32 FILLER_55_2000 ();
 FILLCELL_X32 FILLER_55_2032 ();
 FILLCELL_X32 FILLER_55_2064 ();
 FILLCELL_X16 FILLER_55_2096 ();
 FILLCELL_X2 FILLER_55_2112 ();
 FILLCELL_X1 FILLER_55_2114 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X32 FILLER_56_1592 ();
 FILLCELL_X32 FILLER_56_1624 ();
 FILLCELL_X32 FILLER_56_1656 ();
 FILLCELL_X32 FILLER_56_1688 ();
 FILLCELL_X32 FILLER_56_1720 ();
 FILLCELL_X32 FILLER_56_1752 ();
 FILLCELL_X32 FILLER_56_1784 ();
 FILLCELL_X32 FILLER_56_1816 ();
 FILLCELL_X32 FILLER_56_1848 ();
 FILLCELL_X8 FILLER_56_1880 ();
 FILLCELL_X4 FILLER_56_1888 ();
 FILLCELL_X2 FILLER_56_1892 ();
 FILLCELL_X32 FILLER_56_1895 ();
 FILLCELL_X32 FILLER_56_1927 ();
 FILLCELL_X32 FILLER_56_1959 ();
 FILLCELL_X32 FILLER_56_1991 ();
 FILLCELL_X32 FILLER_56_2023 ();
 FILLCELL_X32 FILLER_56_2055 ();
 FILLCELL_X16 FILLER_56_2087 ();
 FILLCELL_X8 FILLER_56_2103 ();
 FILLCELL_X4 FILLER_56_2111 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X32 FILLER_57_1584 ();
 FILLCELL_X32 FILLER_57_1616 ();
 FILLCELL_X32 FILLER_57_1648 ();
 FILLCELL_X32 FILLER_57_1680 ();
 FILLCELL_X32 FILLER_57_1712 ();
 FILLCELL_X32 FILLER_57_1744 ();
 FILLCELL_X32 FILLER_57_1776 ();
 FILLCELL_X32 FILLER_57_1808 ();
 FILLCELL_X32 FILLER_57_1840 ();
 FILLCELL_X32 FILLER_57_1872 ();
 FILLCELL_X32 FILLER_57_1904 ();
 FILLCELL_X32 FILLER_57_1936 ();
 FILLCELL_X32 FILLER_57_1968 ();
 FILLCELL_X32 FILLER_57_2000 ();
 FILLCELL_X32 FILLER_57_2032 ();
 FILLCELL_X32 FILLER_57_2064 ();
 FILLCELL_X16 FILLER_57_2096 ();
 FILLCELL_X2 FILLER_57_2112 ();
 FILLCELL_X1 FILLER_57_2114 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X32 FILLER_58_1592 ();
 FILLCELL_X32 FILLER_58_1624 ();
 FILLCELL_X32 FILLER_58_1656 ();
 FILLCELL_X32 FILLER_58_1688 ();
 FILLCELL_X32 FILLER_58_1720 ();
 FILLCELL_X32 FILLER_58_1752 ();
 FILLCELL_X32 FILLER_58_1784 ();
 FILLCELL_X32 FILLER_58_1816 ();
 FILLCELL_X32 FILLER_58_1848 ();
 FILLCELL_X8 FILLER_58_1880 ();
 FILLCELL_X4 FILLER_58_1888 ();
 FILLCELL_X2 FILLER_58_1892 ();
 FILLCELL_X32 FILLER_58_1895 ();
 FILLCELL_X32 FILLER_58_1927 ();
 FILLCELL_X32 FILLER_58_1959 ();
 FILLCELL_X32 FILLER_58_1991 ();
 FILLCELL_X32 FILLER_58_2023 ();
 FILLCELL_X32 FILLER_58_2055 ();
 FILLCELL_X16 FILLER_58_2087 ();
 FILLCELL_X8 FILLER_58_2103 ();
 FILLCELL_X4 FILLER_58_2111 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X32 FILLER_59_1584 ();
 FILLCELL_X32 FILLER_59_1616 ();
 FILLCELL_X32 FILLER_59_1648 ();
 FILLCELL_X32 FILLER_59_1680 ();
 FILLCELL_X32 FILLER_59_1712 ();
 FILLCELL_X32 FILLER_59_1744 ();
 FILLCELL_X32 FILLER_59_1776 ();
 FILLCELL_X32 FILLER_59_1808 ();
 FILLCELL_X32 FILLER_59_1840 ();
 FILLCELL_X32 FILLER_59_1872 ();
 FILLCELL_X32 FILLER_59_1904 ();
 FILLCELL_X32 FILLER_59_1936 ();
 FILLCELL_X32 FILLER_59_1968 ();
 FILLCELL_X32 FILLER_59_2000 ();
 FILLCELL_X32 FILLER_59_2032 ();
 FILLCELL_X32 FILLER_59_2064 ();
 FILLCELL_X16 FILLER_59_2096 ();
 FILLCELL_X2 FILLER_59_2112 ();
 FILLCELL_X1 FILLER_59_2114 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X32 FILLER_60_1592 ();
 FILLCELL_X32 FILLER_60_1624 ();
 FILLCELL_X32 FILLER_60_1656 ();
 FILLCELL_X32 FILLER_60_1688 ();
 FILLCELL_X32 FILLER_60_1720 ();
 FILLCELL_X32 FILLER_60_1752 ();
 FILLCELL_X32 FILLER_60_1784 ();
 FILLCELL_X32 FILLER_60_1816 ();
 FILLCELL_X32 FILLER_60_1848 ();
 FILLCELL_X8 FILLER_60_1880 ();
 FILLCELL_X4 FILLER_60_1888 ();
 FILLCELL_X2 FILLER_60_1892 ();
 FILLCELL_X32 FILLER_60_1895 ();
 FILLCELL_X32 FILLER_60_1927 ();
 FILLCELL_X32 FILLER_60_1959 ();
 FILLCELL_X32 FILLER_60_1991 ();
 FILLCELL_X32 FILLER_60_2023 ();
 FILLCELL_X32 FILLER_60_2055 ();
 FILLCELL_X16 FILLER_60_2087 ();
 FILLCELL_X8 FILLER_60_2103 ();
 FILLCELL_X4 FILLER_60_2111 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X32 FILLER_61_1584 ();
 FILLCELL_X32 FILLER_61_1616 ();
 FILLCELL_X32 FILLER_61_1648 ();
 FILLCELL_X32 FILLER_61_1680 ();
 FILLCELL_X32 FILLER_61_1712 ();
 FILLCELL_X32 FILLER_61_1744 ();
 FILLCELL_X32 FILLER_61_1776 ();
 FILLCELL_X32 FILLER_61_1808 ();
 FILLCELL_X32 FILLER_61_1840 ();
 FILLCELL_X32 FILLER_61_1872 ();
 FILLCELL_X32 FILLER_61_1904 ();
 FILLCELL_X32 FILLER_61_1936 ();
 FILLCELL_X32 FILLER_61_1968 ();
 FILLCELL_X32 FILLER_61_2000 ();
 FILLCELL_X32 FILLER_61_2032 ();
 FILLCELL_X32 FILLER_61_2064 ();
 FILLCELL_X16 FILLER_61_2096 ();
 FILLCELL_X2 FILLER_61_2112 ();
 FILLCELL_X1 FILLER_61_2114 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X32 FILLER_62_1592 ();
 FILLCELL_X32 FILLER_62_1624 ();
 FILLCELL_X32 FILLER_62_1656 ();
 FILLCELL_X32 FILLER_62_1688 ();
 FILLCELL_X32 FILLER_62_1720 ();
 FILLCELL_X32 FILLER_62_1752 ();
 FILLCELL_X32 FILLER_62_1784 ();
 FILLCELL_X32 FILLER_62_1816 ();
 FILLCELL_X32 FILLER_62_1848 ();
 FILLCELL_X8 FILLER_62_1880 ();
 FILLCELL_X4 FILLER_62_1888 ();
 FILLCELL_X2 FILLER_62_1892 ();
 FILLCELL_X32 FILLER_62_1895 ();
 FILLCELL_X32 FILLER_62_1927 ();
 FILLCELL_X32 FILLER_62_1959 ();
 FILLCELL_X32 FILLER_62_1991 ();
 FILLCELL_X32 FILLER_62_2023 ();
 FILLCELL_X32 FILLER_62_2055 ();
 FILLCELL_X16 FILLER_62_2087 ();
 FILLCELL_X8 FILLER_62_2103 ();
 FILLCELL_X4 FILLER_62_2111 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X32 FILLER_63_1584 ();
 FILLCELL_X32 FILLER_63_1616 ();
 FILLCELL_X32 FILLER_63_1648 ();
 FILLCELL_X32 FILLER_63_1680 ();
 FILLCELL_X32 FILLER_63_1712 ();
 FILLCELL_X32 FILLER_63_1744 ();
 FILLCELL_X32 FILLER_63_1776 ();
 FILLCELL_X32 FILLER_63_1808 ();
 FILLCELL_X32 FILLER_63_1840 ();
 FILLCELL_X32 FILLER_63_1872 ();
 FILLCELL_X32 FILLER_63_1904 ();
 FILLCELL_X32 FILLER_63_1936 ();
 FILLCELL_X32 FILLER_63_1968 ();
 FILLCELL_X32 FILLER_63_2000 ();
 FILLCELL_X32 FILLER_63_2032 ();
 FILLCELL_X32 FILLER_63_2064 ();
 FILLCELL_X16 FILLER_63_2096 ();
 FILLCELL_X2 FILLER_63_2112 ();
 FILLCELL_X1 FILLER_63_2114 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X32 FILLER_64_1592 ();
 FILLCELL_X32 FILLER_64_1624 ();
 FILLCELL_X32 FILLER_64_1656 ();
 FILLCELL_X32 FILLER_64_1688 ();
 FILLCELL_X32 FILLER_64_1720 ();
 FILLCELL_X32 FILLER_64_1752 ();
 FILLCELL_X32 FILLER_64_1784 ();
 FILLCELL_X32 FILLER_64_1816 ();
 FILLCELL_X32 FILLER_64_1848 ();
 FILLCELL_X8 FILLER_64_1880 ();
 FILLCELL_X4 FILLER_64_1888 ();
 FILLCELL_X2 FILLER_64_1892 ();
 FILLCELL_X32 FILLER_64_1895 ();
 FILLCELL_X32 FILLER_64_1927 ();
 FILLCELL_X32 FILLER_64_1959 ();
 FILLCELL_X32 FILLER_64_1991 ();
 FILLCELL_X32 FILLER_64_2023 ();
 FILLCELL_X32 FILLER_64_2055 ();
 FILLCELL_X16 FILLER_64_2087 ();
 FILLCELL_X8 FILLER_64_2103 ();
 FILLCELL_X4 FILLER_64_2111 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X32 FILLER_65_1584 ();
 FILLCELL_X32 FILLER_65_1616 ();
 FILLCELL_X32 FILLER_65_1648 ();
 FILLCELL_X32 FILLER_65_1680 ();
 FILLCELL_X32 FILLER_65_1712 ();
 FILLCELL_X32 FILLER_65_1744 ();
 FILLCELL_X32 FILLER_65_1776 ();
 FILLCELL_X32 FILLER_65_1808 ();
 FILLCELL_X32 FILLER_65_1840 ();
 FILLCELL_X32 FILLER_65_1872 ();
 FILLCELL_X32 FILLER_65_1904 ();
 FILLCELL_X32 FILLER_65_1936 ();
 FILLCELL_X32 FILLER_65_1968 ();
 FILLCELL_X32 FILLER_65_2000 ();
 FILLCELL_X32 FILLER_65_2032 ();
 FILLCELL_X32 FILLER_65_2064 ();
 FILLCELL_X16 FILLER_65_2096 ();
 FILLCELL_X2 FILLER_65_2112 ();
 FILLCELL_X1 FILLER_65_2114 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X32 FILLER_66_1592 ();
 FILLCELL_X32 FILLER_66_1624 ();
 FILLCELL_X32 FILLER_66_1656 ();
 FILLCELL_X32 FILLER_66_1688 ();
 FILLCELL_X32 FILLER_66_1720 ();
 FILLCELL_X32 FILLER_66_1752 ();
 FILLCELL_X32 FILLER_66_1784 ();
 FILLCELL_X32 FILLER_66_1816 ();
 FILLCELL_X32 FILLER_66_1848 ();
 FILLCELL_X8 FILLER_66_1880 ();
 FILLCELL_X4 FILLER_66_1888 ();
 FILLCELL_X2 FILLER_66_1892 ();
 FILLCELL_X32 FILLER_66_1895 ();
 FILLCELL_X32 FILLER_66_1927 ();
 FILLCELL_X32 FILLER_66_1959 ();
 FILLCELL_X32 FILLER_66_1991 ();
 FILLCELL_X32 FILLER_66_2023 ();
 FILLCELL_X32 FILLER_66_2055 ();
 FILLCELL_X16 FILLER_66_2087 ();
 FILLCELL_X8 FILLER_66_2103 ();
 FILLCELL_X4 FILLER_66_2111 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X32 FILLER_67_801 ();
 FILLCELL_X32 FILLER_67_833 ();
 FILLCELL_X32 FILLER_67_865 ();
 FILLCELL_X32 FILLER_67_897 ();
 FILLCELL_X32 FILLER_67_929 ();
 FILLCELL_X32 FILLER_67_961 ();
 FILLCELL_X32 FILLER_67_993 ();
 FILLCELL_X32 FILLER_67_1025 ();
 FILLCELL_X32 FILLER_67_1057 ();
 FILLCELL_X32 FILLER_67_1089 ();
 FILLCELL_X32 FILLER_67_1121 ();
 FILLCELL_X32 FILLER_67_1153 ();
 FILLCELL_X32 FILLER_67_1185 ();
 FILLCELL_X32 FILLER_67_1217 ();
 FILLCELL_X8 FILLER_67_1249 ();
 FILLCELL_X4 FILLER_67_1257 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X32 FILLER_67_1584 ();
 FILLCELL_X32 FILLER_67_1616 ();
 FILLCELL_X32 FILLER_67_1648 ();
 FILLCELL_X32 FILLER_67_1680 ();
 FILLCELL_X32 FILLER_67_1712 ();
 FILLCELL_X32 FILLER_67_1744 ();
 FILLCELL_X32 FILLER_67_1776 ();
 FILLCELL_X32 FILLER_67_1808 ();
 FILLCELL_X32 FILLER_67_1840 ();
 FILLCELL_X32 FILLER_67_1872 ();
 FILLCELL_X32 FILLER_67_1904 ();
 FILLCELL_X32 FILLER_67_1936 ();
 FILLCELL_X32 FILLER_67_1968 ();
 FILLCELL_X32 FILLER_67_2000 ();
 FILLCELL_X32 FILLER_67_2032 ();
 FILLCELL_X32 FILLER_67_2064 ();
 FILLCELL_X16 FILLER_67_2096 ();
 FILLCELL_X2 FILLER_67_2112 ();
 FILLCELL_X1 FILLER_67_2114 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X32 FILLER_68_952 ();
 FILLCELL_X32 FILLER_68_984 ();
 FILLCELL_X32 FILLER_68_1016 ();
 FILLCELL_X32 FILLER_68_1048 ();
 FILLCELL_X32 FILLER_68_1080 ();
 FILLCELL_X32 FILLER_68_1112 ();
 FILLCELL_X32 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_68_1176 ();
 FILLCELL_X32 FILLER_68_1208 ();
 FILLCELL_X32 FILLER_68_1240 ();
 FILLCELL_X32 FILLER_68_1272 ();
 FILLCELL_X32 FILLER_68_1304 ();
 FILLCELL_X32 FILLER_68_1336 ();
 FILLCELL_X32 FILLER_68_1368 ();
 FILLCELL_X32 FILLER_68_1400 ();
 FILLCELL_X32 FILLER_68_1432 ();
 FILLCELL_X32 FILLER_68_1464 ();
 FILLCELL_X32 FILLER_68_1496 ();
 FILLCELL_X32 FILLER_68_1528 ();
 FILLCELL_X32 FILLER_68_1560 ();
 FILLCELL_X32 FILLER_68_1592 ();
 FILLCELL_X32 FILLER_68_1624 ();
 FILLCELL_X32 FILLER_68_1656 ();
 FILLCELL_X32 FILLER_68_1688 ();
 FILLCELL_X32 FILLER_68_1720 ();
 FILLCELL_X32 FILLER_68_1752 ();
 FILLCELL_X32 FILLER_68_1784 ();
 FILLCELL_X32 FILLER_68_1816 ();
 FILLCELL_X32 FILLER_68_1848 ();
 FILLCELL_X8 FILLER_68_1880 ();
 FILLCELL_X4 FILLER_68_1888 ();
 FILLCELL_X2 FILLER_68_1892 ();
 FILLCELL_X32 FILLER_68_1895 ();
 FILLCELL_X32 FILLER_68_1927 ();
 FILLCELL_X32 FILLER_68_1959 ();
 FILLCELL_X32 FILLER_68_1991 ();
 FILLCELL_X32 FILLER_68_2023 ();
 FILLCELL_X32 FILLER_68_2055 ();
 FILLCELL_X16 FILLER_68_2087 ();
 FILLCELL_X8 FILLER_68_2103 ();
 FILLCELL_X4 FILLER_68_2111 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X32 FILLER_69_833 ();
 FILLCELL_X32 FILLER_69_865 ();
 FILLCELL_X32 FILLER_69_897 ();
 FILLCELL_X32 FILLER_69_929 ();
 FILLCELL_X32 FILLER_69_961 ();
 FILLCELL_X32 FILLER_69_993 ();
 FILLCELL_X32 FILLER_69_1025 ();
 FILLCELL_X32 FILLER_69_1057 ();
 FILLCELL_X32 FILLER_69_1089 ();
 FILLCELL_X32 FILLER_69_1121 ();
 FILLCELL_X32 FILLER_69_1153 ();
 FILLCELL_X32 FILLER_69_1185 ();
 FILLCELL_X32 FILLER_69_1217 ();
 FILLCELL_X8 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1257 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X32 FILLER_69_1584 ();
 FILLCELL_X32 FILLER_69_1616 ();
 FILLCELL_X32 FILLER_69_1648 ();
 FILLCELL_X32 FILLER_69_1680 ();
 FILLCELL_X32 FILLER_69_1712 ();
 FILLCELL_X32 FILLER_69_1744 ();
 FILLCELL_X32 FILLER_69_1776 ();
 FILLCELL_X32 FILLER_69_1808 ();
 FILLCELL_X32 FILLER_69_1840 ();
 FILLCELL_X32 FILLER_69_1872 ();
 FILLCELL_X32 FILLER_69_1904 ();
 FILLCELL_X32 FILLER_69_1936 ();
 FILLCELL_X32 FILLER_69_1968 ();
 FILLCELL_X32 FILLER_69_2000 ();
 FILLCELL_X32 FILLER_69_2032 ();
 FILLCELL_X32 FILLER_69_2064 ();
 FILLCELL_X16 FILLER_69_2096 ();
 FILLCELL_X2 FILLER_69_2112 ();
 FILLCELL_X1 FILLER_69_2114 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X32 FILLER_70_1592 ();
 FILLCELL_X32 FILLER_70_1624 ();
 FILLCELL_X32 FILLER_70_1656 ();
 FILLCELL_X32 FILLER_70_1688 ();
 FILLCELL_X32 FILLER_70_1720 ();
 FILLCELL_X32 FILLER_70_1752 ();
 FILLCELL_X32 FILLER_70_1784 ();
 FILLCELL_X32 FILLER_70_1816 ();
 FILLCELL_X32 FILLER_70_1848 ();
 FILLCELL_X8 FILLER_70_1880 ();
 FILLCELL_X4 FILLER_70_1888 ();
 FILLCELL_X2 FILLER_70_1892 ();
 FILLCELL_X32 FILLER_70_1895 ();
 FILLCELL_X32 FILLER_70_1927 ();
 FILLCELL_X32 FILLER_70_1959 ();
 FILLCELL_X32 FILLER_70_1991 ();
 FILLCELL_X32 FILLER_70_2023 ();
 FILLCELL_X32 FILLER_70_2055 ();
 FILLCELL_X16 FILLER_70_2087 ();
 FILLCELL_X8 FILLER_70_2103 ();
 FILLCELL_X4 FILLER_70_2111 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1584 ();
 FILLCELL_X32 FILLER_71_1616 ();
 FILLCELL_X32 FILLER_71_1648 ();
 FILLCELL_X32 FILLER_71_1680 ();
 FILLCELL_X32 FILLER_71_1712 ();
 FILLCELL_X32 FILLER_71_1744 ();
 FILLCELL_X32 FILLER_71_1776 ();
 FILLCELL_X32 FILLER_71_1808 ();
 FILLCELL_X32 FILLER_71_1840 ();
 FILLCELL_X32 FILLER_71_1872 ();
 FILLCELL_X32 FILLER_71_1904 ();
 FILLCELL_X32 FILLER_71_1936 ();
 FILLCELL_X32 FILLER_71_1968 ();
 FILLCELL_X32 FILLER_71_2000 ();
 FILLCELL_X32 FILLER_71_2032 ();
 FILLCELL_X32 FILLER_71_2064 ();
 FILLCELL_X16 FILLER_71_2096 ();
 FILLCELL_X2 FILLER_71_2112 ();
 FILLCELL_X1 FILLER_71_2114 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X32 FILLER_72_1592 ();
 FILLCELL_X32 FILLER_72_1624 ();
 FILLCELL_X32 FILLER_72_1656 ();
 FILLCELL_X32 FILLER_72_1688 ();
 FILLCELL_X32 FILLER_72_1720 ();
 FILLCELL_X32 FILLER_72_1752 ();
 FILLCELL_X32 FILLER_72_1784 ();
 FILLCELL_X32 FILLER_72_1816 ();
 FILLCELL_X32 FILLER_72_1848 ();
 FILLCELL_X8 FILLER_72_1880 ();
 FILLCELL_X4 FILLER_72_1888 ();
 FILLCELL_X2 FILLER_72_1892 ();
 FILLCELL_X32 FILLER_72_1895 ();
 FILLCELL_X32 FILLER_72_1927 ();
 FILLCELL_X32 FILLER_72_1959 ();
 FILLCELL_X32 FILLER_72_1991 ();
 FILLCELL_X32 FILLER_72_2023 ();
 FILLCELL_X32 FILLER_72_2055 ();
 FILLCELL_X16 FILLER_72_2087 ();
 FILLCELL_X8 FILLER_72_2103 ();
 FILLCELL_X4 FILLER_72_2111 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X32 FILLER_73_1584 ();
 FILLCELL_X32 FILLER_73_1616 ();
 FILLCELL_X32 FILLER_73_1648 ();
 FILLCELL_X32 FILLER_73_1680 ();
 FILLCELL_X32 FILLER_73_1712 ();
 FILLCELL_X32 FILLER_73_1744 ();
 FILLCELL_X32 FILLER_73_1776 ();
 FILLCELL_X32 FILLER_73_1808 ();
 FILLCELL_X32 FILLER_73_1840 ();
 FILLCELL_X32 FILLER_73_1872 ();
 FILLCELL_X32 FILLER_73_1904 ();
 FILLCELL_X32 FILLER_73_1936 ();
 FILLCELL_X32 FILLER_73_1968 ();
 FILLCELL_X32 FILLER_73_2000 ();
 FILLCELL_X32 FILLER_73_2032 ();
 FILLCELL_X32 FILLER_73_2064 ();
 FILLCELL_X16 FILLER_73_2096 ();
 FILLCELL_X2 FILLER_73_2112 ();
 FILLCELL_X1 FILLER_73_2114 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X32 FILLER_74_1592 ();
 FILLCELL_X32 FILLER_74_1624 ();
 FILLCELL_X32 FILLER_74_1656 ();
 FILLCELL_X32 FILLER_74_1688 ();
 FILLCELL_X32 FILLER_74_1720 ();
 FILLCELL_X32 FILLER_74_1752 ();
 FILLCELL_X32 FILLER_74_1784 ();
 FILLCELL_X32 FILLER_74_1816 ();
 FILLCELL_X32 FILLER_74_1848 ();
 FILLCELL_X8 FILLER_74_1880 ();
 FILLCELL_X4 FILLER_74_1888 ();
 FILLCELL_X2 FILLER_74_1892 ();
 FILLCELL_X32 FILLER_74_1895 ();
 FILLCELL_X32 FILLER_74_1927 ();
 FILLCELL_X32 FILLER_74_1959 ();
 FILLCELL_X32 FILLER_74_1991 ();
 FILLCELL_X32 FILLER_74_2023 ();
 FILLCELL_X32 FILLER_74_2055 ();
 FILLCELL_X16 FILLER_74_2087 ();
 FILLCELL_X8 FILLER_74_2103 ();
 FILLCELL_X4 FILLER_74_2111 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X32 FILLER_75_865 ();
 FILLCELL_X32 FILLER_75_897 ();
 FILLCELL_X32 FILLER_75_929 ();
 FILLCELL_X32 FILLER_75_961 ();
 FILLCELL_X32 FILLER_75_993 ();
 FILLCELL_X32 FILLER_75_1025 ();
 FILLCELL_X32 FILLER_75_1057 ();
 FILLCELL_X32 FILLER_75_1089 ();
 FILLCELL_X32 FILLER_75_1121 ();
 FILLCELL_X32 FILLER_75_1153 ();
 FILLCELL_X32 FILLER_75_1185 ();
 FILLCELL_X32 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1249 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X32 FILLER_75_1584 ();
 FILLCELL_X32 FILLER_75_1616 ();
 FILLCELL_X32 FILLER_75_1648 ();
 FILLCELL_X32 FILLER_75_1680 ();
 FILLCELL_X32 FILLER_75_1712 ();
 FILLCELL_X32 FILLER_75_1744 ();
 FILLCELL_X32 FILLER_75_1776 ();
 FILLCELL_X32 FILLER_75_1808 ();
 FILLCELL_X32 FILLER_75_1840 ();
 FILLCELL_X32 FILLER_75_1872 ();
 FILLCELL_X32 FILLER_75_1904 ();
 FILLCELL_X32 FILLER_75_1936 ();
 FILLCELL_X32 FILLER_75_1968 ();
 FILLCELL_X32 FILLER_75_2000 ();
 FILLCELL_X32 FILLER_75_2032 ();
 FILLCELL_X32 FILLER_75_2064 ();
 FILLCELL_X16 FILLER_75_2096 ();
 FILLCELL_X2 FILLER_75_2112 ();
 FILLCELL_X1 FILLER_75_2114 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X32 FILLER_76_952 ();
 FILLCELL_X32 FILLER_76_984 ();
 FILLCELL_X32 FILLER_76_1016 ();
 FILLCELL_X32 FILLER_76_1048 ();
 FILLCELL_X32 FILLER_76_1080 ();
 FILLCELL_X32 FILLER_76_1112 ();
 FILLCELL_X32 FILLER_76_1144 ();
 FILLCELL_X32 FILLER_76_1176 ();
 FILLCELL_X32 FILLER_76_1208 ();
 FILLCELL_X32 FILLER_76_1240 ();
 FILLCELL_X32 FILLER_76_1272 ();
 FILLCELL_X32 FILLER_76_1304 ();
 FILLCELL_X32 FILLER_76_1336 ();
 FILLCELL_X32 FILLER_76_1368 ();
 FILLCELL_X32 FILLER_76_1400 ();
 FILLCELL_X32 FILLER_76_1432 ();
 FILLCELL_X32 FILLER_76_1464 ();
 FILLCELL_X32 FILLER_76_1496 ();
 FILLCELL_X32 FILLER_76_1528 ();
 FILLCELL_X32 FILLER_76_1560 ();
 FILLCELL_X32 FILLER_76_1592 ();
 FILLCELL_X32 FILLER_76_1624 ();
 FILLCELL_X32 FILLER_76_1656 ();
 FILLCELL_X32 FILLER_76_1688 ();
 FILLCELL_X32 FILLER_76_1720 ();
 FILLCELL_X32 FILLER_76_1752 ();
 FILLCELL_X32 FILLER_76_1784 ();
 FILLCELL_X32 FILLER_76_1816 ();
 FILLCELL_X32 FILLER_76_1848 ();
 FILLCELL_X8 FILLER_76_1880 ();
 FILLCELL_X4 FILLER_76_1888 ();
 FILLCELL_X2 FILLER_76_1892 ();
 FILLCELL_X32 FILLER_76_1895 ();
 FILLCELL_X32 FILLER_76_1927 ();
 FILLCELL_X32 FILLER_76_1959 ();
 FILLCELL_X32 FILLER_76_1991 ();
 FILLCELL_X32 FILLER_76_2023 ();
 FILLCELL_X32 FILLER_76_2055 ();
 FILLCELL_X16 FILLER_76_2087 ();
 FILLCELL_X8 FILLER_76_2103 ();
 FILLCELL_X4 FILLER_76_2111 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_961 ();
 FILLCELL_X32 FILLER_77_993 ();
 FILLCELL_X32 FILLER_77_1025 ();
 FILLCELL_X32 FILLER_77_1057 ();
 FILLCELL_X32 FILLER_77_1089 ();
 FILLCELL_X32 FILLER_77_1121 ();
 FILLCELL_X32 FILLER_77_1153 ();
 FILLCELL_X32 FILLER_77_1185 ();
 FILLCELL_X32 FILLER_77_1217 ();
 FILLCELL_X8 FILLER_77_1249 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X32 FILLER_77_1584 ();
 FILLCELL_X32 FILLER_77_1616 ();
 FILLCELL_X32 FILLER_77_1648 ();
 FILLCELL_X32 FILLER_77_1680 ();
 FILLCELL_X32 FILLER_77_1712 ();
 FILLCELL_X32 FILLER_77_1744 ();
 FILLCELL_X32 FILLER_77_1776 ();
 FILLCELL_X32 FILLER_77_1808 ();
 FILLCELL_X32 FILLER_77_1840 ();
 FILLCELL_X32 FILLER_77_1872 ();
 FILLCELL_X32 FILLER_77_1904 ();
 FILLCELL_X32 FILLER_77_1936 ();
 FILLCELL_X32 FILLER_77_1968 ();
 FILLCELL_X32 FILLER_77_2000 ();
 FILLCELL_X32 FILLER_77_2032 ();
 FILLCELL_X32 FILLER_77_2064 ();
 FILLCELL_X16 FILLER_77_2096 ();
 FILLCELL_X2 FILLER_77_2112 ();
 FILLCELL_X1 FILLER_77_2114 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X32 FILLER_78_952 ();
 FILLCELL_X32 FILLER_78_984 ();
 FILLCELL_X32 FILLER_78_1016 ();
 FILLCELL_X32 FILLER_78_1048 ();
 FILLCELL_X32 FILLER_78_1080 ();
 FILLCELL_X32 FILLER_78_1112 ();
 FILLCELL_X32 FILLER_78_1144 ();
 FILLCELL_X32 FILLER_78_1176 ();
 FILLCELL_X32 FILLER_78_1208 ();
 FILLCELL_X32 FILLER_78_1240 ();
 FILLCELL_X32 FILLER_78_1272 ();
 FILLCELL_X32 FILLER_78_1304 ();
 FILLCELL_X32 FILLER_78_1336 ();
 FILLCELL_X32 FILLER_78_1368 ();
 FILLCELL_X32 FILLER_78_1400 ();
 FILLCELL_X32 FILLER_78_1432 ();
 FILLCELL_X32 FILLER_78_1464 ();
 FILLCELL_X32 FILLER_78_1496 ();
 FILLCELL_X32 FILLER_78_1528 ();
 FILLCELL_X32 FILLER_78_1560 ();
 FILLCELL_X32 FILLER_78_1592 ();
 FILLCELL_X32 FILLER_78_1624 ();
 FILLCELL_X32 FILLER_78_1656 ();
 FILLCELL_X32 FILLER_78_1688 ();
 FILLCELL_X32 FILLER_78_1720 ();
 FILLCELL_X32 FILLER_78_1752 ();
 FILLCELL_X32 FILLER_78_1784 ();
 FILLCELL_X32 FILLER_78_1816 ();
 FILLCELL_X32 FILLER_78_1848 ();
 FILLCELL_X8 FILLER_78_1880 ();
 FILLCELL_X4 FILLER_78_1888 ();
 FILLCELL_X2 FILLER_78_1892 ();
 FILLCELL_X32 FILLER_78_1895 ();
 FILLCELL_X32 FILLER_78_1927 ();
 FILLCELL_X32 FILLER_78_1959 ();
 FILLCELL_X32 FILLER_78_1991 ();
 FILLCELL_X32 FILLER_78_2023 ();
 FILLCELL_X32 FILLER_78_2055 ();
 FILLCELL_X16 FILLER_78_2087 ();
 FILLCELL_X8 FILLER_78_2103 ();
 FILLCELL_X4 FILLER_78_2111 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X32 FILLER_79_961 ();
 FILLCELL_X32 FILLER_79_993 ();
 FILLCELL_X32 FILLER_79_1025 ();
 FILLCELL_X32 FILLER_79_1057 ();
 FILLCELL_X32 FILLER_79_1089 ();
 FILLCELL_X32 FILLER_79_1121 ();
 FILLCELL_X32 FILLER_79_1153 ();
 FILLCELL_X32 FILLER_79_1185 ();
 FILLCELL_X32 FILLER_79_1217 ();
 FILLCELL_X8 FILLER_79_1249 ();
 FILLCELL_X4 FILLER_79_1257 ();
 FILLCELL_X2 FILLER_79_1261 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X32 FILLER_79_1584 ();
 FILLCELL_X32 FILLER_79_1616 ();
 FILLCELL_X32 FILLER_79_1648 ();
 FILLCELL_X32 FILLER_79_1680 ();
 FILLCELL_X32 FILLER_79_1712 ();
 FILLCELL_X32 FILLER_79_1744 ();
 FILLCELL_X32 FILLER_79_1776 ();
 FILLCELL_X32 FILLER_79_1808 ();
 FILLCELL_X32 FILLER_79_1840 ();
 FILLCELL_X32 FILLER_79_1872 ();
 FILLCELL_X32 FILLER_79_1904 ();
 FILLCELL_X32 FILLER_79_1936 ();
 FILLCELL_X32 FILLER_79_1968 ();
 FILLCELL_X32 FILLER_79_2000 ();
 FILLCELL_X32 FILLER_79_2032 ();
 FILLCELL_X32 FILLER_79_2064 ();
 FILLCELL_X16 FILLER_79_2096 ();
 FILLCELL_X2 FILLER_79_2112 ();
 FILLCELL_X1 FILLER_79_2114 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X32 FILLER_80_952 ();
 FILLCELL_X32 FILLER_80_984 ();
 FILLCELL_X32 FILLER_80_1016 ();
 FILLCELL_X32 FILLER_80_1048 ();
 FILLCELL_X32 FILLER_80_1080 ();
 FILLCELL_X32 FILLER_80_1112 ();
 FILLCELL_X32 FILLER_80_1144 ();
 FILLCELL_X32 FILLER_80_1176 ();
 FILLCELL_X32 FILLER_80_1208 ();
 FILLCELL_X32 FILLER_80_1240 ();
 FILLCELL_X32 FILLER_80_1272 ();
 FILLCELL_X32 FILLER_80_1304 ();
 FILLCELL_X32 FILLER_80_1336 ();
 FILLCELL_X32 FILLER_80_1368 ();
 FILLCELL_X32 FILLER_80_1400 ();
 FILLCELL_X32 FILLER_80_1432 ();
 FILLCELL_X32 FILLER_80_1464 ();
 FILLCELL_X32 FILLER_80_1496 ();
 FILLCELL_X32 FILLER_80_1528 ();
 FILLCELL_X32 FILLER_80_1560 ();
 FILLCELL_X32 FILLER_80_1592 ();
 FILLCELL_X32 FILLER_80_1624 ();
 FILLCELL_X32 FILLER_80_1656 ();
 FILLCELL_X32 FILLER_80_1688 ();
 FILLCELL_X32 FILLER_80_1720 ();
 FILLCELL_X32 FILLER_80_1752 ();
 FILLCELL_X32 FILLER_80_1784 ();
 FILLCELL_X32 FILLER_80_1816 ();
 FILLCELL_X32 FILLER_80_1848 ();
 FILLCELL_X8 FILLER_80_1880 ();
 FILLCELL_X4 FILLER_80_1888 ();
 FILLCELL_X2 FILLER_80_1892 ();
 FILLCELL_X32 FILLER_80_1895 ();
 FILLCELL_X32 FILLER_80_1927 ();
 FILLCELL_X32 FILLER_80_1959 ();
 FILLCELL_X32 FILLER_80_1991 ();
 FILLCELL_X32 FILLER_80_2023 ();
 FILLCELL_X32 FILLER_80_2055 ();
 FILLCELL_X16 FILLER_80_2087 ();
 FILLCELL_X8 FILLER_80_2103 ();
 FILLCELL_X4 FILLER_80_2111 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X32 FILLER_81_1584 ();
 FILLCELL_X32 FILLER_81_1616 ();
 FILLCELL_X32 FILLER_81_1648 ();
 FILLCELL_X32 FILLER_81_1680 ();
 FILLCELL_X32 FILLER_81_1712 ();
 FILLCELL_X32 FILLER_81_1744 ();
 FILLCELL_X32 FILLER_81_1776 ();
 FILLCELL_X32 FILLER_81_1808 ();
 FILLCELL_X32 FILLER_81_1840 ();
 FILLCELL_X32 FILLER_81_1872 ();
 FILLCELL_X32 FILLER_81_1904 ();
 FILLCELL_X32 FILLER_81_1936 ();
 FILLCELL_X32 FILLER_81_1968 ();
 FILLCELL_X32 FILLER_81_2000 ();
 FILLCELL_X32 FILLER_81_2032 ();
 FILLCELL_X32 FILLER_81_2064 ();
 FILLCELL_X16 FILLER_81_2096 ();
 FILLCELL_X2 FILLER_81_2112 ();
 FILLCELL_X1 FILLER_81_2114 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X32 FILLER_82_1592 ();
 FILLCELL_X32 FILLER_82_1624 ();
 FILLCELL_X32 FILLER_82_1656 ();
 FILLCELL_X32 FILLER_82_1688 ();
 FILLCELL_X32 FILLER_82_1720 ();
 FILLCELL_X32 FILLER_82_1752 ();
 FILLCELL_X32 FILLER_82_1784 ();
 FILLCELL_X32 FILLER_82_1816 ();
 FILLCELL_X32 FILLER_82_1848 ();
 FILLCELL_X8 FILLER_82_1880 ();
 FILLCELL_X4 FILLER_82_1888 ();
 FILLCELL_X2 FILLER_82_1892 ();
 FILLCELL_X32 FILLER_82_1895 ();
 FILLCELL_X32 FILLER_82_1927 ();
 FILLCELL_X32 FILLER_82_1959 ();
 FILLCELL_X32 FILLER_82_1991 ();
 FILLCELL_X32 FILLER_82_2023 ();
 FILLCELL_X32 FILLER_82_2055 ();
 FILLCELL_X16 FILLER_82_2087 ();
 FILLCELL_X8 FILLER_82_2103 ();
 FILLCELL_X4 FILLER_82_2111 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X32 FILLER_83_1584 ();
 FILLCELL_X32 FILLER_83_1616 ();
 FILLCELL_X32 FILLER_83_1648 ();
 FILLCELL_X32 FILLER_83_1680 ();
 FILLCELL_X32 FILLER_83_1712 ();
 FILLCELL_X32 FILLER_83_1744 ();
 FILLCELL_X32 FILLER_83_1776 ();
 FILLCELL_X32 FILLER_83_1808 ();
 FILLCELL_X32 FILLER_83_1840 ();
 FILLCELL_X32 FILLER_83_1872 ();
 FILLCELL_X32 FILLER_83_1904 ();
 FILLCELL_X32 FILLER_83_1936 ();
 FILLCELL_X32 FILLER_83_1968 ();
 FILLCELL_X32 FILLER_83_2000 ();
 FILLCELL_X32 FILLER_83_2032 ();
 FILLCELL_X32 FILLER_83_2064 ();
 FILLCELL_X16 FILLER_83_2096 ();
 FILLCELL_X2 FILLER_83_2112 ();
 FILLCELL_X1 FILLER_83_2114 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X32 FILLER_84_1592 ();
 FILLCELL_X32 FILLER_84_1624 ();
 FILLCELL_X32 FILLER_84_1656 ();
 FILLCELL_X32 FILLER_84_1688 ();
 FILLCELL_X32 FILLER_84_1720 ();
 FILLCELL_X32 FILLER_84_1752 ();
 FILLCELL_X32 FILLER_84_1784 ();
 FILLCELL_X32 FILLER_84_1816 ();
 FILLCELL_X32 FILLER_84_1848 ();
 FILLCELL_X8 FILLER_84_1880 ();
 FILLCELL_X4 FILLER_84_1888 ();
 FILLCELL_X2 FILLER_84_1892 ();
 FILLCELL_X32 FILLER_84_1895 ();
 FILLCELL_X32 FILLER_84_1927 ();
 FILLCELL_X32 FILLER_84_1959 ();
 FILLCELL_X32 FILLER_84_1991 ();
 FILLCELL_X32 FILLER_84_2023 ();
 FILLCELL_X32 FILLER_84_2055 ();
 FILLCELL_X16 FILLER_84_2087 ();
 FILLCELL_X8 FILLER_84_2103 ();
 FILLCELL_X4 FILLER_84_2111 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X32 FILLER_85_1584 ();
 FILLCELL_X32 FILLER_85_1616 ();
 FILLCELL_X32 FILLER_85_1648 ();
 FILLCELL_X32 FILLER_85_1680 ();
 FILLCELL_X32 FILLER_85_1712 ();
 FILLCELL_X32 FILLER_85_1744 ();
 FILLCELL_X32 FILLER_85_1776 ();
 FILLCELL_X32 FILLER_85_1808 ();
 FILLCELL_X32 FILLER_85_1840 ();
 FILLCELL_X32 FILLER_85_1872 ();
 FILLCELL_X32 FILLER_85_1904 ();
 FILLCELL_X32 FILLER_85_1936 ();
 FILLCELL_X32 FILLER_85_1968 ();
 FILLCELL_X32 FILLER_85_2000 ();
 FILLCELL_X32 FILLER_85_2032 ();
 FILLCELL_X32 FILLER_85_2064 ();
 FILLCELL_X16 FILLER_85_2096 ();
 FILLCELL_X2 FILLER_85_2112 ();
 FILLCELL_X1 FILLER_85_2114 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X32 FILLER_86_1592 ();
 FILLCELL_X32 FILLER_86_1624 ();
 FILLCELL_X32 FILLER_86_1656 ();
 FILLCELL_X32 FILLER_86_1688 ();
 FILLCELL_X32 FILLER_86_1720 ();
 FILLCELL_X32 FILLER_86_1752 ();
 FILLCELL_X32 FILLER_86_1784 ();
 FILLCELL_X32 FILLER_86_1816 ();
 FILLCELL_X32 FILLER_86_1848 ();
 FILLCELL_X8 FILLER_86_1880 ();
 FILLCELL_X4 FILLER_86_1888 ();
 FILLCELL_X2 FILLER_86_1892 ();
 FILLCELL_X32 FILLER_86_1895 ();
 FILLCELL_X32 FILLER_86_1927 ();
 FILLCELL_X32 FILLER_86_1959 ();
 FILLCELL_X32 FILLER_86_1991 ();
 FILLCELL_X32 FILLER_86_2023 ();
 FILLCELL_X32 FILLER_86_2055 ();
 FILLCELL_X16 FILLER_86_2087 ();
 FILLCELL_X8 FILLER_86_2103 ();
 FILLCELL_X4 FILLER_86_2111 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X32 FILLER_87_1584 ();
 FILLCELL_X32 FILLER_87_1616 ();
 FILLCELL_X32 FILLER_87_1648 ();
 FILLCELL_X32 FILLER_87_1680 ();
 FILLCELL_X32 FILLER_87_1712 ();
 FILLCELL_X32 FILLER_87_1744 ();
 FILLCELL_X32 FILLER_87_1776 ();
 FILLCELL_X32 FILLER_87_1808 ();
 FILLCELL_X32 FILLER_87_1840 ();
 FILLCELL_X32 FILLER_87_1872 ();
 FILLCELL_X32 FILLER_87_1904 ();
 FILLCELL_X32 FILLER_87_1936 ();
 FILLCELL_X32 FILLER_87_1968 ();
 FILLCELL_X32 FILLER_87_2000 ();
 FILLCELL_X32 FILLER_87_2032 ();
 FILLCELL_X32 FILLER_87_2064 ();
 FILLCELL_X16 FILLER_87_2096 ();
 FILLCELL_X2 FILLER_87_2112 ();
 FILLCELL_X1 FILLER_87_2114 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X32 FILLER_88_1592 ();
 FILLCELL_X32 FILLER_88_1624 ();
 FILLCELL_X32 FILLER_88_1656 ();
 FILLCELL_X32 FILLER_88_1688 ();
 FILLCELL_X32 FILLER_88_1720 ();
 FILLCELL_X32 FILLER_88_1752 ();
 FILLCELL_X32 FILLER_88_1784 ();
 FILLCELL_X32 FILLER_88_1816 ();
 FILLCELL_X32 FILLER_88_1848 ();
 FILLCELL_X8 FILLER_88_1880 ();
 FILLCELL_X4 FILLER_88_1888 ();
 FILLCELL_X2 FILLER_88_1892 ();
 FILLCELL_X32 FILLER_88_1895 ();
 FILLCELL_X32 FILLER_88_1927 ();
 FILLCELL_X32 FILLER_88_1959 ();
 FILLCELL_X32 FILLER_88_1991 ();
 FILLCELL_X32 FILLER_88_2023 ();
 FILLCELL_X32 FILLER_88_2055 ();
 FILLCELL_X16 FILLER_88_2087 ();
 FILLCELL_X8 FILLER_88_2103 ();
 FILLCELL_X4 FILLER_88_2111 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X32 FILLER_89_1584 ();
 FILLCELL_X32 FILLER_89_1616 ();
 FILLCELL_X32 FILLER_89_1648 ();
 FILLCELL_X32 FILLER_89_1680 ();
 FILLCELL_X32 FILLER_89_1712 ();
 FILLCELL_X32 FILLER_89_1744 ();
 FILLCELL_X32 FILLER_89_1776 ();
 FILLCELL_X32 FILLER_89_1808 ();
 FILLCELL_X32 FILLER_89_1840 ();
 FILLCELL_X32 FILLER_89_1872 ();
 FILLCELL_X32 FILLER_89_1904 ();
 FILLCELL_X32 FILLER_89_1936 ();
 FILLCELL_X32 FILLER_89_1968 ();
 FILLCELL_X32 FILLER_89_2000 ();
 FILLCELL_X32 FILLER_89_2032 ();
 FILLCELL_X32 FILLER_89_2064 ();
 FILLCELL_X16 FILLER_89_2096 ();
 FILLCELL_X2 FILLER_89_2112 ();
 FILLCELL_X1 FILLER_89_2114 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X32 FILLER_90_1592 ();
 FILLCELL_X32 FILLER_90_1624 ();
 FILLCELL_X32 FILLER_90_1656 ();
 FILLCELL_X32 FILLER_90_1688 ();
 FILLCELL_X32 FILLER_90_1720 ();
 FILLCELL_X32 FILLER_90_1752 ();
 FILLCELL_X32 FILLER_90_1784 ();
 FILLCELL_X32 FILLER_90_1816 ();
 FILLCELL_X32 FILLER_90_1848 ();
 FILLCELL_X8 FILLER_90_1880 ();
 FILLCELL_X4 FILLER_90_1888 ();
 FILLCELL_X2 FILLER_90_1892 ();
 FILLCELL_X32 FILLER_90_1895 ();
 FILLCELL_X32 FILLER_90_1927 ();
 FILLCELL_X32 FILLER_90_1959 ();
 FILLCELL_X32 FILLER_90_1991 ();
 FILLCELL_X32 FILLER_90_2023 ();
 FILLCELL_X32 FILLER_90_2055 ();
 FILLCELL_X16 FILLER_90_2087 ();
 FILLCELL_X8 FILLER_90_2103 ();
 FILLCELL_X4 FILLER_90_2111 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X32 FILLER_91_1584 ();
 FILLCELL_X32 FILLER_91_1616 ();
 FILLCELL_X32 FILLER_91_1648 ();
 FILLCELL_X32 FILLER_91_1680 ();
 FILLCELL_X32 FILLER_91_1712 ();
 FILLCELL_X32 FILLER_91_1744 ();
 FILLCELL_X32 FILLER_91_1776 ();
 FILLCELL_X32 FILLER_91_1808 ();
 FILLCELL_X32 FILLER_91_1840 ();
 FILLCELL_X32 FILLER_91_1872 ();
 FILLCELL_X32 FILLER_91_1904 ();
 FILLCELL_X32 FILLER_91_1936 ();
 FILLCELL_X32 FILLER_91_1968 ();
 FILLCELL_X32 FILLER_91_2000 ();
 FILLCELL_X32 FILLER_91_2032 ();
 FILLCELL_X32 FILLER_91_2064 ();
 FILLCELL_X16 FILLER_91_2096 ();
 FILLCELL_X2 FILLER_91_2112 ();
 FILLCELL_X1 FILLER_91_2114 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X32 FILLER_92_1592 ();
 FILLCELL_X32 FILLER_92_1624 ();
 FILLCELL_X32 FILLER_92_1656 ();
 FILLCELL_X32 FILLER_92_1688 ();
 FILLCELL_X32 FILLER_92_1720 ();
 FILLCELL_X32 FILLER_92_1752 ();
 FILLCELL_X32 FILLER_92_1784 ();
 FILLCELL_X32 FILLER_92_1816 ();
 FILLCELL_X32 FILLER_92_1848 ();
 FILLCELL_X8 FILLER_92_1880 ();
 FILLCELL_X4 FILLER_92_1888 ();
 FILLCELL_X2 FILLER_92_1892 ();
 FILLCELL_X32 FILLER_92_1895 ();
 FILLCELL_X32 FILLER_92_1927 ();
 FILLCELL_X32 FILLER_92_1959 ();
 FILLCELL_X32 FILLER_92_1991 ();
 FILLCELL_X32 FILLER_92_2023 ();
 FILLCELL_X32 FILLER_92_2055 ();
 FILLCELL_X16 FILLER_92_2087 ();
 FILLCELL_X8 FILLER_92_2103 ();
 FILLCELL_X4 FILLER_92_2111 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X32 FILLER_93_1584 ();
 FILLCELL_X32 FILLER_93_1616 ();
 FILLCELL_X32 FILLER_93_1648 ();
 FILLCELL_X32 FILLER_93_1680 ();
 FILLCELL_X32 FILLER_93_1712 ();
 FILLCELL_X32 FILLER_93_1744 ();
 FILLCELL_X32 FILLER_93_1776 ();
 FILLCELL_X32 FILLER_93_1808 ();
 FILLCELL_X32 FILLER_93_1840 ();
 FILLCELL_X32 FILLER_93_1872 ();
 FILLCELL_X32 FILLER_93_1904 ();
 FILLCELL_X32 FILLER_93_1936 ();
 FILLCELL_X32 FILLER_93_1968 ();
 FILLCELL_X32 FILLER_93_2000 ();
 FILLCELL_X32 FILLER_93_2032 ();
 FILLCELL_X32 FILLER_93_2064 ();
 FILLCELL_X16 FILLER_93_2096 ();
 FILLCELL_X2 FILLER_93_2112 ();
 FILLCELL_X1 FILLER_93_2114 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X32 FILLER_94_1592 ();
 FILLCELL_X32 FILLER_94_1624 ();
 FILLCELL_X32 FILLER_94_1656 ();
 FILLCELL_X32 FILLER_94_1688 ();
 FILLCELL_X32 FILLER_94_1720 ();
 FILLCELL_X32 FILLER_94_1752 ();
 FILLCELL_X32 FILLER_94_1784 ();
 FILLCELL_X32 FILLER_94_1816 ();
 FILLCELL_X32 FILLER_94_1848 ();
 FILLCELL_X8 FILLER_94_1880 ();
 FILLCELL_X4 FILLER_94_1888 ();
 FILLCELL_X2 FILLER_94_1892 ();
 FILLCELL_X32 FILLER_94_1895 ();
 FILLCELL_X32 FILLER_94_1927 ();
 FILLCELL_X32 FILLER_94_1959 ();
 FILLCELL_X32 FILLER_94_1991 ();
 FILLCELL_X32 FILLER_94_2023 ();
 FILLCELL_X32 FILLER_94_2055 ();
 FILLCELL_X16 FILLER_94_2087 ();
 FILLCELL_X8 FILLER_94_2103 ();
 FILLCELL_X4 FILLER_94_2111 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X32 FILLER_95_961 ();
 FILLCELL_X32 FILLER_95_993 ();
 FILLCELL_X32 FILLER_95_1025 ();
 FILLCELL_X32 FILLER_95_1057 ();
 FILLCELL_X32 FILLER_95_1089 ();
 FILLCELL_X32 FILLER_95_1121 ();
 FILLCELL_X32 FILLER_95_1153 ();
 FILLCELL_X32 FILLER_95_1185 ();
 FILLCELL_X32 FILLER_95_1217 ();
 FILLCELL_X8 FILLER_95_1249 ();
 FILLCELL_X4 FILLER_95_1257 ();
 FILLCELL_X2 FILLER_95_1261 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X32 FILLER_95_1584 ();
 FILLCELL_X32 FILLER_95_1616 ();
 FILLCELL_X32 FILLER_95_1648 ();
 FILLCELL_X32 FILLER_95_1680 ();
 FILLCELL_X32 FILLER_95_1712 ();
 FILLCELL_X32 FILLER_95_1744 ();
 FILLCELL_X32 FILLER_95_1776 ();
 FILLCELL_X32 FILLER_95_1808 ();
 FILLCELL_X32 FILLER_95_1840 ();
 FILLCELL_X32 FILLER_95_1872 ();
 FILLCELL_X32 FILLER_95_1904 ();
 FILLCELL_X32 FILLER_95_1936 ();
 FILLCELL_X32 FILLER_95_1968 ();
 FILLCELL_X32 FILLER_95_2000 ();
 FILLCELL_X32 FILLER_95_2032 ();
 FILLCELL_X32 FILLER_95_2064 ();
 FILLCELL_X16 FILLER_95_2096 ();
 FILLCELL_X2 FILLER_95_2112 ();
 FILLCELL_X1 FILLER_95_2114 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X32 FILLER_96_1592 ();
 FILLCELL_X32 FILLER_96_1624 ();
 FILLCELL_X32 FILLER_96_1656 ();
 FILLCELL_X32 FILLER_96_1688 ();
 FILLCELL_X32 FILLER_96_1720 ();
 FILLCELL_X32 FILLER_96_1752 ();
 FILLCELL_X32 FILLER_96_1784 ();
 FILLCELL_X32 FILLER_96_1816 ();
 FILLCELL_X32 FILLER_96_1848 ();
 FILLCELL_X8 FILLER_96_1880 ();
 FILLCELL_X4 FILLER_96_1888 ();
 FILLCELL_X2 FILLER_96_1892 ();
 FILLCELL_X32 FILLER_96_1895 ();
 FILLCELL_X32 FILLER_96_1927 ();
 FILLCELL_X32 FILLER_96_1959 ();
 FILLCELL_X32 FILLER_96_1991 ();
 FILLCELL_X32 FILLER_96_2023 ();
 FILLCELL_X32 FILLER_96_2055 ();
 FILLCELL_X16 FILLER_96_2087 ();
 FILLCELL_X8 FILLER_96_2103 ();
 FILLCELL_X4 FILLER_96_2111 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X32 FILLER_97_961 ();
 FILLCELL_X32 FILLER_97_993 ();
 FILLCELL_X32 FILLER_97_1025 ();
 FILLCELL_X32 FILLER_97_1057 ();
 FILLCELL_X32 FILLER_97_1089 ();
 FILLCELL_X32 FILLER_97_1121 ();
 FILLCELL_X32 FILLER_97_1153 ();
 FILLCELL_X32 FILLER_97_1185 ();
 FILLCELL_X32 FILLER_97_1217 ();
 FILLCELL_X8 FILLER_97_1249 ();
 FILLCELL_X4 FILLER_97_1257 ();
 FILLCELL_X2 FILLER_97_1261 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X32 FILLER_97_1584 ();
 FILLCELL_X32 FILLER_97_1616 ();
 FILLCELL_X32 FILLER_97_1648 ();
 FILLCELL_X32 FILLER_97_1680 ();
 FILLCELL_X32 FILLER_97_1712 ();
 FILLCELL_X32 FILLER_97_1744 ();
 FILLCELL_X32 FILLER_97_1776 ();
 FILLCELL_X32 FILLER_97_1808 ();
 FILLCELL_X32 FILLER_97_1840 ();
 FILLCELL_X32 FILLER_97_1872 ();
 FILLCELL_X32 FILLER_97_1904 ();
 FILLCELL_X32 FILLER_97_1936 ();
 FILLCELL_X32 FILLER_97_1968 ();
 FILLCELL_X32 FILLER_97_2000 ();
 FILLCELL_X32 FILLER_97_2032 ();
 FILLCELL_X32 FILLER_97_2064 ();
 FILLCELL_X16 FILLER_97_2096 ();
 FILLCELL_X2 FILLER_97_2112 ();
 FILLCELL_X1 FILLER_97_2114 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X32 FILLER_98_1304 ();
 FILLCELL_X32 FILLER_98_1336 ();
 FILLCELL_X32 FILLER_98_1368 ();
 FILLCELL_X32 FILLER_98_1400 ();
 FILLCELL_X32 FILLER_98_1432 ();
 FILLCELL_X32 FILLER_98_1464 ();
 FILLCELL_X32 FILLER_98_1496 ();
 FILLCELL_X32 FILLER_98_1528 ();
 FILLCELL_X32 FILLER_98_1560 ();
 FILLCELL_X32 FILLER_98_1592 ();
 FILLCELL_X32 FILLER_98_1624 ();
 FILLCELL_X32 FILLER_98_1656 ();
 FILLCELL_X32 FILLER_98_1688 ();
 FILLCELL_X32 FILLER_98_1720 ();
 FILLCELL_X32 FILLER_98_1752 ();
 FILLCELL_X32 FILLER_98_1784 ();
 FILLCELL_X32 FILLER_98_1816 ();
 FILLCELL_X32 FILLER_98_1848 ();
 FILLCELL_X8 FILLER_98_1880 ();
 FILLCELL_X4 FILLER_98_1888 ();
 FILLCELL_X2 FILLER_98_1892 ();
 FILLCELL_X32 FILLER_98_1895 ();
 FILLCELL_X32 FILLER_98_1927 ();
 FILLCELL_X32 FILLER_98_1959 ();
 FILLCELL_X32 FILLER_98_1991 ();
 FILLCELL_X32 FILLER_98_2023 ();
 FILLCELL_X32 FILLER_98_2055 ();
 FILLCELL_X16 FILLER_98_2087 ();
 FILLCELL_X8 FILLER_98_2103 ();
 FILLCELL_X4 FILLER_98_2111 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X32 FILLER_99_1584 ();
 FILLCELL_X32 FILLER_99_1616 ();
 FILLCELL_X32 FILLER_99_1648 ();
 FILLCELL_X32 FILLER_99_1680 ();
 FILLCELL_X32 FILLER_99_1712 ();
 FILLCELL_X32 FILLER_99_1744 ();
 FILLCELL_X32 FILLER_99_1776 ();
 FILLCELL_X32 FILLER_99_1808 ();
 FILLCELL_X32 FILLER_99_1840 ();
 FILLCELL_X32 FILLER_99_1872 ();
 FILLCELL_X32 FILLER_99_1904 ();
 FILLCELL_X32 FILLER_99_1936 ();
 FILLCELL_X32 FILLER_99_1968 ();
 FILLCELL_X32 FILLER_99_2000 ();
 FILLCELL_X32 FILLER_99_2032 ();
 FILLCELL_X32 FILLER_99_2064 ();
 FILLCELL_X16 FILLER_99_2096 ();
 FILLCELL_X2 FILLER_99_2112 ();
 FILLCELL_X1 FILLER_99_2114 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X32 FILLER_100_952 ();
 FILLCELL_X32 FILLER_100_984 ();
 FILLCELL_X32 FILLER_100_1016 ();
 FILLCELL_X32 FILLER_100_1048 ();
 FILLCELL_X32 FILLER_100_1080 ();
 FILLCELL_X32 FILLER_100_1112 ();
 FILLCELL_X32 FILLER_100_1144 ();
 FILLCELL_X32 FILLER_100_1176 ();
 FILLCELL_X32 FILLER_100_1208 ();
 FILLCELL_X32 FILLER_100_1240 ();
 FILLCELL_X32 FILLER_100_1272 ();
 FILLCELL_X32 FILLER_100_1304 ();
 FILLCELL_X32 FILLER_100_1336 ();
 FILLCELL_X32 FILLER_100_1368 ();
 FILLCELL_X32 FILLER_100_1400 ();
 FILLCELL_X32 FILLER_100_1432 ();
 FILLCELL_X32 FILLER_100_1464 ();
 FILLCELL_X32 FILLER_100_1496 ();
 FILLCELL_X32 FILLER_100_1528 ();
 FILLCELL_X32 FILLER_100_1560 ();
 FILLCELL_X32 FILLER_100_1592 ();
 FILLCELL_X32 FILLER_100_1624 ();
 FILLCELL_X32 FILLER_100_1656 ();
 FILLCELL_X32 FILLER_100_1688 ();
 FILLCELL_X32 FILLER_100_1720 ();
 FILLCELL_X32 FILLER_100_1752 ();
 FILLCELL_X32 FILLER_100_1784 ();
 FILLCELL_X32 FILLER_100_1816 ();
 FILLCELL_X32 FILLER_100_1848 ();
 FILLCELL_X8 FILLER_100_1880 ();
 FILLCELL_X4 FILLER_100_1888 ();
 FILLCELL_X2 FILLER_100_1892 ();
 FILLCELL_X32 FILLER_100_1895 ();
 FILLCELL_X32 FILLER_100_1927 ();
 FILLCELL_X32 FILLER_100_1959 ();
 FILLCELL_X32 FILLER_100_1991 ();
 FILLCELL_X32 FILLER_100_2023 ();
 FILLCELL_X32 FILLER_100_2055 ();
 FILLCELL_X16 FILLER_100_2087 ();
 FILLCELL_X8 FILLER_100_2103 ();
 FILLCELL_X4 FILLER_100_2111 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X32 FILLER_101_1584 ();
 FILLCELL_X32 FILLER_101_1616 ();
 FILLCELL_X32 FILLER_101_1648 ();
 FILLCELL_X32 FILLER_101_1680 ();
 FILLCELL_X32 FILLER_101_1712 ();
 FILLCELL_X32 FILLER_101_1744 ();
 FILLCELL_X32 FILLER_101_1776 ();
 FILLCELL_X32 FILLER_101_1808 ();
 FILLCELL_X32 FILLER_101_1840 ();
 FILLCELL_X32 FILLER_101_1872 ();
 FILLCELL_X32 FILLER_101_1904 ();
 FILLCELL_X32 FILLER_101_1936 ();
 FILLCELL_X32 FILLER_101_1968 ();
 FILLCELL_X32 FILLER_101_2000 ();
 FILLCELL_X32 FILLER_101_2032 ();
 FILLCELL_X32 FILLER_101_2064 ();
 FILLCELL_X16 FILLER_101_2096 ();
 FILLCELL_X2 FILLER_101_2112 ();
 FILLCELL_X1 FILLER_101_2114 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X32 FILLER_102_1304 ();
 FILLCELL_X32 FILLER_102_1336 ();
 FILLCELL_X32 FILLER_102_1368 ();
 FILLCELL_X32 FILLER_102_1400 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X32 FILLER_102_1496 ();
 FILLCELL_X32 FILLER_102_1528 ();
 FILLCELL_X32 FILLER_102_1560 ();
 FILLCELL_X32 FILLER_102_1592 ();
 FILLCELL_X32 FILLER_102_1624 ();
 FILLCELL_X32 FILLER_102_1656 ();
 FILLCELL_X32 FILLER_102_1688 ();
 FILLCELL_X32 FILLER_102_1720 ();
 FILLCELL_X32 FILLER_102_1752 ();
 FILLCELL_X32 FILLER_102_1784 ();
 FILLCELL_X32 FILLER_102_1816 ();
 FILLCELL_X32 FILLER_102_1848 ();
 FILLCELL_X8 FILLER_102_1880 ();
 FILLCELL_X4 FILLER_102_1888 ();
 FILLCELL_X2 FILLER_102_1892 ();
 FILLCELL_X32 FILLER_102_1895 ();
 FILLCELL_X32 FILLER_102_1927 ();
 FILLCELL_X32 FILLER_102_1959 ();
 FILLCELL_X32 FILLER_102_1991 ();
 FILLCELL_X32 FILLER_102_2023 ();
 FILLCELL_X32 FILLER_102_2055 ();
 FILLCELL_X16 FILLER_102_2087 ();
 FILLCELL_X8 FILLER_102_2103 ();
 FILLCELL_X4 FILLER_102_2111 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X32 FILLER_103_1584 ();
 FILLCELL_X32 FILLER_103_1616 ();
 FILLCELL_X32 FILLER_103_1648 ();
 FILLCELL_X32 FILLER_103_1680 ();
 FILLCELL_X32 FILLER_103_1712 ();
 FILLCELL_X32 FILLER_103_1744 ();
 FILLCELL_X32 FILLER_103_1776 ();
 FILLCELL_X32 FILLER_103_1808 ();
 FILLCELL_X32 FILLER_103_1840 ();
 FILLCELL_X32 FILLER_103_1872 ();
 FILLCELL_X32 FILLER_103_1904 ();
 FILLCELL_X32 FILLER_103_1936 ();
 FILLCELL_X32 FILLER_103_1968 ();
 FILLCELL_X32 FILLER_103_2000 ();
 FILLCELL_X32 FILLER_103_2032 ();
 FILLCELL_X32 FILLER_103_2064 ();
 FILLCELL_X16 FILLER_103_2096 ();
 FILLCELL_X2 FILLER_103_2112 ();
 FILLCELL_X1 FILLER_103_2114 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X32 FILLER_104_1304 ();
 FILLCELL_X32 FILLER_104_1336 ();
 FILLCELL_X32 FILLER_104_1368 ();
 FILLCELL_X32 FILLER_104_1400 ();
 FILLCELL_X32 FILLER_104_1432 ();
 FILLCELL_X32 FILLER_104_1464 ();
 FILLCELL_X32 FILLER_104_1496 ();
 FILLCELL_X32 FILLER_104_1528 ();
 FILLCELL_X32 FILLER_104_1560 ();
 FILLCELL_X32 FILLER_104_1592 ();
 FILLCELL_X32 FILLER_104_1624 ();
 FILLCELL_X32 FILLER_104_1656 ();
 FILLCELL_X32 FILLER_104_1688 ();
 FILLCELL_X32 FILLER_104_1720 ();
 FILLCELL_X32 FILLER_104_1752 ();
 FILLCELL_X32 FILLER_104_1784 ();
 FILLCELL_X32 FILLER_104_1816 ();
 FILLCELL_X32 FILLER_104_1848 ();
 FILLCELL_X8 FILLER_104_1880 ();
 FILLCELL_X4 FILLER_104_1888 ();
 FILLCELL_X2 FILLER_104_1892 ();
 FILLCELL_X32 FILLER_104_1895 ();
 FILLCELL_X32 FILLER_104_1927 ();
 FILLCELL_X32 FILLER_104_1959 ();
 FILLCELL_X32 FILLER_104_1991 ();
 FILLCELL_X32 FILLER_104_2023 ();
 FILLCELL_X32 FILLER_104_2055 ();
 FILLCELL_X16 FILLER_104_2087 ();
 FILLCELL_X8 FILLER_104_2103 ();
 FILLCELL_X4 FILLER_104_2111 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X32 FILLER_105_961 ();
 FILLCELL_X32 FILLER_105_993 ();
 FILLCELL_X32 FILLER_105_1025 ();
 FILLCELL_X32 FILLER_105_1057 ();
 FILLCELL_X32 FILLER_105_1089 ();
 FILLCELL_X32 FILLER_105_1121 ();
 FILLCELL_X32 FILLER_105_1153 ();
 FILLCELL_X32 FILLER_105_1185 ();
 FILLCELL_X32 FILLER_105_1217 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X32 FILLER_105_1584 ();
 FILLCELL_X32 FILLER_105_1616 ();
 FILLCELL_X32 FILLER_105_1648 ();
 FILLCELL_X32 FILLER_105_1680 ();
 FILLCELL_X32 FILLER_105_1712 ();
 FILLCELL_X32 FILLER_105_1744 ();
 FILLCELL_X32 FILLER_105_1776 ();
 FILLCELL_X32 FILLER_105_1808 ();
 FILLCELL_X32 FILLER_105_1840 ();
 FILLCELL_X32 FILLER_105_1872 ();
 FILLCELL_X32 FILLER_105_1904 ();
 FILLCELL_X32 FILLER_105_1936 ();
 FILLCELL_X32 FILLER_105_1968 ();
 FILLCELL_X32 FILLER_105_2000 ();
 FILLCELL_X32 FILLER_105_2032 ();
 FILLCELL_X32 FILLER_105_2064 ();
 FILLCELL_X16 FILLER_105_2096 ();
 FILLCELL_X2 FILLER_105_2112 ();
 FILLCELL_X1 FILLER_105_2114 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X32 FILLER_106_1304 ();
 FILLCELL_X32 FILLER_106_1336 ();
 FILLCELL_X32 FILLER_106_1368 ();
 FILLCELL_X32 FILLER_106_1400 ();
 FILLCELL_X32 FILLER_106_1432 ();
 FILLCELL_X32 FILLER_106_1464 ();
 FILLCELL_X32 FILLER_106_1496 ();
 FILLCELL_X32 FILLER_106_1528 ();
 FILLCELL_X32 FILLER_106_1560 ();
 FILLCELL_X32 FILLER_106_1592 ();
 FILLCELL_X32 FILLER_106_1624 ();
 FILLCELL_X32 FILLER_106_1656 ();
 FILLCELL_X32 FILLER_106_1688 ();
 FILLCELL_X32 FILLER_106_1720 ();
 FILLCELL_X32 FILLER_106_1752 ();
 FILLCELL_X32 FILLER_106_1784 ();
 FILLCELL_X32 FILLER_106_1816 ();
 FILLCELL_X32 FILLER_106_1848 ();
 FILLCELL_X8 FILLER_106_1880 ();
 FILLCELL_X4 FILLER_106_1888 ();
 FILLCELL_X2 FILLER_106_1892 ();
 FILLCELL_X32 FILLER_106_1895 ();
 FILLCELL_X32 FILLER_106_1927 ();
 FILLCELL_X32 FILLER_106_1959 ();
 FILLCELL_X32 FILLER_106_1991 ();
 FILLCELL_X32 FILLER_106_2023 ();
 FILLCELL_X32 FILLER_106_2055 ();
 FILLCELL_X16 FILLER_106_2087 ();
 FILLCELL_X8 FILLER_106_2103 ();
 FILLCELL_X4 FILLER_106_2111 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X32 FILLER_107_961 ();
 FILLCELL_X32 FILLER_107_993 ();
 FILLCELL_X32 FILLER_107_1025 ();
 FILLCELL_X32 FILLER_107_1057 ();
 FILLCELL_X32 FILLER_107_1089 ();
 FILLCELL_X32 FILLER_107_1121 ();
 FILLCELL_X32 FILLER_107_1153 ();
 FILLCELL_X32 FILLER_107_1185 ();
 FILLCELL_X32 FILLER_107_1217 ();
 FILLCELL_X8 FILLER_107_1249 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X32 FILLER_107_1584 ();
 FILLCELL_X32 FILLER_107_1616 ();
 FILLCELL_X32 FILLER_107_1648 ();
 FILLCELL_X32 FILLER_107_1680 ();
 FILLCELL_X32 FILLER_107_1712 ();
 FILLCELL_X32 FILLER_107_1744 ();
 FILLCELL_X32 FILLER_107_1776 ();
 FILLCELL_X32 FILLER_107_1808 ();
 FILLCELL_X32 FILLER_107_1840 ();
 FILLCELL_X32 FILLER_107_1872 ();
 FILLCELL_X32 FILLER_107_1904 ();
 FILLCELL_X32 FILLER_107_1936 ();
 FILLCELL_X32 FILLER_107_1968 ();
 FILLCELL_X32 FILLER_107_2000 ();
 FILLCELL_X32 FILLER_107_2032 ();
 FILLCELL_X32 FILLER_107_2064 ();
 FILLCELL_X16 FILLER_107_2096 ();
 FILLCELL_X2 FILLER_107_2112 ();
 FILLCELL_X1 FILLER_107_2114 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X32 FILLER_108_856 ();
 FILLCELL_X32 FILLER_108_888 ();
 FILLCELL_X32 FILLER_108_920 ();
 FILLCELL_X32 FILLER_108_952 ();
 FILLCELL_X32 FILLER_108_984 ();
 FILLCELL_X32 FILLER_108_1016 ();
 FILLCELL_X32 FILLER_108_1048 ();
 FILLCELL_X32 FILLER_108_1080 ();
 FILLCELL_X32 FILLER_108_1112 ();
 FILLCELL_X32 FILLER_108_1144 ();
 FILLCELL_X32 FILLER_108_1176 ();
 FILLCELL_X32 FILLER_108_1208 ();
 FILLCELL_X32 FILLER_108_1240 ();
 FILLCELL_X32 FILLER_108_1272 ();
 FILLCELL_X32 FILLER_108_1304 ();
 FILLCELL_X32 FILLER_108_1336 ();
 FILLCELL_X32 FILLER_108_1368 ();
 FILLCELL_X32 FILLER_108_1400 ();
 FILLCELL_X32 FILLER_108_1432 ();
 FILLCELL_X32 FILLER_108_1464 ();
 FILLCELL_X32 FILLER_108_1496 ();
 FILLCELL_X32 FILLER_108_1528 ();
 FILLCELL_X32 FILLER_108_1560 ();
 FILLCELL_X32 FILLER_108_1592 ();
 FILLCELL_X32 FILLER_108_1624 ();
 FILLCELL_X32 FILLER_108_1656 ();
 FILLCELL_X32 FILLER_108_1688 ();
 FILLCELL_X32 FILLER_108_1720 ();
 FILLCELL_X32 FILLER_108_1752 ();
 FILLCELL_X32 FILLER_108_1784 ();
 FILLCELL_X32 FILLER_108_1816 ();
 FILLCELL_X32 FILLER_108_1848 ();
 FILLCELL_X8 FILLER_108_1880 ();
 FILLCELL_X4 FILLER_108_1888 ();
 FILLCELL_X2 FILLER_108_1892 ();
 FILLCELL_X32 FILLER_108_1895 ();
 FILLCELL_X32 FILLER_108_1927 ();
 FILLCELL_X32 FILLER_108_1959 ();
 FILLCELL_X32 FILLER_108_1991 ();
 FILLCELL_X32 FILLER_108_2023 ();
 FILLCELL_X32 FILLER_108_2055 ();
 FILLCELL_X16 FILLER_108_2087 ();
 FILLCELL_X8 FILLER_108_2103 ();
 FILLCELL_X4 FILLER_108_2111 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X32 FILLER_109_1584 ();
 FILLCELL_X32 FILLER_109_1616 ();
 FILLCELL_X32 FILLER_109_1648 ();
 FILLCELL_X32 FILLER_109_1680 ();
 FILLCELL_X32 FILLER_109_1712 ();
 FILLCELL_X32 FILLER_109_1744 ();
 FILLCELL_X32 FILLER_109_1776 ();
 FILLCELL_X32 FILLER_109_1808 ();
 FILLCELL_X32 FILLER_109_1840 ();
 FILLCELL_X32 FILLER_109_1872 ();
 FILLCELL_X32 FILLER_109_1904 ();
 FILLCELL_X32 FILLER_109_1936 ();
 FILLCELL_X32 FILLER_109_1968 ();
 FILLCELL_X32 FILLER_109_2000 ();
 FILLCELL_X32 FILLER_109_2032 ();
 FILLCELL_X32 FILLER_109_2064 ();
 FILLCELL_X16 FILLER_109_2096 ();
 FILLCELL_X2 FILLER_109_2112 ();
 FILLCELL_X1 FILLER_109_2114 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X32 FILLER_110_952 ();
 FILLCELL_X32 FILLER_110_984 ();
 FILLCELL_X32 FILLER_110_1016 ();
 FILLCELL_X32 FILLER_110_1048 ();
 FILLCELL_X32 FILLER_110_1080 ();
 FILLCELL_X32 FILLER_110_1112 ();
 FILLCELL_X32 FILLER_110_1144 ();
 FILLCELL_X32 FILLER_110_1176 ();
 FILLCELL_X32 FILLER_110_1208 ();
 FILLCELL_X32 FILLER_110_1240 ();
 FILLCELL_X32 FILLER_110_1272 ();
 FILLCELL_X32 FILLER_110_1304 ();
 FILLCELL_X32 FILLER_110_1336 ();
 FILLCELL_X32 FILLER_110_1368 ();
 FILLCELL_X32 FILLER_110_1400 ();
 FILLCELL_X32 FILLER_110_1432 ();
 FILLCELL_X32 FILLER_110_1464 ();
 FILLCELL_X32 FILLER_110_1496 ();
 FILLCELL_X32 FILLER_110_1528 ();
 FILLCELL_X32 FILLER_110_1560 ();
 FILLCELL_X32 FILLER_110_1592 ();
 FILLCELL_X32 FILLER_110_1624 ();
 FILLCELL_X32 FILLER_110_1656 ();
 FILLCELL_X32 FILLER_110_1688 ();
 FILLCELL_X32 FILLER_110_1720 ();
 FILLCELL_X32 FILLER_110_1752 ();
 FILLCELL_X32 FILLER_110_1784 ();
 FILLCELL_X32 FILLER_110_1816 ();
 FILLCELL_X32 FILLER_110_1848 ();
 FILLCELL_X8 FILLER_110_1880 ();
 FILLCELL_X4 FILLER_110_1888 ();
 FILLCELL_X2 FILLER_110_1892 ();
 FILLCELL_X32 FILLER_110_1895 ();
 FILLCELL_X32 FILLER_110_1927 ();
 FILLCELL_X32 FILLER_110_1959 ();
 FILLCELL_X32 FILLER_110_1991 ();
 FILLCELL_X32 FILLER_110_2023 ();
 FILLCELL_X32 FILLER_110_2055 ();
 FILLCELL_X16 FILLER_110_2087 ();
 FILLCELL_X8 FILLER_110_2103 ();
 FILLCELL_X4 FILLER_110_2111 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X32 FILLER_111_961 ();
 FILLCELL_X32 FILLER_111_993 ();
 FILLCELL_X32 FILLER_111_1025 ();
 FILLCELL_X32 FILLER_111_1057 ();
 FILLCELL_X32 FILLER_111_1089 ();
 FILLCELL_X32 FILLER_111_1121 ();
 FILLCELL_X32 FILLER_111_1153 ();
 FILLCELL_X32 FILLER_111_1185 ();
 FILLCELL_X32 FILLER_111_1217 ();
 FILLCELL_X8 FILLER_111_1249 ();
 FILLCELL_X4 FILLER_111_1257 ();
 FILLCELL_X2 FILLER_111_1261 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X32 FILLER_111_1584 ();
 FILLCELL_X32 FILLER_111_1616 ();
 FILLCELL_X32 FILLER_111_1648 ();
 FILLCELL_X32 FILLER_111_1680 ();
 FILLCELL_X32 FILLER_111_1712 ();
 FILLCELL_X32 FILLER_111_1744 ();
 FILLCELL_X32 FILLER_111_1776 ();
 FILLCELL_X32 FILLER_111_1808 ();
 FILLCELL_X32 FILLER_111_1840 ();
 FILLCELL_X32 FILLER_111_1872 ();
 FILLCELL_X32 FILLER_111_1904 ();
 FILLCELL_X32 FILLER_111_1936 ();
 FILLCELL_X32 FILLER_111_1968 ();
 FILLCELL_X32 FILLER_111_2000 ();
 FILLCELL_X32 FILLER_111_2032 ();
 FILLCELL_X32 FILLER_111_2064 ();
 FILLCELL_X16 FILLER_111_2096 ();
 FILLCELL_X2 FILLER_111_2112 ();
 FILLCELL_X1 FILLER_111_2114 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X32 FILLER_112_952 ();
 FILLCELL_X32 FILLER_112_984 ();
 FILLCELL_X32 FILLER_112_1016 ();
 FILLCELL_X32 FILLER_112_1048 ();
 FILLCELL_X32 FILLER_112_1080 ();
 FILLCELL_X32 FILLER_112_1112 ();
 FILLCELL_X32 FILLER_112_1144 ();
 FILLCELL_X32 FILLER_112_1176 ();
 FILLCELL_X32 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_112_1240 ();
 FILLCELL_X32 FILLER_112_1272 ();
 FILLCELL_X32 FILLER_112_1304 ();
 FILLCELL_X32 FILLER_112_1336 ();
 FILLCELL_X32 FILLER_112_1368 ();
 FILLCELL_X32 FILLER_112_1400 ();
 FILLCELL_X32 FILLER_112_1432 ();
 FILLCELL_X32 FILLER_112_1464 ();
 FILLCELL_X32 FILLER_112_1496 ();
 FILLCELL_X32 FILLER_112_1528 ();
 FILLCELL_X32 FILLER_112_1560 ();
 FILLCELL_X32 FILLER_112_1592 ();
 FILLCELL_X32 FILLER_112_1624 ();
 FILLCELL_X32 FILLER_112_1656 ();
 FILLCELL_X32 FILLER_112_1688 ();
 FILLCELL_X32 FILLER_112_1720 ();
 FILLCELL_X32 FILLER_112_1752 ();
 FILLCELL_X32 FILLER_112_1784 ();
 FILLCELL_X32 FILLER_112_1816 ();
 FILLCELL_X32 FILLER_112_1848 ();
 FILLCELL_X8 FILLER_112_1880 ();
 FILLCELL_X4 FILLER_112_1888 ();
 FILLCELL_X2 FILLER_112_1892 ();
 FILLCELL_X32 FILLER_112_1895 ();
 FILLCELL_X32 FILLER_112_1927 ();
 FILLCELL_X32 FILLER_112_1959 ();
 FILLCELL_X32 FILLER_112_1991 ();
 FILLCELL_X32 FILLER_112_2023 ();
 FILLCELL_X32 FILLER_112_2055 ();
 FILLCELL_X16 FILLER_112_2087 ();
 FILLCELL_X8 FILLER_112_2103 ();
 FILLCELL_X4 FILLER_112_2111 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X32 FILLER_113_833 ();
 FILLCELL_X32 FILLER_113_865 ();
 FILLCELL_X32 FILLER_113_897 ();
 FILLCELL_X32 FILLER_113_929 ();
 FILLCELL_X32 FILLER_113_961 ();
 FILLCELL_X32 FILLER_113_993 ();
 FILLCELL_X32 FILLER_113_1025 ();
 FILLCELL_X32 FILLER_113_1057 ();
 FILLCELL_X32 FILLER_113_1089 ();
 FILLCELL_X32 FILLER_113_1121 ();
 FILLCELL_X32 FILLER_113_1153 ();
 FILLCELL_X32 FILLER_113_1185 ();
 FILLCELL_X32 FILLER_113_1217 ();
 FILLCELL_X8 FILLER_113_1249 ();
 FILLCELL_X4 FILLER_113_1257 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X32 FILLER_113_1552 ();
 FILLCELL_X32 FILLER_113_1584 ();
 FILLCELL_X32 FILLER_113_1616 ();
 FILLCELL_X32 FILLER_113_1648 ();
 FILLCELL_X32 FILLER_113_1680 ();
 FILLCELL_X32 FILLER_113_1712 ();
 FILLCELL_X32 FILLER_113_1744 ();
 FILLCELL_X32 FILLER_113_1776 ();
 FILLCELL_X32 FILLER_113_1808 ();
 FILLCELL_X32 FILLER_113_1840 ();
 FILLCELL_X32 FILLER_113_1872 ();
 FILLCELL_X32 FILLER_113_1904 ();
 FILLCELL_X32 FILLER_113_1936 ();
 FILLCELL_X32 FILLER_113_1968 ();
 FILLCELL_X32 FILLER_113_2000 ();
 FILLCELL_X32 FILLER_113_2032 ();
 FILLCELL_X32 FILLER_113_2064 ();
 FILLCELL_X16 FILLER_113_2096 ();
 FILLCELL_X2 FILLER_113_2112 ();
 FILLCELL_X1 FILLER_113_2114 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X32 FILLER_114_952 ();
 FILLCELL_X32 FILLER_114_984 ();
 FILLCELL_X32 FILLER_114_1016 ();
 FILLCELL_X32 FILLER_114_1048 ();
 FILLCELL_X32 FILLER_114_1080 ();
 FILLCELL_X32 FILLER_114_1112 ();
 FILLCELL_X32 FILLER_114_1144 ();
 FILLCELL_X32 FILLER_114_1176 ();
 FILLCELL_X32 FILLER_114_1208 ();
 FILLCELL_X32 FILLER_114_1240 ();
 FILLCELL_X32 FILLER_114_1272 ();
 FILLCELL_X32 FILLER_114_1304 ();
 FILLCELL_X32 FILLER_114_1336 ();
 FILLCELL_X32 FILLER_114_1368 ();
 FILLCELL_X32 FILLER_114_1400 ();
 FILLCELL_X32 FILLER_114_1432 ();
 FILLCELL_X32 FILLER_114_1464 ();
 FILLCELL_X32 FILLER_114_1496 ();
 FILLCELL_X32 FILLER_114_1528 ();
 FILLCELL_X32 FILLER_114_1560 ();
 FILLCELL_X32 FILLER_114_1592 ();
 FILLCELL_X32 FILLER_114_1624 ();
 FILLCELL_X32 FILLER_114_1656 ();
 FILLCELL_X32 FILLER_114_1688 ();
 FILLCELL_X32 FILLER_114_1720 ();
 FILLCELL_X32 FILLER_114_1752 ();
 FILLCELL_X32 FILLER_114_1784 ();
 FILLCELL_X32 FILLER_114_1816 ();
 FILLCELL_X32 FILLER_114_1848 ();
 FILLCELL_X8 FILLER_114_1880 ();
 FILLCELL_X4 FILLER_114_1888 ();
 FILLCELL_X2 FILLER_114_1892 ();
 FILLCELL_X32 FILLER_114_1895 ();
 FILLCELL_X32 FILLER_114_1927 ();
 FILLCELL_X32 FILLER_114_1959 ();
 FILLCELL_X32 FILLER_114_1991 ();
 FILLCELL_X32 FILLER_114_2023 ();
 FILLCELL_X32 FILLER_114_2055 ();
 FILLCELL_X16 FILLER_114_2087 ();
 FILLCELL_X8 FILLER_114_2103 ();
 FILLCELL_X4 FILLER_114_2111 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X32 FILLER_115_801 ();
 FILLCELL_X32 FILLER_115_833 ();
 FILLCELL_X32 FILLER_115_865 ();
 FILLCELL_X32 FILLER_115_897 ();
 FILLCELL_X32 FILLER_115_929 ();
 FILLCELL_X32 FILLER_115_961 ();
 FILLCELL_X32 FILLER_115_993 ();
 FILLCELL_X32 FILLER_115_1025 ();
 FILLCELL_X32 FILLER_115_1057 ();
 FILLCELL_X32 FILLER_115_1089 ();
 FILLCELL_X32 FILLER_115_1121 ();
 FILLCELL_X32 FILLER_115_1153 ();
 FILLCELL_X32 FILLER_115_1185 ();
 FILLCELL_X32 FILLER_115_1217 ();
 FILLCELL_X8 FILLER_115_1249 ();
 FILLCELL_X4 FILLER_115_1257 ();
 FILLCELL_X2 FILLER_115_1261 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X32 FILLER_115_1552 ();
 FILLCELL_X32 FILLER_115_1584 ();
 FILLCELL_X32 FILLER_115_1616 ();
 FILLCELL_X32 FILLER_115_1648 ();
 FILLCELL_X32 FILLER_115_1680 ();
 FILLCELL_X32 FILLER_115_1712 ();
 FILLCELL_X32 FILLER_115_1744 ();
 FILLCELL_X32 FILLER_115_1776 ();
 FILLCELL_X32 FILLER_115_1808 ();
 FILLCELL_X32 FILLER_115_1840 ();
 FILLCELL_X32 FILLER_115_1872 ();
 FILLCELL_X32 FILLER_115_1904 ();
 FILLCELL_X32 FILLER_115_1936 ();
 FILLCELL_X32 FILLER_115_1968 ();
 FILLCELL_X32 FILLER_115_2000 ();
 FILLCELL_X32 FILLER_115_2032 ();
 FILLCELL_X32 FILLER_115_2064 ();
 FILLCELL_X16 FILLER_115_2096 ();
 FILLCELL_X2 FILLER_115_2112 ();
 FILLCELL_X1 FILLER_115_2114 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X32 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_888 ();
 FILLCELL_X32 FILLER_116_920 ();
 FILLCELL_X32 FILLER_116_952 ();
 FILLCELL_X32 FILLER_116_984 ();
 FILLCELL_X32 FILLER_116_1016 ();
 FILLCELL_X32 FILLER_116_1048 ();
 FILLCELL_X32 FILLER_116_1080 ();
 FILLCELL_X32 FILLER_116_1112 ();
 FILLCELL_X32 FILLER_116_1144 ();
 FILLCELL_X32 FILLER_116_1176 ();
 FILLCELL_X32 FILLER_116_1208 ();
 FILLCELL_X32 FILLER_116_1240 ();
 FILLCELL_X32 FILLER_116_1272 ();
 FILLCELL_X32 FILLER_116_1304 ();
 FILLCELL_X32 FILLER_116_1336 ();
 FILLCELL_X32 FILLER_116_1368 ();
 FILLCELL_X32 FILLER_116_1400 ();
 FILLCELL_X32 FILLER_116_1432 ();
 FILLCELL_X32 FILLER_116_1464 ();
 FILLCELL_X32 FILLER_116_1496 ();
 FILLCELL_X32 FILLER_116_1528 ();
 FILLCELL_X32 FILLER_116_1560 ();
 FILLCELL_X32 FILLER_116_1592 ();
 FILLCELL_X32 FILLER_116_1624 ();
 FILLCELL_X32 FILLER_116_1656 ();
 FILLCELL_X32 FILLER_116_1688 ();
 FILLCELL_X32 FILLER_116_1720 ();
 FILLCELL_X32 FILLER_116_1752 ();
 FILLCELL_X32 FILLER_116_1784 ();
 FILLCELL_X32 FILLER_116_1816 ();
 FILLCELL_X32 FILLER_116_1848 ();
 FILLCELL_X8 FILLER_116_1880 ();
 FILLCELL_X4 FILLER_116_1888 ();
 FILLCELL_X2 FILLER_116_1892 ();
 FILLCELL_X32 FILLER_116_1895 ();
 FILLCELL_X32 FILLER_116_1927 ();
 FILLCELL_X32 FILLER_116_1959 ();
 FILLCELL_X32 FILLER_116_1991 ();
 FILLCELL_X32 FILLER_116_2023 ();
 FILLCELL_X32 FILLER_116_2055 ();
 FILLCELL_X16 FILLER_116_2087 ();
 FILLCELL_X8 FILLER_116_2103 ();
 FILLCELL_X4 FILLER_116_2111 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X32 FILLER_117_801 ();
 FILLCELL_X32 FILLER_117_833 ();
 FILLCELL_X32 FILLER_117_865 ();
 FILLCELL_X32 FILLER_117_897 ();
 FILLCELL_X32 FILLER_117_929 ();
 FILLCELL_X32 FILLER_117_961 ();
 FILLCELL_X32 FILLER_117_993 ();
 FILLCELL_X32 FILLER_117_1025 ();
 FILLCELL_X32 FILLER_117_1057 ();
 FILLCELL_X32 FILLER_117_1089 ();
 FILLCELL_X32 FILLER_117_1121 ();
 FILLCELL_X32 FILLER_117_1153 ();
 FILLCELL_X32 FILLER_117_1185 ();
 FILLCELL_X32 FILLER_117_1217 ();
 FILLCELL_X8 FILLER_117_1249 ();
 FILLCELL_X4 FILLER_117_1257 ();
 FILLCELL_X2 FILLER_117_1261 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X32 FILLER_117_1552 ();
 FILLCELL_X32 FILLER_117_1584 ();
 FILLCELL_X32 FILLER_117_1616 ();
 FILLCELL_X32 FILLER_117_1648 ();
 FILLCELL_X32 FILLER_117_1680 ();
 FILLCELL_X32 FILLER_117_1712 ();
 FILLCELL_X32 FILLER_117_1744 ();
 FILLCELL_X32 FILLER_117_1776 ();
 FILLCELL_X32 FILLER_117_1808 ();
 FILLCELL_X32 FILLER_117_1840 ();
 FILLCELL_X32 FILLER_117_1872 ();
 FILLCELL_X32 FILLER_117_1904 ();
 FILLCELL_X32 FILLER_117_1936 ();
 FILLCELL_X32 FILLER_117_1968 ();
 FILLCELL_X32 FILLER_117_2000 ();
 FILLCELL_X32 FILLER_117_2032 ();
 FILLCELL_X32 FILLER_117_2064 ();
 FILLCELL_X16 FILLER_117_2096 ();
 FILLCELL_X2 FILLER_117_2112 ();
 FILLCELL_X1 FILLER_117_2114 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X32 FILLER_118_952 ();
 FILLCELL_X32 FILLER_118_984 ();
 FILLCELL_X32 FILLER_118_1016 ();
 FILLCELL_X32 FILLER_118_1048 ();
 FILLCELL_X32 FILLER_118_1080 ();
 FILLCELL_X32 FILLER_118_1112 ();
 FILLCELL_X32 FILLER_118_1144 ();
 FILLCELL_X32 FILLER_118_1176 ();
 FILLCELL_X32 FILLER_118_1208 ();
 FILLCELL_X32 FILLER_118_1240 ();
 FILLCELL_X32 FILLER_118_1272 ();
 FILLCELL_X32 FILLER_118_1304 ();
 FILLCELL_X32 FILLER_118_1336 ();
 FILLCELL_X32 FILLER_118_1368 ();
 FILLCELL_X32 FILLER_118_1400 ();
 FILLCELL_X32 FILLER_118_1432 ();
 FILLCELL_X32 FILLER_118_1464 ();
 FILLCELL_X32 FILLER_118_1496 ();
 FILLCELL_X32 FILLER_118_1528 ();
 FILLCELL_X32 FILLER_118_1560 ();
 FILLCELL_X32 FILLER_118_1592 ();
 FILLCELL_X32 FILLER_118_1624 ();
 FILLCELL_X32 FILLER_118_1656 ();
 FILLCELL_X32 FILLER_118_1688 ();
 FILLCELL_X32 FILLER_118_1720 ();
 FILLCELL_X32 FILLER_118_1752 ();
 FILLCELL_X32 FILLER_118_1784 ();
 FILLCELL_X32 FILLER_118_1816 ();
 FILLCELL_X32 FILLER_118_1848 ();
 FILLCELL_X8 FILLER_118_1880 ();
 FILLCELL_X4 FILLER_118_1888 ();
 FILLCELL_X2 FILLER_118_1892 ();
 FILLCELL_X32 FILLER_118_1895 ();
 FILLCELL_X32 FILLER_118_1927 ();
 FILLCELL_X32 FILLER_118_1959 ();
 FILLCELL_X32 FILLER_118_1991 ();
 FILLCELL_X32 FILLER_118_2023 ();
 FILLCELL_X32 FILLER_118_2055 ();
 FILLCELL_X16 FILLER_118_2087 ();
 FILLCELL_X8 FILLER_118_2103 ();
 FILLCELL_X4 FILLER_118_2111 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X32 FILLER_119_993 ();
 FILLCELL_X32 FILLER_119_1025 ();
 FILLCELL_X32 FILLER_119_1057 ();
 FILLCELL_X32 FILLER_119_1089 ();
 FILLCELL_X32 FILLER_119_1121 ();
 FILLCELL_X32 FILLER_119_1153 ();
 FILLCELL_X32 FILLER_119_1185 ();
 FILLCELL_X32 FILLER_119_1217 ();
 FILLCELL_X8 FILLER_119_1249 ();
 FILLCELL_X4 FILLER_119_1257 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X32 FILLER_119_1552 ();
 FILLCELL_X32 FILLER_119_1584 ();
 FILLCELL_X32 FILLER_119_1616 ();
 FILLCELL_X32 FILLER_119_1648 ();
 FILLCELL_X32 FILLER_119_1680 ();
 FILLCELL_X32 FILLER_119_1712 ();
 FILLCELL_X32 FILLER_119_1744 ();
 FILLCELL_X32 FILLER_119_1776 ();
 FILLCELL_X32 FILLER_119_1808 ();
 FILLCELL_X32 FILLER_119_1840 ();
 FILLCELL_X32 FILLER_119_1872 ();
 FILLCELL_X32 FILLER_119_1904 ();
 FILLCELL_X32 FILLER_119_1936 ();
 FILLCELL_X32 FILLER_119_1968 ();
 FILLCELL_X32 FILLER_119_2000 ();
 FILLCELL_X32 FILLER_119_2032 ();
 FILLCELL_X32 FILLER_119_2064 ();
 FILLCELL_X16 FILLER_119_2096 ();
 FILLCELL_X2 FILLER_119_2112 ();
 FILLCELL_X1 FILLER_119_2114 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X32 FILLER_120_984 ();
 FILLCELL_X32 FILLER_120_1016 ();
 FILLCELL_X32 FILLER_120_1048 ();
 FILLCELL_X32 FILLER_120_1080 ();
 FILLCELL_X32 FILLER_120_1112 ();
 FILLCELL_X32 FILLER_120_1144 ();
 FILLCELL_X32 FILLER_120_1176 ();
 FILLCELL_X32 FILLER_120_1208 ();
 FILLCELL_X32 FILLER_120_1240 ();
 FILLCELL_X32 FILLER_120_1272 ();
 FILLCELL_X32 FILLER_120_1304 ();
 FILLCELL_X32 FILLER_120_1336 ();
 FILLCELL_X32 FILLER_120_1368 ();
 FILLCELL_X32 FILLER_120_1400 ();
 FILLCELL_X32 FILLER_120_1432 ();
 FILLCELL_X32 FILLER_120_1464 ();
 FILLCELL_X32 FILLER_120_1496 ();
 FILLCELL_X32 FILLER_120_1528 ();
 FILLCELL_X32 FILLER_120_1560 ();
 FILLCELL_X32 FILLER_120_1592 ();
 FILLCELL_X32 FILLER_120_1624 ();
 FILLCELL_X32 FILLER_120_1656 ();
 FILLCELL_X32 FILLER_120_1688 ();
 FILLCELL_X32 FILLER_120_1720 ();
 FILLCELL_X32 FILLER_120_1752 ();
 FILLCELL_X32 FILLER_120_1784 ();
 FILLCELL_X32 FILLER_120_1816 ();
 FILLCELL_X32 FILLER_120_1848 ();
 FILLCELL_X8 FILLER_120_1880 ();
 FILLCELL_X4 FILLER_120_1888 ();
 FILLCELL_X2 FILLER_120_1892 ();
 FILLCELL_X32 FILLER_120_1895 ();
 FILLCELL_X32 FILLER_120_1927 ();
 FILLCELL_X32 FILLER_120_1959 ();
 FILLCELL_X32 FILLER_120_1991 ();
 FILLCELL_X32 FILLER_120_2023 ();
 FILLCELL_X32 FILLER_120_2055 ();
 FILLCELL_X16 FILLER_120_2087 ();
 FILLCELL_X8 FILLER_120_2103 ();
 FILLCELL_X4 FILLER_120_2111 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X32 FILLER_121_993 ();
 FILLCELL_X32 FILLER_121_1025 ();
 FILLCELL_X32 FILLER_121_1057 ();
 FILLCELL_X32 FILLER_121_1089 ();
 FILLCELL_X32 FILLER_121_1121 ();
 FILLCELL_X32 FILLER_121_1153 ();
 FILLCELL_X32 FILLER_121_1185 ();
 FILLCELL_X32 FILLER_121_1217 ();
 FILLCELL_X8 FILLER_121_1249 ();
 FILLCELL_X4 FILLER_121_1257 ();
 FILLCELL_X2 FILLER_121_1261 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X32 FILLER_121_1552 ();
 FILLCELL_X32 FILLER_121_1584 ();
 FILLCELL_X32 FILLER_121_1616 ();
 FILLCELL_X32 FILLER_121_1648 ();
 FILLCELL_X32 FILLER_121_1680 ();
 FILLCELL_X32 FILLER_121_1712 ();
 FILLCELL_X32 FILLER_121_1744 ();
 FILLCELL_X32 FILLER_121_1776 ();
 FILLCELL_X32 FILLER_121_1808 ();
 FILLCELL_X32 FILLER_121_1840 ();
 FILLCELL_X32 FILLER_121_1872 ();
 FILLCELL_X32 FILLER_121_1904 ();
 FILLCELL_X32 FILLER_121_1936 ();
 FILLCELL_X32 FILLER_121_1968 ();
 FILLCELL_X32 FILLER_121_2000 ();
 FILLCELL_X32 FILLER_121_2032 ();
 FILLCELL_X32 FILLER_121_2064 ();
 FILLCELL_X16 FILLER_121_2096 ();
 FILLCELL_X2 FILLER_121_2112 ();
 FILLCELL_X1 FILLER_121_2114 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X32 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_122_1048 ();
 FILLCELL_X32 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1112 ();
 FILLCELL_X32 FILLER_122_1144 ();
 FILLCELL_X32 FILLER_122_1176 ();
 FILLCELL_X32 FILLER_122_1208 ();
 FILLCELL_X32 FILLER_122_1240 ();
 FILLCELL_X32 FILLER_122_1272 ();
 FILLCELL_X32 FILLER_122_1304 ();
 FILLCELL_X32 FILLER_122_1336 ();
 FILLCELL_X32 FILLER_122_1368 ();
 FILLCELL_X32 FILLER_122_1400 ();
 FILLCELL_X32 FILLER_122_1432 ();
 FILLCELL_X32 FILLER_122_1464 ();
 FILLCELL_X32 FILLER_122_1496 ();
 FILLCELL_X32 FILLER_122_1528 ();
 FILLCELL_X32 FILLER_122_1560 ();
 FILLCELL_X32 FILLER_122_1592 ();
 FILLCELL_X32 FILLER_122_1624 ();
 FILLCELL_X32 FILLER_122_1656 ();
 FILLCELL_X32 FILLER_122_1688 ();
 FILLCELL_X32 FILLER_122_1720 ();
 FILLCELL_X32 FILLER_122_1752 ();
 FILLCELL_X32 FILLER_122_1784 ();
 FILLCELL_X32 FILLER_122_1816 ();
 FILLCELL_X32 FILLER_122_1848 ();
 FILLCELL_X8 FILLER_122_1880 ();
 FILLCELL_X4 FILLER_122_1888 ();
 FILLCELL_X2 FILLER_122_1892 ();
 FILLCELL_X32 FILLER_122_1895 ();
 FILLCELL_X32 FILLER_122_1927 ();
 FILLCELL_X32 FILLER_122_1959 ();
 FILLCELL_X32 FILLER_122_1991 ();
 FILLCELL_X32 FILLER_122_2023 ();
 FILLCELL_X32 FILLER_122_2055 ();
 FILLCELL_X16 FILLER_122_2087 ();
 FILLCELL_X8 FILLER_122_2103 ();
 FILLCELL_X4 FILLER_122_2111 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X32 FILLER_123_993 ();
 FILLCELL_X32 FILLER_123_1025 ();
 FILLCELL_X32 FILLER_123_1057 ();
 FILLCELL_X32 FILLER_123_1089 ();
 FILLCELL_X32 FILLER_123_1121 ();
 FILLCELL_X32 FILLER_123_1153 ();
 FILLCELL_X32 FILLER_123_1185 ();
 FILLCELL_X32 FILLER_123_1217 ();
 FILLCELL_X8 FILLER_123_1249 ();
 FILLCELL_X4 FILLER_123_1257 ();
 FILLCELL_X2 FILLER_123_1261 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X32 FILLER_123_1552 ();
 FILLCELL_X32 FILLER_123_1584 ();
 FILLCELL_X32 FILLER_123_1616 ();
 FILLCELL_X32 FILLER_123_1648 ();
 FILLCELL_X32 FILLER_123_1680 ();
 FILLCELL_X32 FILLER_123_1712 ();
 FILLCELL_X32 FILLER_123_1744 ();
 FILLCELL_X32 FILLER_123_1776 ();
 FILLCELL_X32 FILLER_123_1808 ();
 FILLCELL_X32 FILLER_123_1840 ();
 FILLCELL_X32 FILLER_123_1872 ();
 FILLCELL_X32 FILLER_123_1904 ();
 FILLCELL_X32 FILLER_123_1936 ();
 FILLCELL_X32 FILLER_123_1968 ();
 FILLCELL_X32 FILLER_123_2000 ();
 FILLCELL_X32 FILLER_123_2032 ();
 FILLCELL_X32 FILLER_123_2064 ();
 FILLCELL_X16 FILLER_123_2096 ();
 FILLCELL_X2 FILLER_123_2112 ();
 FILLCELL_X1 FILLER_123_2114 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X32 FILLER_124_1144 ();
 FILLCELL_X32 FILLER_124_1176 ();
 FILLCELL_X32 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_124_1240 ();
 FILLCELL_X32 FILLER_124_1272 ();
 FILLCELL_X32 FILLER_124_1304 ();
 FILLCELL_X32 FILLER_124_1336 ();
 FILLCELL_X32 FILLER_124_1368 ();
 FILLCELL_X32 FILLER_124_1400 ();
 FILLCELL_X32 FILLER_124_1432 ();
 FILLCELL_X32 FILLER_124_1464 ();
 FILLCELL_X32 FILLER_124_1496 ();
 FILLCELL_X32 FILLER_124_1528 ();
 FILLCELL_X32 FILLER_124_1560 ();
 FILLCELL_X32 FILLER_124_1592 ();
 FILLCELL_X32 FILLER_124_1624 ();
 FILLCELL_X32 FILLER_124_1656 ();
 FILLCELL_X32 FILLER_124_1688 ();
 FILLCELL_X32 FILLER_124_1720 ();
 FILLCELL_X32 FILLER_124_1752 ();
 FILLCELL_X32 FILLER_124_1784 ();
 FILLCELL_X32 FILLER_124_1816 ();
 FILLCELL_X32 FILLER_124_1848 ();
 FILLCELL_X8 FILLER_124_1880 ();
 FILLCELL_X4 FILLER_124_1888 ();
 FILLCELL_X2 FILLER_124_1892 ();
 FILLCELL_X32 FILLER_124_1895 ();
 FILLCELL_X32 FILLER_124_1927 ();
 FILLCELL_X32 FILLER_124_1959 ();
 FILLCELL_X32 FILLER_124_1991 ();
 FILLCELL_X32 FILLER_124_2023 ();
 FILLCELL_X32 FILLER_124_2055 ();
 FILLCELL_X16 FILLER_124_2087 ();
 FILLCELL_X8 FILLER_124_2103 ();
 FILLCELL_X4 FILLER_124_2111 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X32 FILLER_125_961 ();
 FILLCELL_X32 FILLER_125_993 ();
 FILLCELL_X32 FILLER_125_1025 ();
 FILLCELL_X32 FILLER_125_1057 ();
 FILLCELL_X32 FILLER_125_1089 ();
 FILLCELL_X32 FILLER_125_1121 ();
 FILLCELL_X32 FILLER_125_1153 ();
 FILLCELL_X32 FILLER_125_1185 ();
 FILLCELL_X32 FILLER_125_1217 ();
 FILLCELL_X8 FILLER_125_1249 ();
 FILLCELL_X4 FILLER_125_1257 ();
 FILLCELL_X2 FILLER_125_1261 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X32 FILLER_125_1648 ();
 FILLCELL_X32 FILLER_125_1680 ();
 FILLCELL_X32 FILLER_125_1712 ();
 FILLCELL_X32 FILLER_125_1744 ();
 FILLCELL_X32 FILLER_125_1776 ();
 FILLCELL_X32 FILLER_125_1808 ();
 FILLCELL_X32 FILLER_125_1840 ();
 FILLCELL_X32 FILLER_125_1872 ();
 FILLCELL_X32 FILLER_125_1904 ();
 FILLCELL_X32 FILLER_125_1936 ();
 FILLCELL_X32 FILLER_125_1968 ();
 FILLCELL_X32 FILLER_125_2000 ();
 FILLCELL_X32 FILLER_125_2032 ();
 FILLCELL_X32 FILLER_125_2064 ();
 FILLCELL_X16 FILLER_125_2096 ();
 FILLCELL_X2 FILLER_125_2112 ();
 FILLCELL_X1 FILLER_125_2114 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_126_1048 ();
 FILLCELL_X32 FILLER_126_1080 ();
 FILLCELL_X32 FILLER_126_1112 ();
 FILLCELL_X32 FILLER_126_1144 ();
 FILLCELL_X32 FILLER_126_1176 ();
 FILLCELL_X32 FILLER_126_1208 ();
 FILLCELL_X32 FILLER_126_1240 ();
 FILLCELL_X32 FILLER_126_1272 ();
 FILLCELL_X32 FILLER_126_1304 ();
 FILLCELL_X32 FILLER_126_1336 ();
 FILLCELL_X32 FILLER_126_1368 ();
 FILLCELL_X32 FILLER_126_1400 ();
 FILLCELL_X32 FILLER_126_1432 ();
 FILLCELL_X32 FILLER_126_1464 ();
 FILLCELL_X32 FILLER_126_1496 ();
 FILLCELL_X32 FILLER_126_1528 ();
 FILLCELL_X32 FILLER_126_1560 ();
 FILLCELL_X32 FILLER_126_1592 ();
 FILLCELL_X32 FILLER_126_1624 ();
 FILLCELL_X32 FILLER_126_1656 ();
 FILLCELL_X32 FILLER_126_1688 ();
 FILLCELL_X32 FILLER_126_1720 ();
 FILLCELL_X32 FILLER_126_1752 ();
 FILLCELL_X32 FILLER_126_1784 ();
 FILLCELL_X32 FILLER_126_1816 ();
 FILLCELL_X32 FILLER_126_1848 ();
 FILLCELL_X8 FILLER_126_1880 ();
 FILLCELL_X4 FILLER_126_1888 ();
 FILLCELL_X2 FILLER_126_1892 ();
 FILLCELL_X32 FILLER_126_1895 ();
 FILLCELL_X32 FILLER_126_1927 ();
 FILLCELL_X32 FILLER_126_1959 ();
 FILLCELL_X32 FILLER_126_1991 ();
 FILLCELL_X32 FILLER_126_2023 ();
 FILLCELL_X32 FILLER_126_2055 ();
 FILLCELL_X16 FILLER_126_2087 ();
 FILLCELL_X8 FILLER_126_2103 ();
 FILLCELL_X4 FILLER_126_2111 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X32 FILLER_127_1089 ();
 FILLCELL_X32 FILLER_127_1121 ();
 FILLCELL_X32 FILLER_127_1153 ();
 FILLCELL_X32 FILLER_127_1185 ();
 FILLCELL_X32 FILLER_127_1217 ();
 FILLCELL_X8 FILLER_127_1249 ();
 FILLCELL_X4 FILLER_127_1257 ();
 FILLCELL_X2 FILLER_127_1261 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X32 FILLER_127_1584 ();
 FILLCELL_X32 FILLER_127_1616 ();
 FILLCELL_X32 FILLER_127_1648 ();
 FILLCELL_X32 FILLER_127_1680 ();
 FILLCELL_X32 FILLER_127_1712 ();
 FILLCELL_X32 FILLER_127_1744 ();
 FILLCELL_X32 FILLER_127_1776 ();
 FILLCELL_X32 FILLER_127_1808 ();
 FILLCELL_X32 FILLER_127_1840 ();
 FILLCELL_X32 FILLER_127_1872 ();
 FILLCELL_X32 FILLER_127_1904 ();
 FILLCELL_X32 FILLER_127_1936 ();
 FILLCELL_X32 FILLER_127_1968 ();
 FILLCELL_X32 FILLER_127_2000 ();
 FILLCELL_X32 FILLER_127_2032 ();
 FILLCELL_X32 FILLER_127_2064 ();
 FILLCELL_X4 FILLER_127_2096 ();
 FILLCELL_X1 FILLER_127_2100 ();
 FILLCELL_X8 FILLER_127_2107 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X32 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_128_1048 ();
 FILLCELL_X32 FILLER_128_1080 ();
 FILLCELL_X32 FILLER_128_1112 ();
 FILLCELL_X32 FILLER_128_1144 ();
 FILLCELL_X32 FILLER_128_1176 ();
 FILLCELL_X32 FILLER_128_1208 ();
 FILLCELL_X32 FILLER_128_1240 ();
 FILLCELL_X32 FILLER_128_1272 ();
 FILLCELL_X32 FILLER_128_1304 ();
 FILLCELL_X32 FILLER_128_1336 ();
 FILLCELL_X32 FILLER_128_1368 ();
 FILLCELL_X32 FILLER_128_1400 ();
 FILLCELL_X32 FILLER_128_1432 ();
 FILLCELL_X32 FILLER_128_1464 ();
 FILLCELL_X32 FILLER_128_1496 ();
 FILLCELL_X32 FILLER_128_1528 ();
 FILLCELL_X32 FILLER_128_1560 ();
 FILLCELL_X32 FILLER_128_1592 ();
 FILLCELL_X32 FILLER_128_1624 ();
 FILLCELL_X32 FILLER_128_1656 ();
 FILLCELL_X32 FILLER_128_1688 ();
 FILLCELL_X32 FILLER_128_1720 ();
 FILLCELL_X32 FILLER_128_1752 ();
 FILLCELL_X32 FILLER_128_1784 ();
 FILLCELL_X32 FILLER_128_1816 ();
 FILLCELL_X32 FILLER_128_1848 ();
 FILLCELL_X8 FILLER_128_1880 ();
 FILLCELL_X4 FILLER_128_1888 ();
 FILLCELL_X2 FILLER_128_1892 ();
 FILLCELL_X32 FILLER_128_1895 ();
 FILLCELL_X32 FILLER_128_1927 ();
 FILLCELL_X32 FILLER_128_1959 ();
 FILLCELL_X32 FILLER_128_1991 ();
 FILLCELL_X32 FILLER_128_2023 ();
 FILLCELL_X16 FILLER_128_2055 ();
 FILLCELL_X8 FILLER_128_2071 ();
 FILLCELL_X4 FILLER_128_2079 ();
 FILLCELL_X4 FILLER_128_2096 ();
 FILLCELL_X2 FILLER_128_2100 ();
 FILLCELL_X1 FILLER_128_2102 ();
 FILLCELL_X1 FILLER_128_2106 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_993 ();
 FILLCELL_X32 FILLER_129_1025 ();
 FILLCELL_X32 FILLER_129_1057 ();
 FILLCELL_X32 FILLER_129_1089 ();
 FILLCELL_X32 FILLER_129_1121 ();
 FILLCELL_X32 FILLER_129_1153 ();
 FILLCELL_X32 FILLER_129_1185 ();
 FILLCELL_X32 FILLER_129_1217 ();
 FILLCELL_X8 FILLER_129_1249 ();
 FILLCELL_X4 FILLER_129_1257 ();
 FILLCELL_X2 FILLER_129_1261 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X32 FILLER_129_1584 ();
 FILLCELL_X32 FILLER_129_1616 ();
 FILLCELL_X32 FILLER_129_1648 ();
 FILLCELL_X32 FILLER_129_1680 ();
 FILLCELL_X32 FILLER_129_1712 ();
 FILLCELL_X32 FILLER_129_1744 ();
 FILLCELL_X32 FILLER_129_1776 ();
 FILLCELL_X32 FILLER_129_1808 ();
 FILLCELL_X32 FILLER_129_1840 ();
 FILLCELL_X32 FILLER_129_1872 ();
 FILLCELL_X32 FILLER_129_1904 ();
 FILLCELL_X32 FILLER_129_1936 ();
 FILLCELL_X32 FILLER_129_1968 ();
 FILLCELL_X32 FILLER_129_2000 ();
 FILLCELL_X32 FILLER_129_2032 ();
 FILLCELL_X32 FILLER_129_2064 ();
 FILLCELL_X1 FILLER_129_2096 ();
 FILLCELL_X8 FILLER_129_2103 ();
 FILLCELL_X4 FILLER_129_2111 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X32 FILLER_130_1016 ();
 FILLCELL_X32 FILLER_130_1048 ();
 FILLCELL_X32 FILLER_130_1080 ();
 FILLCELL_X32 FILLER_130_1112 ();
 FILLCELL_X32 FILLER_130_1144 ();
 FILLCELL_X32 FILLER_130_1176 ();
 FILLCELL_X32 FILLER_130_1208 ();
 FILLCELL_X32 FILLER_130_1240 ();
 FILLCELL_X32 FILLER_130_1272 ();
 FILLCELL_X32 FILLER_130_1304 ();
 FILLCELL_X32 FILLER_130_1336 ();
 FILLCELL_X32 FILLER_130_1368 ();
 FILLCELL_X32 FILLER_130_1400 ();
 FILLCELL_X32 FILLER_130_1432 ();
 FILLCELL_X32 FILLER_130_1464 ();
 FILLCELL_X32 FILLER_130_1496 ();
 FILLCELL_X32 FILLER_130_1528 ();
 FILLCELL_X32 FILLER_130_1560 ();
 FILLCELL_X32 FILLER_130_1592 ();
 FILLCELL_X32 FILLER_130_1624 ();
 FILLCELL_X32 FILLER_130_1656 ();
 FILLCELL_X32 FILLER_130_1688 ();
 FILLCELL_X32 FILLER_130_1720 ();
 FILLCELL_X32 FILLER_130_1752 ();
 FILLCELL_X32 FILLER_130_1784 ();
 FILLCELL_X32 FILLER_130_1816 ();
 FILLCELL_X32 FILLER_130_1848 ();
 FILLCELL_X8 FILLER_130_1880 ();
 FILLCELL_X4 FILLER_130_1888 ();
 FILLCELL_X2 FILLER_130_1892 ();
 FILLCELL_X32 FILLER_130_1895 ();
 FILLCELL_X32 FILLER_130_1927 ();
 FILLCELL_X32 FILLER_130_1959 ();
 FILLCELL_X32 FILLER_130_1991 ();
 FILLCELL_X32 FILLER_130_2023 ();
 FILLCELL_X32 FILLER_130_2055 ();
 FILLCELL_X16 FILLER_130_2087 ();
 FILLCELL_X8 FILLER_130_2103 ();
 FILLCELL_X4 FILLER_130_2111 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X32 FILLER_131_993 ();
 FILLCELL_X32 FILLER_131_1025 ();
 FILLCELL_X32 FILLER_131_1057 ();
 FILLCELL_X32 FILLER_131_1089 ();
 FILLCELL_X32 FILLER_131_1121 ();
 FILLCELL_X32 FILLER_131_1153 ();
 FILLCELL_X32 FILLER_131_1185 ();
 FILLCELL_X32 FILLER_131_1217 ();
 FILLCELL_X8 FILLER_131_1249 ();
 FILLCELL_X4 FILLER_131_1257 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X32 FILLER_131_1584 ();
 FILLCELL_X32 FILLER_131_1616 ();
 FILLCELL_X32 FILLER_131_1648 ();
 FILLCELL_X32 FILLER_131_1680 ();
 FILLCELL_X32 FILLER_131_1712 ();
 FILLCELL_X32 FILLER_131_1744 ();
 FILLCELL_X32 FILLER_131_1776 ();
 FILLCELL_X32 FILLER_131_1808 ();
 FILLCELL_X32 FILLER_131_1840 ();
 FILLCELL_X32 FILLER_131_1872 ();
 FILLCELL_X32 FILLER_131_1904 ();
 FILLCELL_X32 FILLER_131_1936 ();
 FILLCELL_X32 FILLER_131_1968 ();
 FILLCELL_X32 FILLER_131_2000 ();
 FILLCELL_X32 FILLER_131_2032 ();
 FILLCELL_X32 FILLER_131_2064 ();
 FILLCELL_X16 FILLER_131_2096 ();
 FILLCELL_X2 FILLER_131_2112 ();
 FILLCELL_X1 FILLER_131_2114 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X32 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_132_1048 ();
 FILLCELL_X32 FILLER_132_1080 ();
 FILLCELL_X32 FILLER_132_1112 ();
 FILLCELL_X32 FILLER_132_1144 ();
 FILLCELL_X32 FILLER_132_1176 ();
 FILLCELL_X32 FILLER_132_1208 ();
 FILLCELL_X32 FILLER_132_1240 ();
 FILLCELL_X32 FILLER_132_1272 ();
 FILLCELL_X32 FILLER_132_1304 ();
 FILLCELL_X32 FILLER_132_1336 ();
 FILLCELL_X32 FILLER_132_1368 ();
 FILLCELL_X32 FILLER_132_1400 ();
 FILLCELL_X32 FILLER_132_1432 ();
 FILLCELL_X32 FILLER_132_1464 ();
 FILLCELL_X32 FILLER_132_1496 ();
 FILLCELL_X32 FILLER_132_1528 ();
 FILLCELL_X32 FILLER_132_1560 ();
 FILLCELL_X32 FILLER_132_1592 ();
 FILLCELL_X32 FILLER_132_1624 ();
 FILLCELL_X32 FILLER_132_1656 ();
 FILLCELL_X32 FILLER_132_1688 ();
 FILLCELL_X32 FILLER_132_1720 ();
 FILLCELL_X32 FILLER_132_1752 ();
 FILLCELL_X32 FILLER_132_1784 ();
 FILLCELL_X32 FILLER_132_1816 ();
 FILLCELL_X32 FILLER_132_1848 ();
 FILLCELL_X8 FILLER_132_1880 ();
 FILLCELL_X4 FILLER_132_1888 ();
 FILLCELL_X2 FILLER_132_1892 ();
 FILLCELL_X32 FILLER_132_1895 ();
 FILLCELL_X32 FILLER_132_1927 ();
 FILLCELL_X32 FILLER_132_1959 ();
 FILLCELL_X32 FILLER_132_1991 ();
 FILLCELL_X32 FILLER_132_2023 ();
 FILLCELL_X32 FILLER_132_2055 ();
 FILLCELL_X16 FILLER_132_2087 ();
 FILLCELL_X8 FILLER_132_2103 ();
 FILLCELL_X4 FILLER_132_2111 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X32 FILLER_133_993 ();
 FILLCELL_X32 FILLER_133_1025 ();
 FILLCELL_X32 FILLER_133_1057 ();
 FILLCELL_X32 FILLER_133_1089 ();
 FILLCELL_X32 FILLER_133_1121 ();
 FILLCELL_X32 FILLER_133_1153 ();
 FILLCELL_X32 FILLER_133_1185 ();
 FILLCELL_X32 FILLER_133_1217 ();
 FILLCELL_X8 FILLER_133_1249 ();
 FILLCELL_X4 FILLER_133_1257 ();
 FILLCELL_X2 FILLER_133_1261 ();
 FILLCELL_X16 FILLER_133_1264 ();
 FILLCELL_X4 FILLER_133_1280 ();
 FILLCELL_X2 FILLER_133_1284 ();
 FILLCELL_X1 FILLER_133_1286 ();
 FILLCELL_X32 FILLER_133_1290 ();
 FILLCELL_X32 FILLER_133_1322 ();
 FILLCELL_X32 FILLER_133_1354 ();
 FILLCELL_X32 FILLER_133_1386 ();
 FILLCELL_X32 FILLER_133_1418 ();
 FILLCELL_X32 FILLER_133_1450 ();
 FILLCELL_X32 FILLER_133_1482 ();
 FILLCELL_X32 FILLER_133_1514 ();
 FILLCELL_X32 FILLER_133_1546 ();
 FILLCELL_X32 FILLER_133_1578 ();
 FILLCELL_X32 FILLER_133_1610 ();
 FILLCELL_X32 FILLER_133_1642 ();
 FILLCELL_X32 FILLER_133_1674 ();
 FILLCELL_X32 FILLER_133_1706 ();
 FILLCELL_X32 FILLER_133_1738 ();
 FILLCELL_X32 FILLER_133_1770 ();
 FILLCELL_X32 FILLER_133_1802 ();
 FILLCELL_X32 FILLER_133_1834 ();
 FILLCELL_X32 FILLER_133_1866 ();
 FILLCELL_X32 FILLER_133_1898 ();
 FILLCELL_X32 FILLER_133_1930 ();
 FILLCELL_X32 FILLER_133_1962 ();
 FILLCELL_X32 FILLER_133_1994 ();
 FILLCELL_X32 FILLER_133_2026 ();
 FILLCELL_X32 FILLER_133_2058 ();
 FILLCELL_X4 FILLER_133_2090 ();
 FILLCELL_X2 FILLER_133_2094 ();
 FILLCELL_X4 FILLER_133_2100 ();
 FILLCELL_X4 FILLER_133_2106 ();
 FILLCELL_X2 FILLER_133_2110 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X8 FILLER_134_984 ();
 FILLCELL_X32 FILLER_134_996 ();
 FILLCELL_X32 FILLER_134_1028 ();
 FILLCELL_X32 FILLER_134_1060 ();
 FILLCELL_X32 FILLER_134_1092 ();
 FILLCELL_X32 FILLER_134_1124 ();
 FILLCELL_X32 FILLER_134_1156 ();
 FILLCELL_X32 FILLER_134_1188 ();
 FILLCELL_X32 FILLER_134_1220 ();
 FILLCELL_X16 FILLER_134_1252 ();
 FILLCELL_X8 FILLER_134_1268 ();
 FILLCELL_X4 FILLER_134_1276 ();
 FILLCELL_X2 FILLER_134_1280 ();
 FILLCELL_X8 FILLER_134_1292 ();
 FILLCELL_X4 FILLER_134_1300 ();
 FILLCELL_X16 FILLER_134_1309 ();
 FILLCELL_X4 FILLER_134_1325 ();
 FILLCELL_X32 FILLER_134_1332 ();
 FILLCELL_X32 FILLER_134_1364 ();
 FILLCELL_X32 FILLER_134_1396 ();
 FILLCELL_X32 FILLER_134_1428 ();
 FILLCELL_X32 FILLER_134_1460 ();
 FILLCELL_X32 FILLER_134_1492 ();
 FILLCELL_X32 FILLER_134_1524 ();
 FILLCELL_X32 FILLER_134_1556 ();
 FILLCELL_X32 FILLER_134_1588 ();
 FILLCELL_X32 FILLER_134_1620 ();
 FILLCELL_X32 FILLER_134_1652 ();
 FILLCELL_X32 FILLER_134_1684 ();
 FILLCELL_X32 FILLER_134_1716 ();
 FILLCELL_X32 FILLER_134_1748 ();
 FILLCELL_X32 FILLER_134_1780 ();
 FILLCELL_X32 FILLER_134_1812 ();
 FILLCELL_X32 FILLER_134_1844 ();
 FILLCELL_X16 FILLER_134_1876 ();
 FILLCELL_X2 FILLER_134_1892 ();
 FILLCELL_X32 FILLER_134_1895 ();
 FILLCELL_X32 FILLER_134_1927 ();
 FILLCELL_X32 FILLER_134_1959 ();
 FILLCELL_X32 FILLER_134_1991 ();
 FILLCELL_X32 FILLER_134_2023 ();
 FILLCELL_X32 FILLER_134_2055 ();
 FILLCELL_X16 FILLER_134_2087 ();
 FILLCELL_X8 FILLER_134_2103 ();
 FILLCELL_X4 FILLER_134_2111 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X16 FILLER_135_929 ();
 FILLCELL_X2 FILLER_135_945 ();
 FILLCELL_X32 FILLER_135_951 ();
 FILLCELL_X32 FILLER_135_983 ();
 FILLCELL_X32 FILLER_135_1015 ();
 FILLCELL_X4 FILLER_135_1047 ();
 FILLCELL_X1 FILLER_135_1051 ();
 FILLCELL_X16 FILLER_135_1059 ();
 FILLCELL_X8 FILLER_135_1075 ();
 FILLCELL_X4 FILLER_135_1083 ();
 FILLCELL_X16 FILLER_135_1094 ();
 FILLCELL_X4 FILLER_135_1110 ();
 FILLCELL_X2 FILLER_135_1114 ();
 FILLCELL_X16 FILLER_135_1140 ();
 FILLCELL_X2 FILLER_135_1156 ();
 FILLCELL_X1 FILLER_135_1158 ();
 FILLCELL_X16 FILLER_135_1167 ();
 FILLCELL_X2 FILLER_135_1183 ();
 FILLCELL_X4 FILLER_135_1198 ();
 FILLCELL_X2 FILLER_135_1202 ();
 FILLCELL_X1 FILLER_135_1204 ();
 FILLCELL_X32 FILLER_135_1227 ();
 FILLCELL_X4 FILLER_135_1259 ();
 FILLCELL_X16 FILLER_135_1264 ();
 FILLCELL_X2 FILLER_135_1280 ();
 FILLCELL_X1 FILLER_135_1282 ();
 FILLCELL_X32 FILLER_135_1309 ();
 FILLCELL_X32 FILLER_135_1341 ();
 FILLCELL_X32 FILLER_135_1373 ();
 FILLCELL_X32 FILLER_135_1405 ();
 FILLCELL_X32 FILLER_135_1437 ();
 FILLCELL_X32 FILLER_135_1469 ();
 FILLCELL_X32 FILLER_135_1501 ();
 FILLCELL_X32 FILLER_135_1533 ();
 FILLCELL_X32 FILLER_135_1565 ();
 FILLCELL_X32 FILLER_135_1597 ();
 FILLCELL_X32 FILLER_135_1629 ();
 FILLCELL_X32 FILLER_135_1661 ();
 FILLCELL_X32 FILLER_135_1693 ();
 FILLCELL_X32 FILLER_135_1725 ();
 FILLCELL_X32 FILLER_135_1757 ();
 FILLCELL_X32 FILLER_135_1789 ();
 FILLCELL_X32 FILLER_135_1821 ();
 FILLCELL_X32 FILLER_135_1853 ();
 FILLCELL_X32 FILLER_135_1885 ();
 FILLCELL_X32 FILLER_135_1917 ();
 FILLCELL_X32 FILLER_135_1949 ();
 FILLCELL_X32 FILLER_135_1981 ();
 FILLCELL_X32 FILLER_135_2013 ();
 FILLCELL_X32 FILLER_135_2045 ();
 FILLCELL_X32 FILLER_135_2077 ();
 FILLCELL_X4 FILLER_135_2109 ();
 FILLCELL_X2 FILLER_135_2113 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X16 FILLER_136_1016 ();
 FILLCELL_X8 FILLER_136_1066 ();
 FILLCELL_X4 FILLER_136_1074 ();
 FILLCELL_X1 FILLER_136_1078 ();
 FILLCELL_X2 FILLER_136_1086 ();
 FILLCELL_X8 FILLER_136_1105 ();
 FILLCELL_X2 FILLER_136_1113 ();
 FILLCELL_X1 FILLER_136_1115 ();
 FILLCELL_X16 FILLER_136_1123 ();
 FILLCELL_X4 FILLER_136_1139 ();
 FILLCELL_X2 FILLER_136_1143 ();
 FILLCELL_X16 FILLER_136_1175 ();
 FILLCELL_X8 FILLER_136_1191 ();
 FILLCELL_X16 FILLER_136_1206 ();
 FILLCELL_X1 FILLER_136_1222 ();
 FILLCELL_X4 FILLER_136_1235 ();
 FILLCELL_X1 FILLER_136_1239 ();
 FILLCELL_X8 FILLER_136_1262 ();
 FILLCELL_X2 FILLER_136_1270 ();
 FILLCELL_X1 FILLER_136_1288 ();
 FILLCELL_X32 FILLER_136_1291 ();
 FILLCELL_X32 FILLER_136_1323 ();
 FILLCELL_X32 FILLER_136_1355 ();
 FILLCELL_X32 FILLER_136_1387 ();
 FILLCELL_X32 FILLER_136_1419 ();
 FILLCELL_X32 FILLER_136_1451 ();
 FILLCELL_X32 FILLER_136_1483 ();
 FILLCELL_X32 FILLER_136_1515 ();
 FILLCELL_X32 FILLER_136_1547 ();
 FILLCELL_X32 FILLER_136_1579 ();
 FILLCELL_X32 FILLER_136_1611 ();
 FILLCELL_X32 FILLER_136_1643 ();
 FILLCELL_X32 FILLER_136_1675 ();
 FILLCELL_X32 FILLER_136_1707 ();
 FILLCELL_X32 FILLER_136_1739 ();
 FILLCELL_X32 FILLER_136_1771 ();
 FILLCELL_X32 FILLER_136_1803 ();
 FILLCELL_X32 FILLER_136_1835 ();
 FILLCELL_X16 FILLER_136_1867 ();
 FILLCELL_X8 FILLER_136_1883 ();
 FILLCELL_X2 FILLER_136_1891 ();
 FILLCELL_X1 FILLER_136_1893 ();
 FILLCELL_X32 FILLER_136_1895 ();
 FILLCELL_X32 FILLER_136_1927 ();
 FILLCELL_X32 FILLER_136_1959 ();
 FILLCELL_X32 FILLER_136_1991 ();
 FILLCELL_X32 FILLER_136_2023 ();
 FILLCELL_X32 FILLER_136_2055 ();
 FILLCELL_X16 FILLER_136_2087 ();
 FILLCELL_X8 FILLER_136_2103 ();
 FILLCELL_X4 FILLER_136_2111 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X32 FILLER_137_801 ();
 FILLCELL_X32 FILLER_137_833 ();
 FILLCELL_X32 FILLER_137_865 ();
 FILLCELL_X32 FILLER_137_897 ();
 FILLCELL_X32 FILLER_137_929 ();
 FILLCELL_X16 FILLER_137_961 ();
 FILLCELL_X8 FILLER_137_977 ();
 FILLCELL_X4 FILLER_137_985 ();
 FILLCELL_X8 FILLER_137_996 ();
 FILLCELL_X4 FILLER_137_1004 ();
 FILLCELL_X2 FILLER_137_1008 ();
 FILLCELL_X8 FILLER_137_1027 ();
 FILLCELL_X4 FILLER_137_1035 ();
 FILLCELL_X2 FILLER_137_1039 ();
 FILLCELL_X1 FILLER_137_1041 ();
 FILLCELL_X4 FILLER_137_1049 ();
 FILLCELL_X1 FILLER_137_1053 ();
 FILLCELL_X8 FILLER_137_1061 ();
 FILLCELL_X4 FILLER_137_1069 ();
 FILLCELL_X1 FILLER_137_1073 ();
 FILLCELL_X2 FILLER_137_1091 ();
 FILLCELL_X8 FILLER_137_1100 ();
 FILLCELL_X2 FILLER_137_1108 ();
 FILLCELL_X1 FILLER_137_1110 ();
 FILLCELL_X1 FILLER_137_1128 ();
 FILLCELL_X8 FILLER_137_1136 ();
 FILLCELL_X4 FILLER_137_1144 ();
 FILLCELL_X2 FILLER_137_1148 ();
 FILLCELL_X1 FILLER_137_1157 ();
 FILLCELL_X32 FILLER_137_1176 ();
 FILLCELL_X8 FILLER_137_1208 ();
 FILLCELL_X4 FILLER_137_1216 ();
 FILLCELL_X2 FILLER_137_1220 ();
 FILLCELL_X1 FILLER_137_1222 ();
 FILLCELL_X16 FILLER_137_1240 ();
 FILLCELL_X4 FILLER_137_1256 ();
 FILLCELL_X2 FILLER_137_1260 ();
 FILLCELL_X1 FILLER_137_1262 ();
 FILLCELL_X8 FILLER_137_1264 ();
 FILLCELL_X1 FILLER_137_1272 ();
 FILLCELL_X32 FILLER_137_1275 ();
 FILLCELL_X32 FILLER_137_1307 ();
 FILLCELL_X32 FILLER_137_1339 ();
 FILLCELL_X32 FILLER_137_1371 ();
 FILLCELL_X32 FILLER_137_1403 ();
 FILLCELL_X32 FILLER_137_1435 ();
 FILLCELL_X32 FILLER_137_1467 ();
 FILLCELL_X32 FILLER_137_1499 ();
 FILLCELL_X32 FILLER_137_1531 ();
 FILLCELL_X32 FILLER_137_1563 ();
 FILLCELL_X32 FILLER_137_1595 ();
 FILLCELL_X32 FILLER_137_1627 ();
 FILLCELL_X32 FILLER_137_1659 ();
 FILLCELL_X32 FILLER_137_1691 ();
 FILLCELL_X32 FILLER_137_1723 ();
 FILLCELL_X32 FILLER_137_1755 ();
 FILLCELL_X32 FILLER_137_1787 ();
 FILLCELL_X32 FILLER_137_1819 ();
 FILLCELL_X32 FILLER_137_1851 ();
 FILLCELL_X32 FILLER_137_1883 ();
 FILLCELL_X32 FILLER_137_1915 ();
 FILLCELL_X32 FILLER_137_1947 ();
 FILLCELL_X32 FILLER_137_1979 ();
 FILLCELL_X32 FILLER_137_2011 ();
 FILLCELL_X32 FILLER_137_2043 ();
 FILLCELL_X32 FILLER_137_2075 ();
 FILLCELL_X8 FILLER_137_2107 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X16 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X32 FILLER_138_824 ();
 FILLCELL_X32 FILLER_138_856 ();
 FILLCELL_X32 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_920 ();
 FILLCELL_X32 FILLER_138_952 ();
 FILLCELL_X1 FILLER_138_984 ();
 FILLCELL_X8 FILLER_138_1002 ();
 FILLCELL_X2 FILLER_138_1010 ();
 FILLCELL_X32 FILLER_138_1026 ();
 FILLCELL_X32 FILLER_138_1058 ();
 FILLCELL_X32 FILLER_138_1090 ();
 FILLCELL_X32 FILLER_138_1122 ();
 FILLCELL_X2 FILLER_138_1154 ();
 FILLCELL_X16 FILLER_138_1161 ();
 FILLCELL_X8 FILLER_138_1177 ();
 FILLCELL_X4 FILLER_138_1185 ();
 FILLCELL_X2 FILLER_138_1214 ();
 FILLCELL_X1 FILLER_138_1216 ();
 FILLCELL_X32 FILLER_138_1227 ();
 FILLCELL_X8 FILLER_138_1259 ();
 FILLCELL_X4 FILLER_138_1267 ();
 FILLCELL_X1 FILLER_138_1271 ();
 FILLCELL_X2 FILLER_138_1282 ();
 FILLCELL_X32 FILLER_138_1301 ();
 FILLCELL_X32 FILLER_138_1333 ();
 FILLCELL_X32 FILLER_138_1365 ();
 FILLCELL_X32 FILLER_138_1397 ();
 FILLCELL_X32 FILLER_138_1429 ();
 FILLCELL_X32 FILLER_138_1461 ();
 FILLCELL_X32 FILLER_138_1493 ();
 FILLCELL_X32 FILLER_138_1525 ();
 FILLCELL_X32 FILLER_138_1557 ();
 FILLCELL_X32 FILLER_138_1589 ();
 FILLCELL_X32 FILLER_138_1621 ();
 FILLCELL_X32 FILLER_138_1653 ();
 FILLCELL_X32 FILLER_138_1685 ();
 FILLCELL_X32 FILLER_138_1717 ();
 FILLCELL_X32 FILLER_138_1749 ();
 FILLCELL_X32 FILLER_138_1781 ();
 FILLCELL_X32 FILLER_138_1813 ();
 FILLCELL_X32 FILLER_138_1845 ();
 FILLCELL_X16 FILLER_138_1877 ();
 FILLCELL_X1 FILLER_138_1893 ();
 FILLCELL_X32 FILLER_138_1895 ();
 FILLCELL_X32 FILLER_138_1927 ();
 FILLCELL_X32 FILLER_138_1959 ();
 FILLCELL_X32 FILLER_138_1991 ();
 FILLCELL_X32 FILLER_138_2023 ();
 FILLCELL_X32 FILLER_138_2055 ();
 FILLCELL_X16 FILLER_138_2087 ();
 FILLCELL_X8 FILLER_138_2103 ();
 FILLCELL_X4 FILLER_138_2111 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X32 FILLER_139_577 ();
 FILLCELL_X32 FILLER_139_609 ();
 FILLCELL_X32 FILLER_139_641 ();
 FILLCELL_X32 FILLER_139_673 ();
 FILLCELL_X32 FILLER_139_705 ();
 FILLCELL_X32 FILLER_139_737 ();
 FILLCELL_X32 FILLER_139_769 ();
 FILLCELL_X32 FILLER_139_801 ();
 FILLCELL_X32 FILLER_139_833 ();
 FILLCELL_X32 FILLER_139_865 ();
 FILLCELL_X32 FILLER_139_897 ();
 FILLCELL_X32 FILLER_139_929 ();
 FILLCELL_X32 FILLER_139_961 ();
 FILLCELL_X32 FILLER_139_993 ();
 FILLCELL_X32 FILLER_139_1025 ();
 FILLCELL_X16 FILLER_139_1057 ();
 FILLCELL_X8 FILLER_139_1073 ();
 FILLCELL_X32 FILLER_139_1088 ();
 FILLCELL_X32 FILLER_139_1120 ();
 FILLCELL_X4 FILLER_139_1152 ();
 FILLCELL_X2 FILLER_139_1156 ();
 FILLCELL_X1 FILLER_139_1158 ();
 FILLCELL_X16 FILLER_139_1161 ();
 FILLCELL_X8 FILLER_139_1177 ();
 FILLCELL_X4 FILLER_139_1185 ();
 FILLCELL_X1 FILLER_139_1189 ();
 FILLCELL_X16 FILLER_139_1197 ();
 FILLCELL_X8 FILLER_139_1213 ();
 FILLCELL_X2 FILLER_139_1221 ();
 FILLCELL_X32 FILLER_139_1229 ();
 FILLCELL_X2 FILLER_139_1261 ();
 FILLCELL_X16 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1289 ();
 FILLCELL_X32 FILLER_139_1321 ();
 FILLCELL_X32 FILLER_139_1353 ();
 FILLCELL_X32 FILLER_139_1385 ();
 FILLCELL_X32 FILLER_139_1417 ();
 FILLCELL_X32 FILLER_139_1449 ();
 FILLCELL_X32 FILLER_139_1481 ();
 FILLCELL_X32 FILLER_139_1513 ();
 FILLCELL_X32 FILLER_139_1545 ();
 FILLCELL_X32 FILLER_139_1577 ();
 FILLCELL_X32 FILLER_139_1609 ();
 FILLCELL_X32 FILLER_139_1641 ();
 FILLCELL_X32 FILLER_139_1673 ();
 FILLCELL_X32 FILLER_139_1705 ();
 FILLCELL_X32 FILLER_139_1737 ();
 FILLCELL_X32 FILLER_139_1769 ();
 FILLCELL_X32 FILLER_139_1801 ();
 FILLCELL_X32 FILLER_139_1833 ();
 FILLCELL_X32 FILLER_139_1865 ();
 FILLCELL_X32 FILLER_139_1897 ();
 FILLCELL_X32 FILLER_139_1929 ();
 FILLCELL_X32 FILLER_139_1961 ();
 FILLCELL_X32 FILLER_139_1993 ();
 FILLCELL_X32 FILLER_139_2025 ();
 FILLCELL_X32 FILLER_139_2057 ();
 FILLCELL_X16 FILLER_139_2089 ();
 FILLCELL_X8 FILLER_139_2105 ();
 FILLCELL_X2 FILLER_139_2113 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X4 FILLER_140_1048 ();
 FILLCELL_X1 FILLER_140_1052 ();
 FILLCELL_X16 FILLER_140_1060 ();
 FILLCELL_X16 FILLER_140_1093 ();
 FILLCELL_X8 FILLER_140_1109 ();
 FILLCELL_X4 FILLER_140_1117 ();
 FILLCELL_X2 FILLER_140_1121 ();
 FILLCELL_X1 FILLER_140_1123 ();
 FILLCELL_X16 FILLER_140_1131 ();
 FILLCELL_X8 FILLER_140_1147 ();
 FILLCELL_X1 FILLER_140_1155 ();
 FILLCELL_X4 FILLER_140_1174 ();
 FILLCELL_X2 FILLER_140_1178 ();
 FILLCELL_X32 FILLER_140_1184 ();
 FILLCELL_X4 FILLER_140_1216 ();
 FILLCELL_X1 FILLER_140_1220 ();
 FILLCELL_X1 FILLER_140_1227 ();
 FILLCELL_X4 FILLER_140_1235 ();
 FILLCELL_X2 FILLER_140_1239 ();
 FILLCELL_X1 FILLER_140_1241 ();
 FILLCELL_X8 FILLER_140_1264 ();
 FILLCELL_X4 FILLER_140_1272 ();
 FILLCELL_X2 FILLER_140_1276 ();
 FILLCELL_X32 FILLER_140_1288 ();
 FILLCELL_X32 FILLER_140_1320 ();
 FILLCELL_X32 FILLER_140_1352 ();
 FILLCELL_X32 FILLER_140_1384 ();
 FILLCELL_X32 FILLER_140_1416 ();
 FILLCELL_X32 FILLER_140_1448 ();
 FILLCELL_X32 FILLER_140_1480 ();
 FILLCELL_X32 FILLER_140_1512 ();
 FILLCELL_X32 FILLER_140_1544 ();
 FILLCELL_X32 FILLER_140_1576 ();
 FILLCELL_X32 FILLER_140_1608 ();
 FILLCELL_X32 FILLER_140_1640 ();
 FILLCELL_X32 FILLER_140_1672 ();
 FILLCELL_X32 FILLER_140_1704 ();
 FILLCELL_X32 FILLER_140_1736 ();
 FILLCELL_X32 FILLER_140_1768 ();
 FILLCELL_X32 FILLER_140_1800 ();
 FILLCELL_X32 FILLER_140_1832 ();
 FILLCELL_X16 FILLER_140_1864 ();
 FILLCELL_X8 FILLER_140_1880 ();
 FILLCELL_X4 FILLER_140_1888 ();
 FILLCELL_X2 FILLER_140_1892 ();
 FILLCELL_X32 FILLER_140_1895 ();
 FILLCELL_X32 FILLER_140_1927 ();
 FILLCELL_X32 FILLER_140_1959 ();
 FILLCELL_X32 FILLER_140_1991 ();
 FILLCELL_X32 FILLER_140_2023 ();
 FILLCELL_X32 FILLER_140_2055 ();
 FILLCELL_X8 FILLER_140_2087 ();
 FILLCELL_X16 FILLER_140_2098 ();
 FILLCELL_X1 FILLER_140_2114 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X8 FILLER_141_993 ();
 FILLCELL_X1 FILLER_141_1001 ();
 FILLCELL_X4 FILLER_141_1026 ();
 FILLCELL_X2 FILLER_141_1030 ();
 FILLCELL_X8 FILLER_141_1073 ();
 FILLCELL_X4 FILLER_141_1081 ();
 FILLCELL_X2 FILLER_141_1085 ();
 FILLCELL_X1 FILLER_141_1087 ();
 FILLCELL_X16 FILLER_141_1095 ();
 FILLCELL_X2 FILLER_141_1111 ();
 FILLCELL_X1 FILLER_141_1113 ();
 FILLCELL_X1 FILLER_141_1155 ();
 FILLCELL_X2 FILLER_141_1174 ();
 FILLCELL_X1 FILLER_141_1176 ();
 FILLCELL_X16 FILLER_141_1200 ();
 FILLCELL_X8 FILLER_141_1216 ();
 FILLCELL_X4 FILLER_141_1224 ();
 FILLCELL_X16 FILLER_141_1235 ();
 FILLCELL_X8 FILLER_141_1251 ();
 FILLCELL_X4 FILLER_141_1259 ();
 FILLCELL_X8 FILLER_141_1264 ();
 FILLCELL_X4 FILLER_141_1272 ();
 FILLCELL_X1 FILLER_141_1276 ();
 FILLCELL_X32 FILLER_141_1297 ();
 FILLCELL_X32 FILLER_141_1329 ();
 FILLCELL_X32 FILLER_141_1361 ();
 FILLCELL_X32 FILLER_141_1393 ();
 FILLCELL_X32 FILLER_141_1425 ();
 FILLCELL_X32 FILLER_141_1457 ();
 FILLCELL_X32 FILLER_141_1489 ();
 FILLCELL_X32 FILLER_141_1521 ();
 FILLCELL_X32 FILLER_141_1553 ();
 FILLCELL_X32 FILLER_141_1585 ();
 FILLCELL_X32 FILLER_141_1617 ();
 FILLCELL_X32 FILLER_141_1649 ();
 FILLCELL_X32 FILLER_141_1681 ();
 FILLCELL_X32 FILLER_141_1713 ();
 FILLCELL_X32 FILLER_141_1745 ();
 FILLCELL_X32 FILLER_141_1777 ();
 FILLCELL_X32 FILLER_141_1809 ();
 FILLCELL_X32 FILLER_141_1841 ();
 FILLCELL_X32 FILLER_141_1873 ();
 FILLCELL_X32 FILLER_141_1905 ();
 FILLCELL_X32 FILLER_141_1937 ();
 FILLCELL_X32 FILLER_141_1969 ();
 FILLCELL_X32 FILLER_141_2001 ();
 FILLCELL_X32 FILLER_141_2033 ();
 FILLCELL_X32 FILLER_141_2065 ();
 FILLCELL_X16 FILLER_141_2097 ();
 FILLCELL_X2 FILLER_141_2113 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X16 FILLER_142_952 ();
 FILLCELL_X8 FILLER_142_968 ();
 FILLCELL_X2 FILLER_142_976 ();
 FILLCELL_X1 FILLER_142_978 ();
 FILLCELL_X8 FILLER_142_1003 ();
 FILLCELL_X4 FILLER_142_1011 ();
 FILLCELL_X1 FILLER_142_1015 ();
 FILLCELL_X2 FILLER_142_1023 ();
 FILLCELL_X1 FILLER_142_1025 ();
 FILLCELL_X16 FILLER_142_1031 ();
 FILLCELL_X4 FILLER_142_1047 ();
 FILLCELL_X1 FILLER_142_1058 ();
 FILLCELL_X16 FILLER_142_1068 ();
 FILLCELL_X2 FILLER_142_1084 ();
 FILLCELL_X1 FILLER_142_1086 ();
 FILLCELL_X16 FILLER_142_1104 ();
 FILLCELL_X8 FILLER_142_1120 ();
 FILLCELL_X4 FILLER_142_1128 ();
 FILLCELL_X1 FILLER_142_1132 ();
 FILLCELL_X32 FILLER_142_1140 ();
 FILLCELL_X16 FILLER_142_1172 ();
 FILLCELL_X8 FILLER_142_1188 ();
 FILLCELL_X2 FILLER_142_1196 ();
 FILLCELL_X1 FILLER_142_1198 ();
 FILLCELL_X16 FILLER_142_1206 ();
 FILLCELL_X8 FILLER_142_1222 ();
 FILLCELL_X4 FILLER_142_1230 ();
 FILLCELL_X2 FILLER_142_1234 ();
 FILLCELL_X1 FILLER_142_1236 ();
 FILLCELL_X4 FILLER_142_1257 ();
 FILLCELL_X2 FILLER_142_1261 ();
 FILLCELL_X4 FILLER_142_1272 ();
 FILLCELL_X1 FILLER_142_1276 ();
 FILLCELL_X32 FILLER_142_1295 ();
 FILLCELL_X32 FILLER_142_1327 ();
 FILLCELL_X32 FILLER_142_1359 ();
 FILLCELL_X32 FILLER_142_1391 ();
 FILLCELL_X32 FILLER_142_1423 ();
 FILLCELL_X32 FILLER_142_1455 ();
 FILLCELL_X32 FILLER_142_1487 ();
 FILLCELL_X32 FILLER_142_1519 ();
 FILLCELL_X32 FILLER_142_1551 ();
 FILLCELL_X32 FILLER_142_1583 ();
 FILLCELL_X32 FILLER_142_1615 ();
 FILLCELL_X32 FILLER_142_1647 ();
 FILLCELL_X32 FILLER_142_1679 ();
 FILLCELL_X32 FILLER_142_1711 ();
 FILLCELL_X32 FILLER_142_1743 ();
 FILLCELL_X32 FILLER_142_1775 ();
 FILLCELL_X32 FILLER_142_1807 ();
 FILLCELL_X32 FILLER_142_1839 ();
 FILLCELL_X16 FILLER_142_1871 ();
 FILLCELL_X4 FILLER_142_1887 ();
 FILLCELL_X2 FILLER_142_1891 ();
 FILLCELL_X1 FILLER_142_1893 ();
 FILLCELL_X32 FILLER_142_1895 ();
 FILLCELL_X32 FILLER_142_1927 ();
 FILLCELL_X32 FILLER_142_1959 ();
 FILLCELL_X32 FILLER_142_1991 ();
 FILLCELL_X32 FILLER_142_2023 ();
 FILLCELL_X32 FILLER_142_2055 ();
 FILLCELL_X8 FILLER_142_2087 ();
 FILLCELL_X2 FILLER_142_2095 ();
 FILLCELL_X8 FILLER_142_2100 ();
 FILLCELL_X4 FILLER_142_2108 ();
 FILLCELL_X2 FILLER_142_2112 ();
 FILLCELL_X1 FILLER_142_2114 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X4 FILLER_143_1089 ();
 FILLCELL_X1 FILLER_143_1093 ();
 FILLCELL_X16 FILLER_143_1109 ();
 FILLCELL_X8 FILLER_143_1125 ();
 FILLCELL_X2 FILLER_143_1133 ();
 FILLCELL_X32 FILLER_143_1140 ();
 FILLCELL_X32 FILLER_143_1172 ();
 FILLCELL_X2 FILLER_143_1204 ();
 FILLCELL_X32 FILLER_143_1226 ();
 FILLCELL_X4 FILLER_143_1258 ();
 FILLCELL_X1 FILLER_143_1262 ();
 FILLCELL_X4 FILLER_143_1264 ();
 FILLCELL_X1 FILLER_143_1268 ();
 FILLCELL_X32 FILLER_143_1289 ();
 FILLCELL_X32 FILLER_143_1321 ();
 FILLCELL_X32 FILLER_143_1353 ();
 FILLCELL_X32 FILLER_143_1385 ();
 FILLCELL_X32 FILLER_143_1417 ();
 FILLCELL_X32 FILLER_143_1449 ();
 FILLCELL_X32 FILLER_143_1481 ();
 FILLCELL_X32 FILLER_143_1513 ();
 FILLCELL_X32 FILLER_143_1545 ();
 FILLCELL_X32 FILLER_143_1577 ();
 FILLCELL_X32 FILLER_143_1609 ();
 FILLCELL_X32 FILLER_143_1641 ();
 FILLCELL_X32 FILLER_143_1673 ();
 FILLCELL_X32 FILLER_143_1705 ();
 FILLCELL_X32 FILLER_143_1737 ();
 FILLCELL_X32 FILLER_143_1769 ();
 FILLCELL_X32 FILLER_143_1801 ();
 FILLCELL_X32 FILLER_143_1833 ();
 FILLCELL_X32 FILLER_143_1865 ();
 FILLCELL_X32 FILLER_143_1897 ();
 FILLCELL_X32 FILLER_143_1929 ();
 FILLCELL_X32 FILLER_143_1961 ();
 FILLCELL_X32 FILLER_143_1993 ();
 FILLCELL_X32 FILLER_143_2025 ();
 FILLCELL_X32 FILLER_143_2057 ();
 FILLCELL_X16 FILLER_143_2089 ();
 FILLCELL_X8 FILLER_143_2105 ();
 FILLCELL_X2 FILLER_143_2113 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X8 FILLER_144_984 ();
 FILLCELL_X4 FILLER_144_992 ();
 FILLCELL_X2 FILLER_144_996 ();
 FILLCELL_X8 FILLER_144_1005 ();
 FILLCELL_X4 FILLER_144_1013 ();
 FILLCELL_X8 FILLER_144_1024 ();
 FILLCELL_X4 FILLER_144_1032 ();
 FILLCELL_X1 FILLER_144_1036 ();
 FILLCELL_X16 FILLER_144_1044 ();
 FILLCELL_X8 FILLER_144_1060 ();
 FILLCELL_X4 FILLER_144_1068 ();
 FILLCELL_X32 FILLER_144_1079 ();
 FILLCELL_X16 FILLER_144_1111 ();
 FILLCELL_X8 FILLER_144_1127 ();
 FILLCELL_X2 FILLER_144_1135 ();
 FILLCELL_X8 FILLER_144_1140 ();
 FILLCELL_X2 FILLER_144_1148 ();
 FILLCELL_X1 FILLER_144_1150 ();
 FILLCELL_X8 FILLER_144_1158 ();
 FILLCELL_X4 FILLER_144_1166 ();
 FILLCELL_X2 FILLER_144_1170 ();
 FILLCELL_X32 FILLER_144_1179 ();
 FILLCELL_X32 FILLER_144_1211 ();
 FILLCELL_X32 FILLER_144_1243 ();
 FILLCELL_X32 FILLER_144_1275 ();
 FILLCELL_X32 FILLER_144_1307 ();
 FILLCELL_X32 FILLER_144_1339 ();
 FILLCELL_X32 FILLER_144_1371 ();
 FILLCELL_X32 FILLER_144_1403 ();
 FILLCELL_X32 FILLER_144_1435 ();
 FILLCELL_X32 FILLER_144_1467 ();
 FILLCELL_X32 FILLER_144_1499 ();
 FILLCELL_X32 FILLER_144_1531 ();
 FILLCELL_X32 FILLER_144_1563 ();
 FILLCELL_X32 FILLER_144_1595 ();
 FILLCELL_X32 FILLER_144_1627 ();
 FILLCELL_X32 FILLER_144_1659 ();
 FILLCELL_X32 FILLER_144_1691 ();
 FILLCELL_X32 FILLER_144_1723 ();
 FILLCELL_X32 FILLER_144_1755 ();
 FILLCELL_X32 FILLER_144_1787 ();
 FILLCELL_X32 FILLER_144_1819 ();
 FILLCELL_X32 FILLER_144_1851 ();
 FILLCELL_X8 FILLER_144_1883 ();
 FILLCELL_X2 FILLER_144_1891 ();
 FILLCELL_X1 FILLER_144_1893 ();
 FILLCELL_X32 FILLER_144_1895 ();
 FILLCELL_X32 FILLER_144_1927 ();
 FILLCELL_X32 FILLER_144_1959 ();
 FILLCELL_X32 FILLER_144_1991 ();
 FILLCELL_X32 FILLER_144_2023 ();
 FILLCELL_X32 FILLER_144_2055 ();
 FILLCELL_X16 FILLER_144_2087 ();
 FILLCELL_X8 FILLER_144_2103 ();
 FILLCELL_X4 FILLER_144_2111 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X8 FILLER_145_961 ();
 FILLCELL_X4 FILLER_145_969 ();
 FILLCELL_X4 FILLER_145_980 ();
 FILLCELL_X2 FILLER_145_984 ();
 FILLCELL_X2 FILLER_145_1010 ();
 FILLCELL_X4 FILLER_145_1029 ();
 FILLCELL_X1 FILLER_145_1033 ();
 FILLCELL_X8 FILLER_145_1051 ();
 FILLCELL_X4 FILLER_145_1059 ();
 FILLCELL_X2 FILLER_145_1063 ();
 FILLCELL_X4 FILLER_145_1089 ();
 FILLCELL_X2 FILLER_145_1093 ();
 FILLCELL_X4 FILLER_145_1100 ();
 FILLCELL_X2 FILLER_145_1104 ();
 FILLCELL_X1 FILLER_145_1106 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X16 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1233 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X32 FILLER_145_1584 ();
 FILLCELL_X32 FILLER_145_1616 ();
 FILLCELL_X32 FILLER_145_1648 ();
 FILLCELL_X32 FILLER_145_1680 ();
 FILLCELL_X32 FILLER_145_1712 ();
 FILLCELL_X32 FILLER_145_1744 ();
 FILLCELL_X32 FILLER_145_1776 ();
 FILLCELL_X32 FILLER_145_1808 ();
 FILLCELL_X32 FILLER_145_1840 ();
 FILLCELL_X32 FILLER_145_1872 ();
 FILLCELL_X32 FILLER_145_1904 ();
 FILLCELL_X32 FILLER_145_1936 ();
 FILLCELL_X32 FILLER_145_1968 ();
 FILLCELL_X32 FILLER_145_2000 ();
 FILLCELL_X32 FILLER_145_2032 ();
 FILLCELL_X32 FILLER_145_2064 ();
 FILLCELL_X16 FILLER_145_2096 ();
 FILLCELL_X2 FILLER_145_2112 ();
 FILLCELL_X1 FILLER_145_2114 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X16 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_985 ();
 FILLCELL_X16 FILLER_146_1017 ();
 FILLCELL_X32 FILLER_146_1045 ();
 FILLCELL_X16 FILLER_146_1077 ();
 FILLCELL_X2 FILLER_146_1093 ();
 FILLCELL_X4 FILLER_146_1098 ();
 FILLCELL_X1 FILLER_146_1102 ();
 FILLCELL_X1 FILLER_146_1127 ();
 FILLCELL_X32 FILLER_146_1145 ();
 FILLCELL_X32 FILLER_146_1177 ();
 FILLCELL_X16 FILLER_146_1209 ();
 FILLCELL_X16 FILLER_146_1245 ();
 FILLCELL_X32 FILLER_146_1283 ();
 FILLCELL_X32 FILLER_146_1315 ();
 FILLCELL_X32 FILLER_146_1347 ();
 FILLCELL_X32 FILLER_146_1379 ();
 FILLCELL_X32 FILLER_146_1411 ();
 FILLCELL_X32 FILLER_146_1443 ();
 FILLCELL_X32 FILLER_146_1475 ();
 FILLCELL_X32 FILLER_146_1507 ();
 FILLCELL_X32 FILLER_146_1539 ();
 FILLCELL_X32 FILLER_146_1571 ();
 FILLCELL_X32 FILLER_146_1603 ();
 FILLCELL_X32 FILLER_146_1635 ();
 FILLCELL_X32 FILLER_146_1667 ();
 FILLCELL_X32 FILLER_146_1699 ();
 FILLCELL_X32 FILLER_146_1731 ();
 FILLCELL_X32 FILLER_146_1763 ();
 FILLCELL_X32 FILLER_146_1795 ();
 FILLCELL_X32 FILLER_146_1827 ();
 FILLCELL_X32 FILLER_146_1859 ();
 FILLCELL_X2 FILLER_146_1891 ();
 FILLCELL_X1 FILLER_146_1893 ();
 FILLCELL_X32 FILLER_146_1895 ();
 FILLCELL_X32 FILLER_146_1927 ();
 FILLCELL_X32 FILLER_146_1959 ();
 FILLCELL_X32 FILLER_146_1991 ();
 FILLCELL_X32 FILLER_146_2023 ();
 FILLCELL_X32 FILLER_146_2055 ();
 FILLCELL_X16 FILLER_146_2087 ();
 FILLCELL_X8 FILLER_146_2103 ();
 FILLCELL_X4 FILLER_146_2111 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X16 FILLER_147_993 ();
 FILLCELL_X4 FILLER_147_1009 ();
 FILLCELL_X32 FILLER_147_1017 ();
 FILLCELL_X16 FILLER_147_1049 ();
 FILLCELL_X4 FILLER_147_1065 ();
 FILLCELL_X32 FILLER_147_1093 ();
 FILLCELL_X32 FILLER_147_1125 ();
 FILLCELL_X32 FILLER_147_1157 ();
 FILLCELL_X32 FILLER_147_1189 ();
 FILLCELL_X2 FILLER_147_1221 ();
 FILLCELL_X1 FILLER_147_1223 ();
 FILLCELL_X16 FILLER_147_1244 ();
 FILLCELL_X2 FILLER_147_1260 ();
 FILLCELL_X1 FILLER_147_1262 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X32 FILLER_147_1584 ();
 FILLCELL_X32 FILLER_147_1616 ();
 FILLCELL_X32 FILLER_147_1648 ();
 FILLCELL_X32 FILLER_147_1680 ();
 FILLCELL_X32 FILLER_147_1712 ();
 FILLCELL_X32 FILLER_147_1744 ();
 FILLCELL_X32 FILLER_147_1776 ();
 FILLCELL_X32 FILLER_147_1808 ();
 FILLCELL_X32 FILLER_147_1840 ();
 FILLCELL_X32 FILLER_147_1872 ();
 FILLCELL_X32 FILLER_147_1904 ();
 FILLCELL_X32 FILLER_147_1936 ();
 FILLCELL_X32 FILLER_147_1968 ();
 FILLCELL_X32 FILLER_147_2000 ();
 FILLCELL_X32 FILLER_147_2032 ();
 FILLCELL_X32 FILLER_147_2064 ();
 FILLCELL_X16 FILLER_147_2096 ();
 FILLCELL_X2 FILLER_147_2112 ();
 FILLCELL_X1 FILLER_147_2114 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X8 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_964 ();
 FILLCELL_X32 FILLER_148_996 ();
 FILLCELL_X32 FILLER_148_1028 ();
 FILLCELL_X32 FILLER_148_1060 ();
 FILLCELL_X32 FILLER_148_1092 ();
 FILLCELL_X16 FILLER_148_1124 ();
 FILLCELL_X32 FILLER_148_1147 ();
 FILLCELL_X4 FILLER_148_1179 ();
 FILLCELL_X2 FILLER_148_1183 ();
 FILLCELL_X1 FILLER_148_1185 ();
 FILLCELL_X32 FILLER_148_1214 ();
 FILLCELL_X32 FILLER_148_1266 ();
 FILLCELL_X32 FILLER_148_1298 ();
 FILLCELL_X32 FILLER_148_1330 ();
 FILLCELL_X32 FILLER_148_1362 ();
 FILLCELL_X32 FILLER_148_1394 ();
 FILLCELL_X32 FILLER_148_1426 ();
 FILLCELL_X32 FILLER_148_1458 ();
 FILLCELL_X32 FILLER_148_1490 ();
 FILLCELL_X32 FILLER_148_1522 ();
 FILLCELL_X32 FILLER_148_1554 ();
 FILLCELL_X32 FILLER_148_1586 ();
 FILLCELL_X32 FILLER_148_1618 ();
 FILLCELL_X32 FILLER_148_1650 ();
 FILLCELL_X32 FILLER_148_1682 ();
 FILLCELL_X32 FILLER_148_1714 ();
 FILLCELL_X32 FILLER_148_1746 ();
 FILLCELL_X32 FILLER_148_1778 ();
 FILLCELL_X32 FILLER_148_1810 ();
 FILLCELL_X32 FILLER_148_1842 ();
 FILLCELL_X16 FILLER_148_1874 ();
 FILLCELL_X4 FILLER_148_1890 ();
 FILLCELL_X32 FILLER_148_1895 ();
 FILLCELL_X32 FILLER_148_1927 ();
 FILLCELL_X32 FILLER_148_1959 ();
 FILLCELL_X32 FILLER_148_1991 ();
 FILLCELL_X32 FILLER_148_2023 ();
 FILLCELL_X32 FILLER_148_2055 ();
 FILLCELL_X16 FILLER_148_2087 ();
 FILLCELL_X8 FILLER_148_2103 ();
 FILLCELL_X4 FILLER_148_2111 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X4 FILLER_149_993 ();
 FILLCELL_X2 FILLER_149_997 ();
 FILLCELL_X32 FILLER_149_1023 ();
 FILLCELL_X32 FILLER_149_1055 ();
 FILLCELL_X2 FILLER_149_1087 ();
 FILLCELL_X8 FILLER_149_1096 ();
 FILLCELL_X1 FILLER_149_1104 ();
 FILLCELL_X16 FILLER_149_1112 ();
 FILLCELL_X4 FILLER_149_1128 ();
 FILLCELL_X2 FILLER_149_1132 ();
 FILLCELL_X1 FILLER_149_1134 ();
 FILLCELL_X1 FILLER_149_1152 ();
 FILLCELL_X32 FILLER_149_1177 ();
 FILLCELL_X16 FILLER_149_1209 ();
 FILLCELL_X4 FILLER_149_1225 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X32 FILLER_149_1584 ();
 FILLCELL_X32 FILLER_149_1616 ();
 FILLCELL_X32 FILLER_149_1648 ();
 FILLCELL_X32 FILLER_149_1680 ();
 FILLCELL_X32 FILLER_149_1712 ();
 FILLCELL_X32 FILLER_149_1744 ();
 FILLCELL_X32 FILLER_149_1776 ();
 FILLCELL_X32 FILLER_149_1808 ();
 FILLCELL_X32 FILLER_149_1840 ();
 FILLCELL_X32 FILLER_149_1872 ();
 FILLCELL_X32 FILLER_149_1904 ();
 FILLCELL_X32 FILLER_149_1936 ();
 FILLCELL_X32 FILLER_149_1968 ();
 FILLCELL_X32 FILLER_149_2000 ();
 FILLCELL_X32 FILLER_149_2032 ();
 FILLCELL_X32 FILLER_149_2064 ();
 FILLCELL_X16 FILLER_149_2096 ();
 FILLCELL_X2 FILLER_149_2112 ();
 FILLCELL_X1 FILLER_149_2114 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X16 FILLER_150_952 ();
 FILLCELL_X8 FILLER_150_968 ();
 FILLCELL_X4 FILLER_150_976 ();
 FILLCELL_X2 FILLER_150_980 ();
 FILLCELL_X8 FILLER_150_1006 ();
 FILLCELL_X1 FILLER_150_1014 ();
 FILLCELL_X8 FILLER_150_1022 ();
 FILLCELL_X2 FILLER_150_1030 ();
 FILLCELL_X1 FILLER_150_1032 ();
 FILLCELL_X8 FILLER_150_1040 ();
 FILLCELL_X4 FILLER_150_1048 ();
 FILLCELL_X1 FILLER_150_1052 ();
 FILLCELL_X2 FILLER_150_1060 ();
 FILLCELL_X1 FILLER_150_1062 ();
 FILLCELL_X8 FILLER_150_1070 ();
 FILLCELL_X4 FILLER_150_1078 ();
 FILLCELL_X2 FILLER_150_1082 ();
 FILLCELL_X1 FILLER_150_1084 ();
 FILLCELL_X2 FILLER_150_1102 ();
 FILLCELL_X16 FILLER_150_1121 ();
 FILLCELL_X4 FILLER_150_1137 ();
 FILLCELL_X2 FILLER_150_1141 ();
 FILLCELL_X32 FILLER_150_1150 ();
 FILLCELL_X2 FILLER_150_1182 ();
 FILLCELL_X32 FILLER_150_1204 ();
 FILLCELL_X16 FILLER_150_1236 ();
 FILLCELL_X32 FILLER_150_1274 ();
 FILLCELL_X32 FILLER_150_1306 ();
 FILLCELL_X32 FILLER_150_1338 ();
 FILLCELL_X32 FILLER_150_1370 ();
 FILLCELL_X32 FILLER_150_1402 ();
 FILLCELL_X32 FILLER_150_1434 ();
 FILLCELL_X32 FILLER_150_1466 ();
 FILLCELL_X32 FILLER_150_1498 ();
 FILLCELL_X32 FILLER_150_1530 ();
 FILLCELL_X32 FILLER_150_1562 ();
 FILLCELL_X32 FILLER_150_1594 ();
 FILLCELL_X32 FILLER_150_1626 ();
 FILLCELL_X32 FILLER_150_1658 ();
 FILLCELL_X32 FILLER_150_1690 ();
 FILLCELL_X32 FILLER_150_1722 ();
 FILLCELL_X32 FILLER_150_1754 ();
 FILLCELL_X32 FILLER_150_1786 ();
 FILLCELL_X32 FILLER_150_1818 ();
 FILLCELL_X32 FILLER_150_1850 ();
 FILLCELL_X8 FILLER_150_1882 ();
 FILLCELL_X4 FILLER_150_1890 ();
 FILLCELL_X32 FILLER_150_1895 ();
 FILLCELL_X32 FILLER_150_1927 ();
 FILLCELL_X32 FILLER_150_1959 ();
 FILLCELL_X32 FILLER_150_1991 ();
 FILLCELL_X32 FILLER_150_2023 ();
 FILLCELL_X32 FILLER_150_2055 ();
 FILLCELL_X16 FILLER_150_2087 ();
 FILLCELL_X8 FILLER_150_2103 ();
 FILLCELL_X4 FILLER_150_2111 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X4 FILLER_151_1025 ();
 FILLCELL_X1 FILLER_151_1029 ();
 FILLCELL_X8 FILLER_151_1047 ();
 FILLCELL_X32 FILLER_151_1072 ();
 FILLCELL_X32 FILLER_151_1111 ();
 FILLCELL_X32 FILLER_151_1143 ();
 FILLCELL_X16 FILLER_151_1175 ();
 FILLCELL_X8 FILLER_151_1191 ();
 FILLCELL_X1 FILLER_151_1199 ();
 FILLCELL_X32 FILLER_151_1220 ();
 FILLCELL_X8 FILLER_151_1252 ();
 FILLCELL_X2 FILLER_151_1260 ();
 FILLCELL_X1 FILLER_151_1262 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X32 FILLER_151_1648 ();
 FILLCELL_X32 FILLER_151_1680 ();
 FILLCELL_X32 FILLER_151_1712 ();
 FILLCELL_X32 FILLER_151_1744 ();
 FILLCELL_X32 FILLER_151_1776 ();
 FILLCELL_X32 FILLER_151_1808 ();
 FILLCELL_X32 FILLER_151_1840 ();
 FILLCELL_X32 FILLER_151_1872 ();
 FILLCELL_X32 FILLER_151_1904 ();
 FILLCELL_X32 FILLER_151_1936 ();
 FILLCELL_X32 FILLER_151_1968 ();
 FILLCELL_X32 FILLER_151_2000 ();
 FILLCELL_X32 FILLER_151_2032 ();
 FILLCELL_X32 FILLER_151_2064 ();
 FILLCELL_X16 FILLER_151_2096 ();
 FILLCELL_X2 FILLER_151_2112 ();
 FILLCELL_X1 FILLER_151_2114 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X4 FILLER_152_1080 ();
 FILLCELL_X2 FILLER_152_1084 ();
 FILLCELL_X32 FILLER_152_1093 ();
 FILLCELL_X8 FILLER_152_1125 ();
 FILLCELL_X4 FILLER_152_1133 ();
 FILLCELL_X1 FILLER_152_1137 ();
 FILLCELL_X4 FILLER_152_1150 ();
 FILLCELL_X1 FILLER_152_1154 ();
 FILLCELL_X32 FILLER_152_1162 ();
 FILLCELL_X32 FILLER_152_1194 ();
 FILLCELL_X8 FILLER_152_1226 ();
 FILLCELL_X2 FILLER_152_1234 ();
 FILLCELL_X8 FILLER_152_1256 ();
 FILLCELL_X32 FILLER_152_1286 ();
 FILLCELL_X32 FILLER_152_1318 ();
 FILLCELL_X32 FILLER_152_1350 ();
 FILLCELL_X32 FILLER_152_1382 ();
 FILLCELL_X32 FILLER_152_1414 ();
 FILLCELL_X32 FILLER_152_1446 ();
 FILLCELL_X32 FILLER_152_1478 ();
 FILLCELL_X32 FILLER_152_1510 ();
 FILLCELL_X32 FILLER_152_1542 ();
 FILLCELL_X32 FILLER_152_1574 ();
 FILLCELL_X32 FILLER_152_1606 ();
 FILLCELL_X32 FILLER_152_1638 ();
 FILLCELL_X32 FILLER_152_1670 ();
 FILLCELL_X32 FILLER_152_1702 ();
 FILLCELL_X32 FILLER_152_1734 ();
 FILLCELL_X32 FILLER_152_1766 ();
 FILLCELL_X32 FILLER_152_1798 ();
 FILLCELL_X32 FILLER_152_1830 ();
 FILLCELL_X32 FILLER_152_1862 ();
 FILLCELL_X32 FILLER_152_1895 ();
 FILLCELL_X32 FILLER_152_1927 ();
 FILLCELL_X32 FILLER_152_1959 ();
 FILLCELL_X32 FILLER_152_1991 ();
 FILLCELL_X32 FILLER_152_2023 ();
 FILLCELL_X32 FILLER_152_2055 ();
 FILLCELL_X16 FILLER_152_2087 ();
 FILLCELL_X8 FILLER_152_2103 ();
 FILLCELL_X4 FILLER_152_2111 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X16 FILLER_153_961 ();
 FILLCELL_X16 FILLER_153_984 ();
 FILLCELL_X2 FILLER_153_1000 ();
 FILLCELL_X1 FILLER_153_1002 ();
 FILLCELL_X4 FILLER_153_1010 ();
 FILLCELL_X4 FILLER_153_1021 ();
 FILLCELL_X1 FILLER_153_1025 ();
 FILLCELL_X4 FILLER_153_1031 ();
 FILLCELL_X8 FILLER_153_1071 ();
 FILLCELL_X4 FILLER_153_1079 ();
 FILLCELL_X4 FILLER_153_1100 ();
 FILLCELL_X8 FILLER_153_1109 ();
 FILLCELL_X2 FILLER_153_1117 ();
 FILLCELL_X1 FILLER_153_1119 ();
 FILLCELL_X8 FILLER_153_1123 ();
 FILLCELL_X2 FILLER_153_1131 ();
 FILLCELL_X1 FILLER_153_1133 ();
 FILLCELL_X32 FILLER_153_1175 ();
 FILLCELL_X4 FILLER_153_1207 ();
 FILLCELL_X1 FILLER_153_1211 ();
 FILLCELL_X8 FILLER_153_1234 ();
 FILLCELL_X1 FILLER_153_1242 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X32 FILLER_153_1584 ();
 FILLCELL_X32 FILLER_153_1616 ();
 FILLCELL_X32 FILLER_153_1648 ();
 FILLCELL_X32 FILLER_153_1680 ();
 FILLCELL_X32 FILLER_153_1712 ();
 FILLCELL_X32 FILLER_153_1744 ();
 FILLCELL_X32 FILLER_153_1776 ();
 FILLCELL_X32 FILLER_153_1808 ();
 FILLCELL_X32 FILLER_153_1840 ();
 FILLCELL_X32 FILLER_153_1872 ();
 FILLCELL_X32 FILLER_153_1904 ();
 FILLCELL_X32 FILLER_153_1936 ();
 FILLCELL_X32 FILLER_153_1968 ();
 FILLCELL_X32 FILLER_153_2000 ();
 FILLCELL_X32 FILLER_153_2032 ();
 FILLCELL_X32 FILLER_153_2064 ();
 FILLCELL_X16 FILLER_153_2096 ();
 FILLCELL_X2 FILLER_153_2112 ();
 FILLCELL_X1 FILLER_153_2114 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X16 FILLER_154_952 ();
 FILLCELL_X2 FILLER_154_968 ();
 FILLCELL_X1 FILLER_154_970 ();
 FILLCELL_X4 FILLER_154_988 ();
 FILLCELL_X1 FILLER_154_992 ();
 FILLCELL_X8 FILLER_154_1000 ();
 FILLCELL_X2 FILLER_154_1008 ();
 FILLCELL_X1 FILLER_154_1010 ();
 FILLCELL_X32 FILLER_154_1028 ();
 FILLCELL_X4 FILLER_154_1060 ();
 FILLCELL_X2 FILLER_154_1064 ();
 FILLCELL_X8 FILLER_154_1097 ();
 FILLCELL_X2 FILLER_154_1105 ();
 FILLCELL_X32 FILLER_154_1110 ();
 FILLCELL_X32 FILLER_154_1142 ();
 FILLCELL_X32 FILLER_154_1174 ();
 FILLCELL_X32 FILLER_154_1206 ();
 FILLCELL_X32 FILLER_154_1238 ();
 FILLCELL_X32 FILLER_154_1270 ();
 FILLCELL_X32 FILLER_154_1302 ();
 FILLCELL_X32 FILLER_154_1334 ();
 FILLCELL_X32 FILLER_154_1366 ();
 FILLCELL_X32 FILLER_154_1398 ();
 FILLCELL_X32 FILLER_154_1430 ();
 FILLCELL_X32 FILLER_154_1462 ();
 FILLCELL_X32 FILLER_154_1494 ();
 FILLCELL_X32 FILLER_154_1526 ();
 FILLCELL_X32 FILLER_154_1558 ();
 FILLCELL_X32 FILLER_154_1590 ();
 FILLCELL_X32 FILLER_154_1622 ();
 FILLCELL_X32 FILLER_154_1654 ();
 FILLCELL_X32 FILLER_154_1686 ();
 FILLCELL_X32 FILLER_154_1718 ();
 FILLCELL_X32 FILLER_154_1750 ();
 FILLCELL_X32 FILLER_154_1782 ();
 FILLCELL_X32 FILLER_154_1814 ();
 FILLCELL_X32 FILLER_154_1846 ();
 FILLCELL_X16 FILLER_154_1878 ();
 FILLCELL_X32 FILLER_154_1895 ();
 FILLCELL_X32 FILLER_154_1927 ();
 FILLCELL_X32 FILLER_154_1959 ();
 FILLCELL_X32 FILLER_154_1991 ();
 FILLCELL_X32 FILLER_154_2023 ();
 FILLCELL_X32 FILLER_154_2055 ();
 FILLCELL_X16 FILLER_154_2087 ();
 FILLCELL_X8 FILLER_154_2103 ();
 FILLCELL_X4 FILLER_154_2111 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X16 FILLER_155_929 ();
 FILLCELL_X8 FILLER_155_945 ();
 FILLCELL_X4 FILLER_155_953 ();
 FILLCELL_X2 FILLER_155_957 ();
 FILLCELL_X1 FILLER_155_959 ();
 FILLCELL_X16 FILLER_155_964 ();
 FILLCELL_X8 FILLER_155_980 ();
 FILLCELL_X4 FILLER_155_988 ();
 FILLCELL_X32 FILLER_155_1009 ();
 FILLCELL_X32 FILLER_155_1041 ();
 FILLCELL_X32 FILLER_155_1073 ();
 FILLCELL_X4 FILLER_155_1105 ();
 FILLCELL_X2 FILLER_155_1109 ();
 FILLCELL_X32 FILLER_155_1135 ();
 FILLCELL_X32 FILLER_155_1167 ();
 FILLCELL_X16 FILLER_155_1199 ();
 FILLCELL_X1 FILLER_155_1215 ();
 FILLCELL_X4 FILLER_155_1225 ();
 FILLCELL_X1 FILLER_155_1229 ();
 FILLCELL_X8 FILLER_155_1252 ();
 FILLCELL_X2 FILLER_155_1260 ();
 FILLCELL_X1 FILLER_155_1262 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X32 FILLER_155_1584 ();
 FILLCELL_X32 FILLER_155_1616 ();
 FILLCELL_X32 FILLER_155_1648 ();
 FILLCELL_X32 FILLER_155_1680 ();
 FILLCELL_X32 FILLER_155_1712 ();
 FILLCELL_X32 FILLER_155_1744 ();
 FILLCELL_X32 FILLER_155_1776 ();
 FILLCELL_X32 FILLER_155_1808 ();
 FILLCELL_X32 FILLER_155_1840 ();
 FILLCELL_X32 FILLER_155_1872 ();
 FILLCELL_X32 FILLER_155_1904 ();
 FILLCELL_X32 FILLER_155_1936 ();
 FILLCELL_X32 FILLER_155_1968 ();
 FILLCELL_X32 FILLER_155_2000 ();
 FILLCELL_X32 FILLER_155_2032 ();
 FILLCELL_X32 FILLER_155_2064 ();
 FILLCELL_X16 FILLER_155_2096 ();
 FILLCELL_X2 FILLER_155_2112 ();
 FILLCELL_X1 FILLER_155_2114 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X16 FILLER_156_1080 ();
 FILLCELL_X1 FILLER_156_1096 ();
 FILLCELL_X16 FILLER_156_1121 ();
 FILLCELL_X8 FILLER_156_1137 ();
 FILLCELL_X4 FILLER_156_1152 ();
 FILLCELL_X16 FILLER_156_1163 ();
 FILLCELL_X8 FILLER_156_1179 ();
 FILLCELL_X2 FILLER_156_1187 ();
 FILLCELL_X1 FILLER_156_1189 ();
 FILLCELL_X8 FILLER_156_1212 ();
 FILLCELL_X2 FILLER_156_1220 ();
 FILLCELL_X1 FILLER_156_1222 ();
 FILLCELL_X32 FILLER_156_1243 ();
 FILLCELL_X32 FILLER_156_1275 ();
 FILLCELL_X32 FILLER_156_1307 ();
 FILLCELL_X32 FILLER_156_1339 ();
 FILLCELL_X32 FILLER_156_1371 ();
 FILLCELL_X32 FILLER_156_1403 ();
 FILLCELL_X32 FILLER_156_1435 ();
 FILLCELL_X32 FILLER_156_1467 ();
 FILLCELL_X32 FILLER_156_1499 ();
 FILLCELL_X32 FILLER_156_1531 ();
 FILLCELL_X32 FILLER_156_1563 ();
 FILLCELL_X32 FILLER_156_1595 ();
 FILLCELL_X32 FILLER_156_1627 ();
 FILLCELL_X32 FILLER_156_1659 ();
 FILLCELL_X32 FILLER_156_1691 ();
 FILLCELL_X32 FILLER_156_1723 ();
 FILLCELL_X32 FILLER_156_1755 ();
 FILLCELL_X32 FILLER_156_1787 ();
 FILLCELL_X32 FILLER_156_1819 ();
 FILLCELL_X32 FILLER_156_1851 ();
 FILLCELL_X8 FILLER_156_1883 ();
 FILLCELL_X2 FILLER_156_1891 ();
 FILLCELL_X1 FILLER_156_1893 ();
 FILLCELL_X32 FILLER_156_1895 ();
 FILLCELL_X32 FILLER_156_1927 ();
 FILLCELL_X32 FILLER_156_1959 ();
 FILLCELL_X32 FILLER_156_1991 ();
 FILLCELL_X32 FILLER_156_2023 ();
 FILLCELL_X32 FILLER_156_2055 ();
 FILLCELL_X16 FILLER_156_2087 ();
 FILLCELL_X8 FILLER_156_2103 ();
 FILLCELL_X4 FILLER_156_2111 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X16 FILLER_157_929 ();
 FILLCELL_X1 FILLER_157_945 ();
 FILLCELL_X32 FILLER_157_950 ();
 FILLCELL_X32 FILLER_157_982 ();
 FILLCELL_X32 FILLER_157_1014 ();
 FILLCELL_X16 FILLER_157_1046 ();
 FILLCELL_X4 FILLER_157_1062 ();
 FILLCELL_X16 FILLER_157_1080 ();
 FILLCELL_X8 FILLER_157_1096 ();
 FILLCELL_X4 FILLER_157_1104 ();
 FILLCELL_X2 FILLER_157_1108 ();
 FILLCELL_X16 FILLER_157_1117 ();
 FILLCELL_X8 FILLER_157_1133 ();
 FILLCELL_X1 FILLER_157_1141 ();
 FILLCELL_X8 FILLER_157_1176 ();
 FILLCELL_X4 FILLER_157_1184 ();
 FILLCELL_X16 FILLER_157_1194 ();
 FILLCELL_X2 FILLER_157_1210 ();
 FILLCELL_X16 FILLER_157_1232 ();
 FILLCELL_X8 FILLER_157_1248 ();
 FILLCELL_X4 FILLER_157_1256 ();
 FILLCELL_X2 FILLER_157_1260 ();
 FILLCELL_X1 FILLER_157_1262 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X32 FILLER_157_1584 ();
 FILLCELL_X32 FILLER_157_1616 ();
 FILLCELL_X32 FILLER_157_1648 ();
 FILLCELL_X32 FILLER_157_1680 ();
 FILLCELL_X32 FILLER_157_1712 ();
 FILLCELL_X32 FILLER_157_1744 ();
 FILLCELL_X32 FILLER_157_1776 ();
 FILLCELL_X32 FILLER_157_1808 ();
 FILLCELL_X32 FILLER_157_1840 ();
 FILLCELL_X32 FILLER_157_1872 ();
 FILLCELL_X32 FILLER_157_1904 ();
 FILLCELL_X32 FILLER_157_1936 ();
 FILLCELL_X32 FILLER_157_1968 ();
 FILLCELL_X32 FILLER_157_2000 ();
 FILLCELL_X32 FILLER_157_2032 ();
 FILLCELL_X32 FILLER_157_2064 ();
 FILLCELL_X16 FILLER_157_2096 ();
 FILLCELL_X2 FILLER_157_2112 ();
 FILLCELL_X1 FILLER_157_2114 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X16 FILLER_158_952 ();
 FILLCELL_X4 FILLER_158_968 ();
 FILLCELL_X16 FILLER_158_979 ();
 FILLCELL_X8 FILLER_158_995 ();
 FILLCELL_X16 FILLER_158_1034 ();
 FILLCELL_X1 FILLER_158_1050 ();
 FILLCELL_X32 FILLER_158_1085 ();
 FILLCELL_X16 FILLER_158_1117 ();
 FILLCELL_X8 FILLER_158_1133 ();
 FILLCELL_X4 FILLER_158_1141 ();
 FILLCELL_X1 FILLER_158_1145 ();
 FILLCELL_X32 FILLER_158_1153 ();
 FILLCELL_X2 FILLER_158_1185 ();
 FILLCELL_X32 FILLER_158_1193 ();
 FILLCELL_X32 FILLER_158_1225 ();
 FILLCELL_X32 FILLER_158_1257 ();
 FILLCELL_X32 FILLER_158_1289 ();
 FILLCELL_X32 FILLER_158_1321 ();
 FILLCELL_X32 FILLER_158_1353 ();
 FILLCELL_X32 FILLER_158_1385 ();
 FILLCELL_X32 FILLER_158_1417 ();
 FILLCELL_X32 FILLER_158_1449 ();
 FILLCELL_X32 FILLER_158_1481 ();
 FILLCELL_X32 FILLER_158_1513 ();
 FILLCELL_X32 FILLER_158_1545 ();
 FILLCELL_X32 FILLER_158_1577 ();
 FILLCELL_X32 FILLER_158_1609 ();
 FILLCELL_X32 FILLER_158_1641 ();
 FILLCELL_X32 FILLER_158_1673 ();
 FILLCELL_X32 FILLER_158_1705 ();
 FILLCELL_X32 FILLER_158_1737 ();
 FILLCELL_X32 FILLER_158_1769 ();
 FILLCELL_X32 FILLER_158_1801 ();
 FILLCELL_X32 FILLER_158_1833 ();
 FILLCELL_X16 FILLER_158_1865 ();
 FILLCELL_X8 FILLER_158_1881 ();
 FILLCELL_X4 FILLER_158_1889 ();
 FILLCELL_X1 FILLER_158_1893 ();
 FILLCELL_X32 FILLER_158_1895 ();
 FILLCELL_X32 FILLER_158_1927 ();
 FILLCELL_X32 FILLER_158_1959 ();
 FILLCELL_X32 FILLER_158_1991 ();
 FILLCELL_X32 FILLER_158_2023 ();
 FILLCELL_X32 FILLER_158_2055 ();
 FILLCELL_X16 FILLER_158_2087 ();
 FILLCELL_X8 FILLER_158_2103 ();
 FILLCELL_X4 FILLER_158_2111 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X8 FILLER_159_929 ();
 FILLCELL_X16 FILLER_159_941 ();
 FILLCELL_X8 FILLER_159_957 ();
 FILLCELL_X1 FILLER_159_965 ();
 FILLCELL_X2 FILLER_159_1007 ();
 FILLCELL_X1 FILLER_159_1009 ();
 FILLCELL_X32 FILLER_159_1039 ();
 FILLCELL_X2 FILLER_159_1071 ();
 FILLCELL_X1 FILLER_159_1073 ();
 FILLCELL_X16 FILLER_159_1081 ();
 FILLCELL_X4 FILLER_159_1097 ();
 FILLCELL_X4 FILLER_159_1104 ();
 FILLCELL_X2 FILLER_159_1108 ();
 FILLCELL_X1 FILLER_159_1110 ();
 FILLCELL_X2 FILLER_159_1116 ();
 FILLCELL_X8 FILLER_159_1125 ();
 FILLCELL_X4 FILLER_159_1133 ();
 FILLCELL_X1 FILLER_159_1137 ();
 FILLCELL_X32 FILLER_159_1145 ();
 FILLCELL_X8 FILLER_159_1177 ();
 FILLCELL_X4 FILLER_159_1185 ();
 FILLCELL_X16 FILLER_159_1245 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X32 FILLER_159_1584 ();
 FILLCELL_X32 FILLER_159_1616 ();
 FILLCELL_X32 FILLER_159_1648 ();
 FILLCELL_X32 FILLER_159_1680 ();
 FILLCELL_X32 FILLER_159_1712 ();
 FILLCELL_X32 FILLER_159_1744 ();
 FILLCELL_X32 FILLER_159_1776 ();
 FILLCELL_X32 FILLER_159_1808 ();
 FILLCELL_X32 FILLER_159_1840 ();
 FILLCELL_X32 FILLER_159_1872 ();
 FILLCELL_X32 FILLER_159_1904 ();
 FILLCELL_X32 FILLER_159_1936 ();
 FILLCELL_X32 FILLER_159_1968 ();
 FILLCELL_X32 FILLER_159_2000 ();
 FILLCELL_X32 FILLER_159_2032 ();
 FILLCELL_X32 FILLER_159_2064 ();
 FILLCELL_X16 FILLER_159_2096 ();
 FILLCELL_X2 FILLER_159_2112 ();
 FILLCELL_X1 FILLER_159_2114 ();
 FILLCELL_X8 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_34 ();
 FILLCELL_X32 FILLER_160_66 ();
 FILLCELL_X32 FILLER_160_98 ();
 FILLCELL_X32 FILLER_160_130 ();
 FILLCELL_X32 FILLER_160_162 ();
 FILLCELL_X32 FILLER_160_194 ();
 FILLCELL_X32 FILLER_160_226 ();
 FILLCELL_X32 FILLER_160_258 ();
 FILLCELL_X32 FILLER_160_290 ();
 FILLCELL_X32 FILLER_160_322 ();
 FILLCELL_X32 FILLER_160_354 ();
 FILLCELL_X32 FILLER_160_386 ();
 FILLCELL_X32 FILLER_160_418 ();
 FILLCELL_X32 FILLER_160_450 ();
 FILLCELL_X32 FILLER_160_482 ();
 FILLCELL_X32 FILLER_160_514 ();
 FILLCELL_X32 FILLER_160_546 ();
 FILLCELL_X32 FILLER_160_578 ();
 FILLCELL_X16 FILLER_160_610 ();
 FILLCELL_X4 FILLER_160_626 ();
 FILLCELL_X1 FILLER_160_630 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X2 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1025 ();
 FILLCELL_X32 FILLER_160_1057 ();
 FILLCELL_X8 FILLER_160_1089 ();
 FILLCELL_X2 FILLER_160_1097 ();
 FILLCELL_X4 FILLER_160_1106 ();
 FILLCELL_X2 FILLER_160_1110 ();
 FILLCELL_X2 FILLER_160_1119 ();
 FILLCELL_X32 FILLER_160_1138 ();
 FILLCELL_X4 FILLER_160_1170 ();
 FILLCELL_X2 FILLER_160_1174 ();
 FILLCELL_X1 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1184 ();
 FILLCELL_X32 FILLER_160_1244 ();
 FILLCELL_X32 FILLER_160_1276 ();
 FILLCELL_X32 FILLER_160_1308 ();
 FILLCELL_X32 FILLER_160_1340 ();
 FILLCELL_X32 FILLER_160_1372 ();
 FILLCELL_X32 FILLER_160_1404 ();
 FILLCELL_X32 FILLER_160_1436 ();
 FILLCELL_X32 FILLER_160_1468 ();
 FILLCELL_X32 FILLER_160_1500 ();
 FILLCELL_X32 FILLER_160_1532 ();
 FILLCELL_X32 FILLER_160_1564 ();
 FILLCELL_X32 FILLER_160_1596 ();
 FILLCELL_X32 FILLER_160_1628 ();
 FILLCELL_X32 FILLER_160_1660 ();
 FILLCELL_X32 FILLER_160_1692 ();
 FILLCELL_X32 FILLER_160_1724 ();
 FILLCELL_X32 FILLER_160_1756 ();
 FILLCELL_X32 FILLER_160_1788 ();
 FILLCELL_X32 FILLER_160_1820 ();
 FILLCELL_X32 FILLER_160_1852 ();
 FILLCELL_X8 FILLER_160_1884 ();
 FILLCELL_X2 FILLER_160_1892 ();
 FILLCELL_X32 FILLER_160_1895 ();
 FILLCELL_X32 FILLER_160_1927 ();
 FILLCELL_X32 FILLER_160_1959 ();
 FILLCELL_X32 FILLER_160_1991 ();
 FILLCELL_X32 FILLER_160_2023 ();
 FILLCELL_X32 FILLER_160_2055 ();
 FILLCELL_X16 FILLER_160_2087 ();
 FILLCELL_X8 FILLER_160_2103 ();
 FILLCELL_X4 FILLER_160_2111 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X4 FILLER_161_993 ();
 FILLCELL_X2 FILLER_161_997 ();
 FILLCELL_X1 FILLER_161_999 ();
 FILLCELL_X32 FILLER_161_1007 ();
 FILLCELL_X8 FILLER_161_1039 ();
 FILLCELL_X4 FILLER_161_1047 ();
 FILLCELL_X1 FILLER_161_1051 ();
 FILLCELL_X16 FILLER_161_1059 ();
 FILLCELL_X2 FILLER_161_1075 ();
 FILLCELL_X8 FILLER_161_1084 ();
 FILLCELL_X2 FILLER_161_1092 ();
 FILLCELL_X1 FILLER_161_1094 ();
 FILLCELL_X32 FILLER_161_1112 ();
 FILLCELL_X4 FILLER_161_1144 ();
 FILLCELL_X2 FILLER_161_1148 ();
 FILLCELL_X4 FILLER_161_1174 ();
 FILLCELL_X2 FILLER_161_1178 ();
 FILLCELL_X1 FILLER_161_1180 ();
 FILLCELL_X16 FILLER_161_1188 ();
 FILLCELL_X8 FILLER_161_1204 ();
 FILLCELL_X4 FILLER_161_1212 ();
 FILLCELL_X2 FILLER_161_1216 ();
 FILLCELL_X1 FILLER_161_1218 ();
 FILLCELL_X16 FILLER_161_1236 ();
 FILLCELL_X8 FILLER_161_1252 ();
 FILLCELL_X2 FILLER_161_1260 ();
 FILLCELL_X1 FILLER_161_1262 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X32 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1520 ();
 FILLCELL_X32 FILLER_161_1552 ();
 FILLCELL_X32 FILLER_161_1584 ();
 FILLCELL_X32 FILLER_161_1616 ();
 FILLCELL_X32 FILLER_161_1648 ();
 FILLCELL_X32 FILLER_161_1680 ();
 FILLCELL_X32 FILLER_161_1712 ();
 FILLCELL_X32 FILLER_161_1744 ();
 FILLCELL_X32 FILLER_161_1776 ();
 FILLCELL_X32 FILLER_161_1808 ();
 FILLCELL_X32 FILLER_161_1840 ();
 FILLCELL_X32 FILLER_161_1872 ();
 FILLCELL_X32 FILLER_161_1904 ();
 FILLCELL_X32 FILLER_161_1936 ();
 FILLCELL_X32 FILLER_161_1968 ();
 FILLCELL_X32 FILLER_161_2000 ();
 FILLCELL_X32 FILLER_161_2032 ();
 FILLCELL_X32 FILLER_161_2064 ();
 FILLCELL_X16 FILLER_161_2096 ();
 FILLCELL_X2 FILLER_161_2112 ();
 FILLCELL_X1 FILLER_161_2114 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X16 FILLER_162_952 ();
 FILLCELL_X8 FILLER_162_968 ();
 FILLCELL_X1 FILLER_162_976 ();
 FILLCELL_X8 FILLER_162_984 ();
 FILLCELL_X4 FILLER_162_992 ();
 FILLCELL_X1 FILLER_162_996 ();
 FILLCELL_X16 FILLER_162_1014 ();
 FILLCELL_X4 FILLER_162_1030 ();
 FILLCELL_X4 FILLER_162_1041 ();
 FILLCELL_X1 FILLER_162_1045 ();
 FILLCELL_X8 FILLER_162_1063 ();
 FILLCELL_X1 FILLER_162_1071 ();
 FILLCELL_X4 FILLER_162_1089 ();
 FILLCELL_X2 FILLER_162_1093 ();
 FILLCELL_X16 FILLER_162_1100 ();
 FILLCELL_X8 FILLER_162_1116 ();
 FILLCELL_X4 FILLER_162_1124 ();
 FILLCELL_X4 FILLER_162_1154 ();
 FILLCELL_X8 FILLER_162_1165 ();
 FILLCELL_X4 FILLER_162_1173 ();
 FILLCELL_X2 FILLER_162_1177 ();
 FILLCELL_X1 FILLER_162_1179 ();
 FILLCELL_X8 FILLER_162_1184 ();
 FILLCELL_X1 FILLER_162_1192 ();
 FILLCELL_X32 FILLER_162_1199 ();
 FILLCELL_X32 FILLER_162_1231 ();
 FILLCELL_X32 FILLER_162_1263 ();
 FILLCELL_X32 FILLER_162_1295 ();
 FILLCELL_X32 FILLER_162_1327 ();
 FILLCELL_X32 FILLER_162_1359 ();
 FILLCELL_X32 FILLER_162_1391 ();
 FILLCELL_X32 FILLER_162_1423 ();
 FILLCELL_X32 FILLER_162_1455 ();
 FILLCELL_X32 FILLER_162_1487 ();
 FILLCELL_X32 FILLER_162_1519 ();
 FILLCELL_X32 FILLER_162_1551 ();
 FILLCELL_X32 FILLER_162_1583 ();
 FILLCELL_X32 FILLER_162_1615 ();
 FILLCELL_X32 FILLER_162_1647 ();
 FILLCELL_X32 FILLER_162_1679 ();
 FILLCELL_X32 FILLER_162_1711 ();
 FILLCELL_X32 FILLER_162_1743 ();
 FILLCELL_X32 FILLER_162_1775 ();
 FILLCELL_X32 FILLER_162_1807 ();
 FILLCELL_X32 FILLER_162_1839 ();
 FILLCELL_X16 FILLER_162_1871 ();
 FILLCELL_X4 FILLER_162_1887 ();
 FILLCELL_X2 FILLER_162_1891 ();
 FILLCELL_X1 FILLER_162_1893 ();
 FILLCELL_X32 FILLER_162_1895 ();
 FILLCELL_X32 FILLER_162_1927 ();
 FILLCELL_X32 FILLER_162_1959 ();
 FILLCELL_X32 FILLER_162_1991 ();
 FILLCELL_X32 FILLER_162_2023 ();
 FILLCELL_X32 FILLER_162_2055 ();
 FILLCELL_X16 FILLER_162_2087 ();
 FILLCELL_X8 FILLER_162_2103 ();
 FILLCELL_X4 FILLER_162_2111 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X8 FILLER_163_961 ();
 FILLCELL_X4 FILLER_163_969 ();
 FILLCELL_X1 FILLER_163_973 ();
 FILLCELL_X8 FILLER_163_991 ();
 FILLCELL_X4 FILLER_163_999 ();
 FILLCELL_X1 FILLER_163_1003 ();
 FILLCELL_X16 FILLER_163_1011 ();
 FILLCELL_X2 FILLER_163_1027 ();
 FILLCELL_X16 FILLER_163_1034 ();
 FILLCELL_X4 FILLER_163_1050 ();
 FILLCELL_X2 FILLER_163_1054 ();
 FILLCELL_X16 FILLER_163_1063 ();
 FILLCELL_X4 FILLER_163_1079 ();
 FILLCELL_X4 FILLER_163_1090 ();
 FILLCELL_X1 FILLER_163_1094 ();
 FILLCELL_X16 FILLER_163_1098 ();
 FILLCELL_X1 FILLER_163_1114 ();
 FILLCELL_X2 FILLER_163_1123 ();
 FILLCELL_X1 FILLER_163_1125 ();
 FILLCELL_X2 FILLER_163_1147 ();
 FILLCELL_X16 FILLER_163_1156 ();
 FILLCELL_X8 FILLER_163_1172 ();
 FILLCELL_X1 FILLER_163_1180 ();
 FILLCELL_X16 FILLER_163_1194 ();
 FILLCELL_X8 FILLER_163_1210 ();
 FILLCELL_X2 FILLER_163_1218 ();
 FILLCELL_X1 FILLER_163_1227 ();
 FILLCELL_X8 FILLER_163_1250 ();
 FILLCELL_X4 FILLER_163_1258 ();
 FILLCELL_X1 FILLER_163_1262 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X32 FILLER_163_1584 ();
 FILLCELL_X32 FILLER_163_1616 ();
 FILLCELL_X32 FILLER_163_1648 ();
 FILLCELL_X32 FILLER_163_1680 ();
 FILLCELL_X32 FILLER_163_1712 ();
 FILLCELL_X32 FILLER_163_1744 ();
 FILLCELL_X32 FILLER_163_1776 ();
 FILLCELL_X32 FILLER_163_1808 ();
 FILLCELL_X32 FILLER_163_1840 ();
 FILLCELL_X32 FILLER_163_1872 ();
 FILLCELL_X32 FILLER_163_1904 ();
 FILLCELL_X32 FILLER_163_1936 ();
 FILLCELL_X32 FILLER_163_1968 ();
 FILLCELL_X32 FILLER_163_2000 ();
 FILLCELL_X32 FILLER_163_2032 ();
 FILLCELL_X32 FILLER_163_2064 ();
 FILLCELL_X16 FILLER_163_2096 ();
 FILLCELL_X2 FILLER_163_2112 ();
 FILLCELL_X1 FILLER_163_2114 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X8 FILLER_164_984 ();
 FILLCELL_X2 FILLER_164_992 ();
 FILLCELL_X4 FILLER_164_1018 ();
 FILLCELL_X2 FILLER_164_1022 ();
 FILLCELL_X16 FILLER_164_1031 ();
 FILLCELL_X4 FILLER_164_1047 ();
 FILLCELL_X2 FILLER_164_1051 ();
 FILLCELL_X16 FILLER_164_1060 ();
 FILLCELL_X4 FILLER_164_1076 ();
 FILLCELL_X1 FILLER_164_1080 ();
 FILLCELL_X8 FILLER_164_1088 ();
 FILLCELL_X1 FILLER_164_1096 ();
 FILLCELL_X4 FILLER_164_1104 ();
 FILLCELL_X2 FILLER_164_1108 ();
 FILLCELL_X1 FILLER_164_1110 ();
 FILLCELL_X32 FILLER_164_1118 ();
 FILLCELL_X8 FILLER_164_1167 ();
 FILLCELL_X2 FILLER_164_1175 ();
 FILLCELL_X16 FILLER_164_1202 ();
 FILLCELL_X4 FILLER_164_1218 ();
 FILLCELL_X32 FILLER_164_1231 ();
 FILLCELL_X32 FILLER_164_1263 ();
 FILLCELL_X32 FILLER_164_1295 ();
 FILLCELL_X32 FILLER_164_1327 ();
 FILLCELL_X32 FILLER_164_1359 ();
 FILLCELL_X32 FILLER_164_1391 ();
 FILLCELL_X32 FILLER_164_1423 ();
 FILLCELL_X32 FILLER_164_1455 ();
 FILLCELL_X32 FILLER_164_1487 ();
 FILLCELL_X32 FILLER_164_1519 ();
 FILLCELL_X32 FILLER_164_1551 ();
 FILLCELL_X32 FILLER_164_1583 ();
 FILLCELL_X32 FILLER_164_1615 ();
 FILLCELL_X32 FILLER_164_1647 ();
 FILLCELL_X32 FILLER_164_1679 ();
 FILLCELL_X32 FILLER_164_1711 ();
 FILLCELL_X32 FILLER_164_1743 ();
 FILLCELL_X32 FILLER_164_1775 ();
 FILLCELL_X32 FILLER_164_1807 ();
 FILLCELL_X32 FILLER_164_1839 ();
 FILLCELL_X16 FILLER_164_1871 ();
 FILLCELL_X4 FILLER_164_1887 ();
 FILLCELL_X2 FILLER_164_1891 ();
 FILLCELL_X1 FILLER_164_1893 ();
 FILLCELL_X32 FILLER_164_1895 ();
 FILLCELL_X32 FILLER_164_1927 ();
 FILLCELL_X32 FILLER_164_1959 ();
 FILLCELL_X32 FILLER_164_1991 ();
 FILLCELL_X32 FILLER_164_2023 ();
 FILLCELL_X32 FILLER_164_2055 ();
 FILLCELL_X16 FILLER_164_2087 ();
 FILLCELL_X8 FILLER_164_2103 ();
 FILLCELL_X4 FILLER_164_2111 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X8 FILLER_165_993 ();
 FILLCELL_X4 FILLER_165_1001 ();
 FILLCELL_X1 FILLER_165_1005 ();
 FILLCELL_X16 FILLER_165_1030 ();
 FILLCELL_X2 FILLER_165_1046 ();
 FILLCELL_X4 FILLER_165_1065 ();
 FILLCELL_X32 FILLER_165_1086 ();
 FILLCELL_X4 FILLER_165_1118 ();
 FILLCELL_X1 FILLER_165_1122 ();
 FILLCELL_X32 FILLER_165_1130 ();
 FILLCELL_X32 FILLER_165_1162 ();
 FILLCELL_X8 FILLER_165_1194 ();
 FILLCELL_X1 FILLER_165_1202 ();
 FILLCELL_X32 FILLER_165_1218 ();
 FILLCELL_X8 FILLER_165_1250 ();
 FILLCELL_X4 FILLER_165_1258 ();
 FILLCELL_X1 FILLER_165_1262 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X32 FILLER_165_1584 ();
 FILLCELL_X32 FILLER_165_1616 ();
 FILLCELL_X32 FILLER_165_1648 ();
 FILLCELL_X32 FILLER_165_1680 ();
 FILLCELL_X32 FILLER_165_1712 ();
 FILLCELL_X32 FILLER_165_1744 ();
 FILLCELL_X32 FILLER_165_1776 ();
 FILLCELL_X32 FILLER_165_1808 ();
 FILLCELL_X32 FILLER_165_1840 ();
 FILLCELL_X32 FILLER_165_1872 ();
 FILLCELL_X32 FILLER_165_1904 ();
 FILLCELL_X32 FILLER_165_1936 ();
 FILLCELL_X32 FILLER_165_1968 ();
 FILLCELL_X32 FILLER_165_2000 ();
 FILLCELL_X32 FILLER_165_2032 ();
 FILLCELL_X32 FILLER_165_2064 ();
 FILLCELL_X16 FILLER_165_2096 ();
 FILLCELL_X2 FILLER_165_2112 ();
 FILLCELL_X1 FILLER_165_2114 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X16 FILLER_166_1048 ();
 FILLCELL_X4 FILLER_166_1064 ();
 FILLCELL_X2 FILLER_166_1068 ();
 FILLCELL_X16 FILLER_166_1074 ();
 FILLCELL_X8 FILLER_166_1090 ();
 FILLCELL_X4 FILLER_166_1115 ();
 FILLCELL_X2 FILLER_166_1119 ();
 FILLCELL_X1 FILLER_166_1121 ();
 FILLCELL_X32 FILLER_166_1139 ();
 FILLCELL_X16 FILLER_166_1171 ();
 FILLCELL_X4 FILLER_166_1187 ();
 FILLCELL_X8 FILLER_166_1201 ();
 FILLCELL_X2 FILLER_166_1209 ();
 FILLCELL_X32 FILLER_166_1227 ();
 FILLCELL_X32 FILLER_166_1259 ();
 FILLCELL_X32 FILLER_166_1291 ();
 FILLCELL_X32 FILLER_166_1323 ();
 FILLCELL_X32 FILLER_166_1355 ();
 FILLCELL_X32 FILLER_166_1387 ();
 FILLCELL_X32 FILLER_166_1419 ();
 FILLCELL_X32 FILLER_166_1451 ();
 FILLCELL_X32 FILLER_166_1483 ();
 FILLCELL_X32 FILLER_166_1515 ();
 FILLCELL_X32 FILLER_166_1547 ();
 FILLCELL_X32 FILLER_166_1579 ();
 FILLCELL_X32 FILLER_166_1611 ();
 FILLCELL_X32 FILLER_166_1643 ();
 FILLCELL_X32 FILLER_166_1675 ();
 FILLCELL_X32 FILLER_166_1707 ();
 FILLCELL_X32 FILLER_166_1739 ();
 FILLCELL_X32 FILLER_166_1771 ();
 FILLCELL_X32 FILLER_166_1803 ();
 FILLCELL_X32 FILLER_166_1835 ();
 FILLCELL_X16 FILLER_166_1867 ();
 FILLCELL_X8 FILLER_166_1883 ();
 FILLCELL_X2 FILLER_166_1891 ();
 FILLCELL_X1 FILLER_166_1893 ();
 FILLCELL_X32 FILLER_166_1895 ();
 FILLCELL_X32 FILLER_166_1927 ();
 FILLCELL_X32 FILLER_166_1959 ();
 FILLCELL_X32 FILLER_166_1991 ();
 FILLCELL_X32 FILLER_166_2023 ();
 FILLCELL_X32 FILLER_166_2055 ();
 FILLCELL_X16 FILLER_166_2087 ();
 FILLCELL_X8 FILLER_166_2103 ();
 FILLCELL_X4 FILLER_166_2111 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X32 FILLER_167_801 ();
 FILLCELL_X32 FILLER_167_833 ();
 FILLCELL_X32 FILLER_167_865 ();
 FILLCELL_X32 FILLER_167_897 ();
 FILLCELL_X32 FILLER_167_929 ();
 FILLCELL_X32 FILLER_167_961 ();
 FILLCELL_X32 FILLER_167_993 ();
 FILLCELL_X32 FILLER_167_1025 ();
 FILLCELL_X32 FILLER_167_1057 ();
 FILLCELL_X32 FILLER_167_1089 ();
 FILLCELL_X16 FILLER_167_1121 ();
 FILLCELL_X4 FILLER_167_1137 ();
 FILLCELL_X2 FILLER_167_1141 ();
 FILLCELL_X1 FILLER_167_1143 ();
 FILLCELL_X2 FILLER_167_1171 ();
 FILLCELL_X4 FILLER_167_1178 ();
 FILLCELL_X1 FILLER_167_1182 ();
 FILLCELL_X8 FILLER_167_1198 ();
 FILLCELL_X4 FILLER_167_1206 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X8 FILLER_167_1249 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X32 FILLER_167_1584 ();
 FILLCELL_X32 FILLER_167_1616 ();
 FILLCELL_X32 FILLER_167_1648 ();
 FILLCELL_X32 FILLER_167_1680 ();
 FILLCELL_X32 FILLER_167_1712 ();
 FILLCELL_X32 FILLER_167_1744 ();
 FILLCELL_X32 FILLER_167_1776 ();
 FILLCELL_X32 FILLER_167_1808 ();
 FILLCELL_X32 FILLER_167_1840 ();
 FILLCELL_X32 FILLER_167_1872 ();
 FILLCELL_X32 FILLER_167_1904 ();
 FILLCELL_X32 FILLER_167_1936 ();
 FILLCELL_X32 FILLER_167_1968 ();
 FILLCELL_X32 FILLER_167_2000 ();
 FILLCELL_X32 FILLER_167_2032 ();
 FILLCELL_X32 FILLER_167_2064 ();
 FILLCELL_X16 FILLER_167_2096 ();
 FILLCELL_X2 FILLER_167_2112 ();
 FILLCELL_X1 FILLER_167_2114 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X4 FILLER_168_1176 ();
 FILLCELL_X16 FILLER_168_1187 ();
 FILLCELL_X8 FILLER_168_1203 ();
 FILLCELL_X4 FILLER_168_1211 ();
 FILLCELL_X32 FILLER_168_1233 ();
 FILLCELL_X32 FILLER_168_1265 ();
 FILLCELL_X32 FILLER_168_1297 ();
 FILLCELL_X32 FILLER_168_1329 ();
 FILLCELL_X32 FILLER_168_1361 ();
 FILLCELL_X32 FILLER_168_1393 ();
 FILLCELL_X32 FILLER_168_1425 ();
 FILLCELL_X32 FILLER_168_1457 ();
 FILLCELL_X32 FILLER_168_1489 ();
 FILLCELL_X32 FILLER_168_1521 ();
 FILLCELL_X32 FILLER_168_1553 ();
 FILLCELL_X32 FILLER_168_1585 ();
 FILLCELL_X32 FILLER_168_1617 ();
 FILLCELL_X32 FILLER_168_1649 ();
 FILLCELL_X32 FILLER_168_1681 ();
 FILLCELL_X32 FILLER_168_1713 ();
 FILLCELL_X32 FILLER_168_1745 ();
 FILLCELL_X32 FILLER_168_1777 ();
 FILLCELL_X32 FILLER_168_1809 ();
 FILLCELL_X32 FILLER_168_1841 ();
 FILLCELL_X16 FILLER_168_1873 ();
 FILLCELL_X4 FILLER_168_1889 ();
 FILLCELL_X1 FILLER_168_1893 ();
 FILLCELL_X32 FILLER_168_1895 ();
 FILLCELL_X32 FILLER_168_1927 ();
 FILLCELL_X32 FILLER_168_1959 ();
 FILLCELL_X32 FILLER_168_1991 ();
 FILLCELL_X32 FILLER_168_2023 ();
 FILLCELL_X32 FILLER_168_2055 ();
 FILLCELL_X16 FILLER_168_2087 ();
 FILLCELL_X8 FILLER_168_2103 ();
 FILLCELL_X4 FILLER_168_2111 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X32 FILLER_169_577 ();
 FILLCELL_X32 FILLER_169_609 ();
 FILLCELL_X32 FILLER_169_641 ();
 FILLCELL_X32 FILLER_169_673 ();
 FILLCELL_X32 FILLER_169_705 ();
 FILLCELL_X32 FILLER_169_737 ();
 FILLCELL_X32 FILLER_169_769 ();
 FILLCELL_X32 FILLER_169_801 ();
 FILLCELL_X32 FILLER_169_833 ();
 FILLCELL_X32 FILLER_169_865 ();
 FILLCELL_X32 FILLER_169_897 ();
 FILLCELL_X32 FILLER_169_929 ();
 FILLCELL_X32 FILLER_169_961 ();
 FILLCELL_X32 FILLER_169_993 ();
 FILLCELL_X32 FILLER_169_1025 ();
 FILLCELL_X32 FILLER_169_1057 ();
 FILLCELL_X8 FILLER_169_1089 ();
 FILLCELL_X4 FILLER_169_1097 ();
 FILLCELL_X8 FILLER_169_1108 ();
 FILLCELL_X2 FILLER_169_1116 ();
 FILLCELL_X1 FILLER_169_1118 ();
 FILLCELL_X32 FILLER_169_1126 ();
 FILLCELL_X16 FILLER_169_1158 ();
 FILLCELL_X4 FILLER_169_1174 ();
 FILLCELL_X2 FILLER_169_1178 ();
 FILLCELL_X16 FILLER_169_1200 ();
 FILLCELL_X1 FILLER_169_1216 ();
 FILLCELL_X32 FILLER_169_1229 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X32 FILLER_169_1584 ();
 FILLCELL_X32 FILLER_169_1616 ();
 FILLCELL_X32 FILLER_169_1648 ();
 FILLCELL_X32 FILLER_169_1680 ();
 FILLCELL_X32 FILLER_169_1712 ();
 FILLCELL_X32 FILLER_169_1744 ();
 FILLCELL_X32 FILLER_169_1776 ();
 FILLCELL_X32 FILLER_169_1808 ();
 FILLCELL_X32 FILLER_169_1840 ();
 FILLCELL_X32 FILLER_169_1872 ();
 FILLCELL_X32 FILLER_169_1904 ();
 FILLCELL_X32 FILLER_169_1936 ();
 FILLCELL_X32 FILLER_169_1968 ();
 FILLCELL_X32 FILLER_169_2000 ();
 FILLCELL_X32 FILLER_169_2032 ();
 FILLCELL_X32 FILLER_169_2064 ();
 FILLCELL_X16 FILLER_169_2096 ();
 FILLCELL_X2 FILLER_169_2112 ();
 FILLCELL_X1 FILLER_169_2114 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X32 FILLER_170_1048 ();
 FILLCELL_X16 FILLER_170_1080 ();
 FILLCELL_X2 FILLER_170_1096 ();
 FILLCELL_X1 FILLER_170_1098 ();
 FILLCELL_X2 FILLER_170_1121 ();
 FILLCELL_X32 FILLER_170_1145 ();
 FILLCELL_X32 FILLER_170_1177 ();
 FILLCELL_X4 FILLER_170_1209 ();
 FILLCELL_X32 FILLER_170_1229 ();
 FILLCELL_X32 FILLER_170_1261 ();
 FILLCELL_X32 FILLER_170_1293 ();
 FILLCELL_X32 FILLER_170_1325 ();
 FILLCELL_X32 FILLER_170_1357 ();
 FILLCELL_X32 FILLER_170_1389 ();
 FILLCELL_X32 FILLER_170_1421 ();
 FILLCELL_X32 FILLER_170_1453 ();
 FILLCELL_X32 FILLER_170_1485 ();
 FILLCELL_X32 FILLER_170_1517 ();
 FILLCELL_X32 FILLER_170_1549 ();
 FILLCELL_X32 FILLER_170_1581 ();
 FILLCELL_X32 FILLER_170_1613 ();
 FILLCELL_X32 FILLER_170_1645 ();
 FILLCELL_X32 FILLER_170_1677 ();
 FILLCELL_X32 FILLER_170_1709 ();
 FILLCELL_X32 FILLER_170_1741 ();
 FILLCELL_X32 FILLER_170_1773 ();
 FILLCELL_X32 FILLER_170_1805 ();
 FILLCELL_X32 FILLER_170_1837 ();
 FILLCELL_X16 FILLER_170_1869 ();
 FILLCELL_X8 FILLER_170_1885 ();
 FILLCELL_X1 FILLER_170_1893 ();
 FILLCELL_X32 FILLER_170_1895 ();
 FILLCELL_X32 FILLER_170_1927 ();
 FILLCELL_X32 FILLER_170_1959 ();
 FILLCELL_X32 FILLER_170_1991 ();
 FILLCELL_X32 FILLER_170_2023 ();
 FILLCELL_X32 FILLER_170_2055 ();
 FILLCELL_X16 FILLER_170_2087 ();
 FILLCELL_X8 FILLER_170_2103 ();
 FILLCELL_X4 FILLER_170_2111 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X32 FILLER_171_353 ();
 FILLCELL_X32 FILLER_171_385 ();
 FILLCELL_X32 FILLER_171_417 ();
 FILLCELL_X32 FILLER_171_449 ();
 FILLCELL_X32 FILLER_171_481 ();
 FILLCELL_X32 FILLER_171_513 ();
 FILLCELL_X32 FILLER_171_545 ();
 FILLCELL_X32 FILLER_171_577 ();
 FILLCELL_X32 FILLER_171_609 ();
 FILLCELL_X32 FILLER_171_641 ();
 FILLCELL_X32 FILLER_171_673 ();
 FILLCELL_X32 FILLER_171_705 ();
 FILLCELL_X32 FILLER_171_737 ();
 FILLCELL_X32 FILLER_171_769 ();
 FILLCELL_X32 FILLER_171_801 ();
 FILLCELL_X32 FILLER_171_833 ();
 FILLCELL_X32 FILLER_171_865 ();
 FILLCELL_X32 FILLER_171_897 ();
 FILLCELL_X32 FILLER_171_929 ();
 FILLCELL_X32 FILLER_171_961 ();
 FILLCELL_X32 FILLER_171_993 ();
 FILLCELL_X32 FILLER_171_1025 ();
 FILLCELL_X32 FILLER_171_1057 ();
 FILLCELL_X32 FILLER_171_1089 ();
 FILLCELL_X32 FILLER_171_1121 ();
 FILLCELL_X32 FILLER_171_1153 ();
 FILLCELL_X16 FILLER_171_1185 ();
 FILLCELL_X8 FILLER_171_1201 ();
 FILLCELL_X2 FILLER_171_1209 ();
 FILLCELL_X32 FILLER_171_1220 ();
 FILLCELL_X8 FILLER_171_1252 ();
 FILLCELL_X2 FILLER_171_1260 ();
 FILLCELL_X1 FILLER_171_1262 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X32 FILLER_171_1584 ();
 FILLCELL_X32 FILLER_171_1616 ();
 FILLCELL_X32 FILLER_171_1648 ();
 FILLCELL_X32 FILLER_171_1680 ();
 FILLCELL_X32 FILLER_171_1712 ();
 FILLCELL_X32 FILLER_171_1744 ();
 FILLCELL_X32 FILLER_171_1776 ();
 FILLCELL_X32 FILLER_171_1808 ();
 FILLCELL_X32 FILLER_171_1840 ();
 FILLCELL_X32 FILLER_171_1872 ();
 FILLCELL_X32 FILLER_171_1904 ();
 FILLCELL_X32 FILLER_171_1936 ();
 FILLCELL_X32 FILLER_171_1968 ();
 FILLCELL_X32 FILLER_171_2000 ();
 FILLCELL_X32 FILLER_171_2032 ();
 FILLCELL_X32 FILLER_171_2064 ();
 FILLCELL_X16 FILLER_171_2096 ();
 FILLCELL_X2 FILLER_171_2112 ();
 FILLCELL_X1 FILLER_171_2114 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X16 FILLER_172_1080 ();
 FILLCELL_X4 FILLER_172_1096 ();
 FILLCELL_X16 FILLER_172_1107 ();
 FILLCELL_X2 FILLER_172_1123 ();
 FILLCELL_X32 FILLER_172_1132 ();
 FILLCELL_X32 FILLER_172_1164 ();
 FILLCELL_X32 FILLER_172_1196 ();
 FILLCELL_X32 FILLER_172_1228 ();
 FILLCELL_X32 FILLER_172_1260 ();
 FILLCELL_X32 FILLER_172_1292 ();
 FILLCELL_X32 FILLER_172_1324 ();
 FILLCELL_X32 FILLER_172_1356 ();
 FILLCELL_X32 FILLER_172_1388 ();
 FILLCELL_X32 FILLER_172_1420 ();
 FILLCELL_X32 FILLER_172_1452 ();
 FILLCELL_X32 FILLER_172_1484 ();
 FILLCELL_X32 FILLER_172_1516 ();
 FILLCELL_X32 FILLER_172_1548 ();
 FILLCELL_X32 FILLER_172_1580 ();
 FILLCELL_X32 FILLER_172_1612 ();
 FILLCELL_X32 FILLER_172_1644 ();
 FILLCELL_X32 FILLER_172_1676 ();
 FILLCELL_X32 FILLER_172_1708 ();
 FILLCELL_X32 FILLER_172_1740 ();
 FILLCELL_X32 FILLER_172_1772 ();
 FILLCELL_X32 FILLER_172_1804 ();
 FILLCELL_X32 FILLER_172_1836 ();
 FILLCELL_X16 FILLER_172_1868 ();
 FILLCELL_X8 FILLER_172_1884 ();
 FILLCELL_X2 FILLER_172_1892 ();
 FILLCELL_X32 FILLER_172_1895 ();
 FILLCELL_X32 FILLER_172_1927 ();
 FILLCELL_X32 FILLER_172_1959 ();
 FILLCELL_X32 FILLER_172_1991 ();
 FILLCELL_X32 FILLER_172_2023 ();
 FILLCELL_X32 FILLER_172_2055 ();
 FILLCELL_X16 FILLER_172_2087 ();
 FILLCELL_X8 FILLER_172_2103 ();
 FILLCELL_X4 FILLER_172_2111 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X8 FILLER_173_1089 ();
 FILLCELL_X2 FILLER_173_1097 ();
 FILLCELL_X4 FILLER_173_1121 ();
 FILLCELL_X2 FILLER_173_1125 ();
 FILLCELL_X1 FILLER_173_1127 ();
 FILLCELL_X32 FILLER_173_1150 ();
 FILLCELL_X32 FILLER_173_1182 ();
 FILLCELL_X32 FILLER_173_1214 ();
 FILLCELL_X16 FILLER_173_1246 ();
 FILLCELL_X1 FILLER_173_1262 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X32 FILLER_173_1584 ();
 FILLCELL_X32 FILLER_173_1616 ();
 FILLCELL_X32 FILLER_173_1648 ();
 FILLCELL_X32 FILLER_173_1680 ();
 FILLCELL_X32 FILLER_173_1712 ();
 FILLCELL_X32 FILLER_173_1744 ();
 FILLCELL_X32 FILLER_173_1776 ();
 FILLCELL_X32 FILLER_173_1808 ();
 FILLCELL_X32 FILLER_173_1840 ();
 FILLCELL_X32 FILLER_173_1872 ();
 FILLCELL_X32 FILLER_173_1904 ();
 FILLCELL_X32 FILLER_173_1936 ();
 FILLCELL_X32 FILLER_173_1968 ();
 FILLCELL_X32 FILLER_173_2000 ();
 FILLCELL_X32 FILLER_173_2032 ();
 FILLCELL_X32 FILLER_173_2064 ();
 FILLCELL_X16 FILLER_173_2096 ();
 FILLCELL_X2 FILLER_173_2112 ();
 FILLCELL_X1 FILLER_173_2114 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X32 FILLER_174_1304 ();
 FILLCELL_X32 FILLER_174_1336 ();
 FILLCELL_X32 FILLER_174_1368 ();
 FILLCELL_X32 FILLER_174_1400 ();
 FILLCELL_X32 FILLER_174_1432 ();
 FILLCELL_X32 FILLER_174_1464 ();
 FILLCELL_X32 FILLER_174_1496 ();
 FILLCELL_X32 FILLER_174_1528 ();
 FILLCELL_X32 FILLER_174_1560 ();
 FILLCELL_X32 FILLER_174_1592 ();
 FILLCELL_X32 FILLER_174_1624 ();
 FILLCELL_X32 FILLER_174_1656 ();
 FILLCELL_X32 FILLER_174_1688 ();
 FILLCELL_X32 FILLER_174_1720 ();
 FILLCELL_X32 FILLER_174_1752 ();
 FILLCELL_X32 FILLER_174_1784 ();
 FILLCELL_X32 FILLER_174_1816 ();
 FILLCELL_X32 FILLER_174_1848 ();
 FILLCELL_X8 FILLER_174_1880 ();
 FILLCELL_X4 FILLER_174_1888 ();
 FILLCELL_X2 FILLER_174_1892 ();
 FILLCELL_X32 FILLER_174_1895 ();
 FILLCELL_X32 FILLER_174_1927 ();
 FILLCELL_X32 FILLER_174_1959 ();
 FILLCELL_X32 FILLER_174_1991 ();
 FILLCELL_X32 FILLER_174_2023 ();
 FILLCELL_X32 FILLER_174_2055 ();
 FILLCELL_X16 FILLER_174_2087 ();
 FILLCELL_X8 FILLER_174_2103 ();
 FILLCELL_X4 FILLER_174_2111 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X32 FILLER_175_385 ();
 FILLCELL_X32 FILLER_175_417 ();
 FILLCELL_X32 FILLER_175_449 ();
 FILLCELL_X32 FILLER_175_481 ();
 FILLCELL_X32 FILLER_175_513 ();
 FILLCELL_X32 FILLER_175_545 ();
 FILLCELL_X32 FILLER_175_577 ();
 FILLCELL_X32 FILLER_175_609 ();
 FILLCELL_X32 FILLER_175_641 ();
 FILLCELL_X32 FILLER_175_673 ();
 FILLCELL_X32 FILLER_175_705 ();
 FILLCELL_X32 FILLER_175_737 ();
 FILLCELL_X32 FILLER_175_769 ();
 FILLCELL_X32 FILLER_175_801 ();
 FILLCELL_X32 FILLER_175_833 ();
 FILLCELL_X32 FILLER_175_865 ();
 FILLCELL_X32 FILLER_175_897 ();
 FILLCELL_X32 FILLER_175_929 ();
 FILLCELL_X32 FILLER_175_961 ();
 FILLCELL_X32 FILLER_175_993 ();
 FILLCELL_X32 FILLER_175_1025 ();
 FILLCELL_X32 FILLER_175_1057 ();
 FILLCELL_X32 FILLER_175_1089 ();
 FILLCELL_X32 FILLER_175_1121 ();
 FILLCELL_X32 FILLER_175_1153 ();
 FILLCELL_X32 FILLER_175_1185 ();
 FILLCELL_X32 FILLER_175_1217 ();
 FILLCELL_X8 FILLER_175_1249 ();
 FILLCELL_X4 FILLER_175_1257 ();
 FILLCELL_X2 FILLER_175_1261 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X32 FILLER_175_1584 ();
 FILLCELL_X32 FILLER_175_1616 ();
 FILLCELL_X32 FILLER_175_1648 ();
 FILLCELL_X32 FILLER_175_1680 ();
 FILLCELL_X32 FILLER_175_1712 ();
 FILLCELL_X32 FILLER_175_1744 ();
 FILLCELL_X32 FILLER_175_1776 ();
 FILLCELL_X32 FILLER_175_1808 ();
 FILLCELL_X32 FILLER_175_1840 ();
 FILLCELL_X32 FILLER_175_1872 ();
 FILLCELL_X32 FILLER_175_1904 ();
 FILLCELL_X32 FILLER_175_1936 ();
 FILLCELL_X32 FILLER_175_1968 ();
 FILLCELL_X32 FILLER_175_2000 ();
 FILLCELL_X32 FILLER_175_2032 ();
 FILLCELL_X32 FILLER_175_2064 ();
 FILLCELL_X16 FILLER_175_2096 ();
 FILLCELL_X2 FILLER_175_2112 ();
 FILLCELL_X1 FILLER_175_2114 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X32 FILLER_176_353 ();
 FILLCELL_X32 FILLER_176_385 ();
 FILLCELL_X32 FILLER_176_417 ();
 FILLCELL_X32 FILLER_176_449 ();
 FILLCELL_X32 FILLER_176_481 ();
 FILLCELL_X32 FILLER_176_513 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X32 FILLER_176_577 ();
 FILLCELL_X16 FILLER_176_609 ();
 FILLCELL_X4 FILLER_176_625 ();
 FILLCELL_X2 FILLER_176_629 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X16 FILLER_176_1080 ();
 FILLCELL_X4 FILLER_176_1096 ();
 FILLCELL_X2 FILLER_176_1100 ();
 FILLCELL_X8 FILLER_176_1109 ();
 FILLCELL_X4 FILLER_176_1117 ();
 FILLCELL_X32 FILLER_176_1128 ();
 FILLCELL_X32 FILLER_176_1160 ();
 FILLCELL_X32 FILLER_176_1192 ();
 FILLCELL_X32 FILLER_176_1224 ();
 FILLCELL_X32 FILLER_176_1256 ();
 FILLCELL_X32 FILLER_176_1288 ();
 FILLCELL_X32 FILLER_176_1320 ();
 FILLCELL_X32 FILLER_176_1352 ();
 FILLCELL_X32 FILLER_176_1384 ();
 FILLCELL_X32 FILLER_176_1416 ();
 FILLCELL_X32 FILLER_176_1448 ();
 FILLCELL_X32 FILLER_176_1480 ();
 FILLCELL_X32 FILLER_176_1512 ();
 FILLCELL_X32 FILLER_176_1544 ();
 FILLCELL_X32 FILLER_176_1576 ();
 FILLCELL_X32 FILLER_176_1608 ();
 FILLCELL_X32 FILLER_176_1640 ();
 FILLCELL_X32 FILLER_176_1672 ();
 FILLCELL_X32 FILLER_176_1704 ();
 FILLCELL_X32 FILLER_176_1736 ();
 FILLCELL_X32 FILLER_176_1768 ();
 FILLCELL_X32 FILLER_176_1800 ();
 FILLCELL_X32 FILLER_176_1832 ();
 FILLCELL_X16 FILLER_176_1864 ();
 FILLCELL_X8 FILLER_176_1880 ();
 FILLCELL_X4 FILLER_176_1888 ();
 FILLCELL_X2 FILLER_176_1892 ();
 FILLCELL_X32 FILLER_176_1895 ();
 FILLCELL_X32 FILLER_176_1927 ();
 FILLCELL_X32 FILLER_176_1959 ();
 FILLCELL_X32 FILLER_176_1991 ();
 FILLCELL_X32 FILLER_176_2023 ();
 FILLCELL_X32 FILLER_176_2055 ();
 FILLCELL_X16 FILLER_176_2087 ();
 FILLCELL_X8 FILLER_176_2103 ();
 FILLCELL_X4 FILLER_176_2111 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X8 FILLER_177_1089 ();
 FILLCELL_X2 FILLER_177_1097 ();
 FILLCELL_X32 FILLER_177_1143 ();
 FILLCELL_X32 FILLER_177_1175 ();
 FILLCELL_X32 FILLER_177_1207 ();
 FILLCELL_X16 FILLER_177_1239 ();
 FILLCELL_X8 FILLER_177_1255 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X32 FILLER_177_1584 ();
 FILLCELL_X32 FILLER_177_1616 ();
 FILLCELL_X32 FILLER_177_1648 ();
 FILLCELL_X32 FILLER_177_1680 ();
 FILLCELL_X32 FILLER_177_1712 ();
 FILLCELL_X32 FILLER_177_1744 ();
 FILLCELL_X32 FILLER_177_1776 ();
 FILLCELL_X32 FILLER_177_1808 ();
 FILLCELL_X32 FILLER_177_1840 ();
 FILLCELL_X32 FILLER_177_1872 ();
 FILLCELL_X32 FILLER_177_1904 ();
 FILLCELL_X32 FILLER_177_1936 ();
 FILLCELL_X32 FILLER_177_1968 ();
 FILLCELL_X32 FILLER_177_2000 ();
 FILLCELL_X32 FILLER_177_2032 ();
 FILLCELL_X32 FILLER_177_2064 ();
 FILLCELL_X16 FILLER_177_2096 ();
 FILLCELL_X2 FILLER_177_2112 ();
 FILLCELL_X1 FILLER_177_2114 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X32 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1144 ();
 FILLCELL_X32 FILLER_178_1176 ();
 FILLCELL_X32 FILLER_178_1208 ();
 FILLCELL_X32 FILLER_178_1240 ();
 FILLCELL_X32 FILLER_178_1272 ();
 FILLCELL_X32 FILLER_178_1304 ();
 FILLCELL_X32 FILLER_178_1336 ();
 FILLCELL_X32 FILLER_178_1368 ();
 FILLCELL_X32 FILLER_178_1400 ();
 FILLCELL_X32 FILLER_178_1432 ();
 FILLCELL_X32 FILLER_178_1464 ();
 FILLCELL_X32 FILLER_178_1496 ();
 FILLCELL_X32 FILLER_178_1528 ();
 FILLCELL_X32 FILLER_178_1560 ();
 FILLCELL_X32 FILLER_178_1592 ();
 FILLCELL_X32 FILLER_178_1624 ();
 FILLCELL_X32 FILLER_178_1656 ();
 FILLCELL_X32 FILLER_178_1688 ();
 FILLCELL_X32 FILLER_178_1720 ();
 FILLCELL_X32 FILLER_178_1752 ();
 FILLCELL_X32 FILLER_178_1784 ();
 FILLCELL_X32 FILLER_178_1816 ();
 FILLCELL_X32 FILLER_178_1848 ();
 FILLCELL_X8 FILLER_178_1880 ();
 FILLCELL_X4 FILLER_178_1888 ();
 FILLCELL_X2 FILLER_178_1892 ();
 FILLCELL_X32 FILLER_178_1895 ();
 FILLCELL_X32 FILLER_178_1927 ();
 FILLCELL_X32 FILLER_178_1959 ();
 FILLCELL_X32 FILLER_178_1991 ();
 FILLCELL_X32 FILLER_178_2023 ();
 FILLCELL_X32 FILLER_178_2055 ();
 FILLCELL_X16 FILLER_178_2087 ();
 FILLCELL_X8 FILLER_178_2103 ();
 FILLCELL_X4 FILLER_178_2111 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X32 FILLER_179_1089 ();
 FILLCELL_X32 FILLER_179_1121 ();
 FILLCELL_X32 FILLER_179_1153 ();
 FILLCELL_X32 FILLER_179_1185 ();
 FILLCELL_X32 FILLER_179_1217 ();
 FILLCELL_X8 FILLER_179_1249 ();
 FILLCELL_X4 FILLER_179_1257 ();
 FILLCELL_X2 FILLER_179_1261 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X32 FILLER_179_1584 ();
 FILLCELL_X32 FILLER_179_1616 ();
 FILLCELL_X32 FILLER_179_1648 ();
 FILLCELL_X32 FILLER_179_1680 ();
 FILLCELL_X32 FILLER_179_1712 ();
 FILLCELL_X32 FILLER_179_1744 ();
 FILLCELL_X32 FILLER_179_1776 ();
 FILLCELL_X32 FILLER_179_1808 ();
 FILLCELL_X32 FILLER_179_1840 ();
 FILLCELL_X32 FILLER_179_1872 ();
 FILLCELL_X32 FILLER_179_1904 ();
 FILLCELL_X32 FILLER_179_1936 ();
 FILLCELL_X32 FILLER_179_1968 ();
 FILLCELL_X32 FILLER_179_2000 ();
 FILLCELL_X32 FILLER_179_2032 ();
 FILLCELL_X32 FILLER_179_2064 ();
 FILLCELL_X16 FILLER_179_2096 ();
 FILLCELL_X2 FILLER_179_2112 ();
 FILLCELL_X1 FILLER_179_2114 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X32 FILLER_180_353 ();
 FILLCELL_X32 FILLER_180_385 ();
 FILLCELL_X32 FILLER_180_417 ();
 FILLCELL_X32 FILLER_180_449 ();
 FILLCELL_X32 FILLER_180_481 ();
 FILLCELL_X32 FILLER_180_513 ();
 FILLCELL_X32 FILLER_180_545 ();
 FILLCELL_X32 FILLER_180_577 ();
 FILLCELL_X16 FILLER_180_609 ();
 FILLCELL_X4 FILLER_180_625 ();
 FILLCELL_X2 FILLER_180_629 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X32 FILLER_180_1080 ();
 FILLCELL_X32 FILLER_180_1112 ();
 FILLCELL_X32 FILLER_180_1144 ();
 FILLCELL_X32 FILLER_180_1176 ();
 FILLCELL_X32 FILLER_180_1208 ();
 FILLCELL_X32 FILLER_180_1240 ();
 FILLCELL_X32 FILLER_180_1272 ();
 FILLCELL_X32 FILLER_180_1304 ();
 FILLCELL_X32 FILLER_180_1336 ();
 FILLCELL_X32 FILLER_180_1368 ();
 FILLCELL_X32 FILLER_180_1400 ();
 FILLCELL_X32 FILLER_180_1432 ();
 FILLCELL_X32 FILLER_180_1464 ();
 FILLCELL_X32 FILLER_180_1496 ();
 FILLCELL_X32 FILLER_180_1528 ();
 FILLCELL_X32 FILLER_180_1560 ();
 FILLCELL_X32 FILLER_180_1592 ();
 FILLCELL_X32 FILLER_180_1624 ();
 FILLCELL_X32 FILLER_180_1656 ();
 FILLCELL_X32 FILLER_180_1688 ();
 FILLCELL_X32 FILLER_180_1720 ();
 FILLCELL_X32 FILLER_180_1752 ();
 FILLCELL_X32 FILLER_180_1784 ();
 FILLCELL_X32 FILLER_180_1816 ();
 FILLCELL_X32 FILLER_180_1848 ();
 FILLCELL_X8 FILLER_180_1880 ();
 FILLCELL_X4 FILLER_180_1888 ();
 FILLCELL_X2 FILLER_180_1892 ();
 FILLCELL_X32 FILLER_180_1895 ();
 FILLCELL_X32 FILLER_180_1927 ();
 FILLCELL_X32 FILLER_180_1959 ();
 FILLCELL_X32 FILLER_180_1991 ();
 FILLCELL_X32 FILLER_180_2023 ();
 FILLCELL_X32 FILLER_180_2055 ();
 FILLCELL_X16 FILLER_180_2087 ();
 FILLCELL_X8 FILLER_180_2103 ();
 FILLCELL_X4 FILLER_180_2111 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X32 FILLER_181_1089 ();
 FILLCELL_X32 FILLER_181_1121 ();
 FILLCELL_X32 FILLER_181_1153 ();
 FILLCELL_X32 FILLER_181_1185 ();
 FILLCELL_X32 FILLER_181_1217 ();
 FILLCELL_X8 FILLER_181_1249 ();
 FILLCELL_X4 FILLER_181_1257 ();
 FILLCELL_X2 FILLER_181_1261 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X32 FILLER_181_1584 ();
 FILLCELL_X32 FILLER_181_1616 ();
 FILLCELL_X32 FILLER_181_1648 ();
 FILLCELL_X32 FILLER_181_1680 ();
 FILLCELL_X32 FILLER_181_1712 ();
 FILLCELL_X32 FILLER_181_1744 ();
 FILLCELL_X32 FILLER_181_1776 ();
 FILLCELL_X32 FILLER_181_1808 ();
 FILLCELL_X32 FILLER_181_1840 ();
 FILLCELL_X32 FILLER_181_1872 ();
 FILLCELL_X32 FILLER_181_1904 ();
 FILLCELL_X32 FILLER_181_1936 ();
 FILLCELL_X32 FILLER_181_1968 ();
 FILLCELL_X32 FILLER_181_2000 ();
 FILLCELL_X32 FILLER_181_2032 ();
 FILLCELL_X32 FILLER_181_2064 ();
 FILLCELL_X16 FILLER_181_2096 ();
 FILLCELL_X2 FILLER_181_2112 ();
 FILLCELL_X1 FILLER_181_2114 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X32 FILLER_182_1080 ();
 FILLCELL_X32 FILLER_182_1112 ();
 FILLCELL_X32 FILLER_182_1144 ();
 FILLCELL_X32 FILLER_182_1176 ();
 FILLCELL_X32 FILLER_182_1208 ();
 FILLCELL_X32 FILLER_182_1240 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X32 FILLER_182_1400 ();
 FILLCELL_X32 FILLER_182_1432 ();
 FILLCELL_X32 FILLER_182_1464 ();
 FILLCELL_X32 FILLER_182_1496 ();
 FILLCELL_X32 FILLER_182_1528 ();
 FILLCELL_X32 FILLER_182_1560 ();
 FILLCELL_X32 FILLER_182_1592 ();
 FILLCELL_X32 FILLER_182_1624 ();
 FILLCELL_X32 FILLER_182_1656 ();
 FILLCELL_X32 FILLER_182_1688 ();
 FILLCELL_X32 FILLER_182_1720 ();
 FILLCELL_X32 FILLER_182_1752 ();
 FILLCELL_X32 FILLER_182_1784 ();
 FILLCELL_X32 FILLER_182_1816 ();
 FILLCELL_X32 FILLER_182_1848 ();
 FILLCELL_X8 FILLER_182_1880 ();
 FILLCELL_X4 FILLER_182_1888 ();
 FILLCELL_X2 FILLER_182_1892 ();
 FILLCELL_X32 FILLER_182_1895 ();
 FILLCELL_X32 FILLER_182_1927 ();
 FILLCELL_X32 FILLER_182_1959 ();
 FILLCELL_X32 FILLER_182_1991 ();
 FILLCELL_X32 FILLER_182_2023 ();
 FILLCELL_X32 FILLER_182_2055 ();
 FILLCELL_X16 FILLER_182_2087 ();
 FILLCELL_X8 FILLER_182_2103 ();
 FILLCELL_X4 FILLER_182_2111 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X32 FILLER_183_1089 ();
 FILLCELL_X32 FILLER_183_1121 ();
 FILLCELL_X32 FILLER_183_1153 ();
 FILLCELL_X32 FILLER_183_1185 ();
 FILLCELL_X32 FILLER_183_1217 ();
 FILLCELL_X8 FILLER_183_1249 ();
 FILLCELL_X4 FILLER_183_1257 ();
 FILLCELL_X2 FILLER_183_1261 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X32 FILLER_183_1584 ();
 FILLCELL_X32 FILLER_183_1616 ();
 FILLCELL_X32 FILLER_183_1648 ();
 FILLCELL_X32 FILLER_183_1680 ();
 FILLCELL_X32 FILLER_183_1712 ();
 FILLCELL_X32 FILLER_183_1744 ();
 FILLCELL_X32 FILLER_183_1776 ();
 FILLCELL_X32 FILLER_183_1808 ();
 FILLCELL_X32 FILLER_183_1840 ();
 FILLCELL_X32 FILLER_183_1872 ();
 FILLCELL_X32 FILLER_183_1904 ();
 FILLCELL_X32 FILLER_183_1936 ();
 FILLCELL_X32 FILLER_183_1968 ();
 FILLCELL_X32 FILLER_183_2000 ();
 FILLCELL_X32 FILLER_183_2032 ();
 FILLCELL_X32 FILLER_183_2064 ();
 FILLCELL_X16 FILLER_183_2096 ();
 FILLCELL_X2 FILLER_183_2112 ();
 FILLCELL_X1 FILLER_183_2114 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X32 FILLER_184_1144 ();
 FILLCELL_X32 FILLER_184_1176 ();
 FILLCELL_X32 FILLER_184_1208 ();
 FILLCELL_X32 FILLER_184_1240 ();
 FILLCELL_X32 FILLER_184_1272 ();
 FILLCELL_X32 FILLER_184_1304 ();
 FILLCELL_X32 FILLER_184_1336 ();
 FILLCELL_X32 FILLER_184_1368 ();
 FILLCELL_X32 FILLER_184_1400 ();
 FILLCELL_X32 FILLER_184_1432 ();
 FILLCELL_X32 FILLER_184_1464 ();
 FILLCELL_X32 FILLER_184_1496 ();
 FILLCELL_X32 FILLER_184_1528 ();
 FILLCELL_X32 FILLER_184_1560 ();
 FILLCELL_X32 FILLER_184_1592 ();
 FILLCELL_X32 FILLER_184_1624 ();
 FILLCELL_X32 FILLER_184_1656 ();
 FILLCELL_X32 FILLER_184_1688 ();
 FILLCELL_X32 FILLER_184_1720 ();
 FILLCELL_X32 FILLER_184_1752 ();
 FILLCELL_X32 FILLER_184_1784 ();
 FILLCELL_X32 FILLER_184_1816 ();
 FILLCELL_X32 FILLER_184_1848 ();
 FILLCELL_X8 FILLER_184_1880 ();
 FILLCELL_X4 FILLER_184_1888 ();
 FILLCELL_X2 FILLER_184_1892 ();
 FILLCELL_X32 FILLER_184_1895 ();
 FILLCELL_X32 FILLER_184_1927 ();
 FILLCELL_X32 FILLER_184_1959 ();
 FILLCELL_X32 FILLER_184_1991 ();
 FILLCELL_X32 FILLER_184_2023 ();
 FILLCELL_X32 FILLER_184_2055 ();
 FILLCELL_X16 FILLER_184_2087 ();
 FILLCELL_X8 FILLER_184_2103 ();
 FILLCELL_X4 FILLER_184_2111 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X32 FILLER_185_1185 ();
 FILLCELL_X32 FILLER_185_1217 ();
 FILLCELL_X8 FILLER_185_1249 ();
 FILLCELL_X4 FILLER_185_1257 ();
 FILLCELL_X2 FILLER_185_1261 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X32 FILLER_185_1584 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X32 FILLER_185_1648 ();
 FILLCELL_X32 FILLER_185_1680 ();
 FILLCELL_X32 FILLER_185_1712 ();
 FILLCELL_X32 FILLER_185_1744 ();
 FILLCELL_X32 FILLER_185_1776 ();
 FILLCELL_X32 FILLER_185_1808 ();
 FILLCELL_X32 FILLER_185_1840 ();
 FILLCELL_X32 FILLER_185_1872 ();
 FILLCELL_X32 FILLER_185_1904 ();
 FILLCELL_X32 FILLER_185_1936 ();
 FILLCELL_X32 FILLER_185_1968 ();
 FILLCELL_X32 FILLER_185_2000 ();
 FILLCELL_X32 FILLER_185_2032 ();
 FILLCELL_X32 FILLER_185_2064 ();
 FILLCELL_X16 FILLER_185_2096 ();
 FILLCELL_X2 FILLER_185_2112 ();
 FILLCELL_X1 FILLER_185_2114 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X32 FILLER_186_1240 ();
 FILLCELL_X32 FILLER_186_1272 ();
 FILLCELL_X32 FILLER_186_1304 ();
 FILLCELL_X32 FILLER_186_1336 ();
 FILLCELL_X32 FILLER_186_1368 ();
 FILLCELL_X32 FILLER_186_1400 ();
 FILLCELL_X32 FILLER_186_1432 ();
 FILLCELL_X32 FILLER_186_1464 ();
 FILLCELL_X32 FILLER_186_1496 ();
 FILLCELL_X32 FILLER_186_1528 ();
 FILLCELL_X32 FILLER_186_1560 ();
 FILLCELL_X32 FILLER_186_1592 ();
 FILLCELL_X32 FILLER_186_1624 ();
 FILLCELL_X32 FILLER_186_1656 ();
 FILLCELL_X32 FILLER_186_1688 ();
 FILLCELL_X32 FILLER_186_1720 ();
 FILLCELL_X32 FILLER_186_1752 ();
 FILLCELL_X32 FILLER_186_1784 ();
 FILLCELL_X32 FILLER_186_1816 ();
 FILLCELL_X32 FILLER_186_1848 ();
 FILLCELL_X8 FILLER_186_1880 ();
 FILLCELL_X4 FILLER_186_1888 ();
 FILLCELL_X2 FILLER_186_1892 ();
 FILLCELL_X32 FILLER_186_1895 ();
 FILLCELL_X32 FILLER_186_1927 ();
 FILLCELL_X32 FILLER_186_1959 ();
 FILLCELL_X32 FILLER_186_1991 ();
 FILLCELL_X32 FILLER_186_2023 ();
 FILLCELL_X32 FILLER_186_2055 ();
 FILLCELL_X16 FILLER_186_2087 ();
 FILLCELL_X8 FILLER_186_2103 ();
 FILLCELL_X4 FILLER_186_2111 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X32 FILLER_187_1217 ();
 FILLCELL_X8 FILLER_187_1249 ();
 FILLCELL_X4 FILLER_187_1257 ();
 FILLCELL_X2 FILLER_187_1261 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X32 FILLER_187_1584 ();
 FILLCELL_X32 FILLER_187_1616 ();
 FILLCELL_X32 FILLER_187_1648 ();
 FILLCELL_X32 FILLER_187_1680 ();
 FILLCELL_X32 FILLER_187_1712 ();
 FILLCELL_X32 FILLER_187_1744 ();
 FILLCELL_X32 FILLER_187_1776 ();
 FILLCELL_X32 FILLER_187_1808 ();
 FILLCELL_X32 FILLER_187_1840 ();
 FILLCELL_X32 FILLER_187_1872 ();
 FILLCELL_X32 FILLER_187_1904 ();
 FILLCELL_X32 FILLER_187_1936 ();
 FILLCELL_X32 FILLER_187_1968 ();
 FILLCELL_X32 FILLER_187_2000 ();
 FILLCELL_X32 FILLER_187_2032 ();
 FILLCELL_X32 FILLER_187_2064 ();
 FILLCELL_X16 FILLER_187_2096 ();
 FILLCELL_X2 FILLER_187_2112 ();
 FILLCELL_X1 FILLER_187_2114 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X32 FILLER_188_1240 ();
 FILLCELL_X32 FILLER_188_1272 ();
 FILLCELL_X32 FILLER_188_1304 ();
 FILLCELL_X32 FILLER_188_1336 ();
 FILLCELL_X32 FILLER_188_1368 ();
 FILLCELL_X32 FILLER_188_1400 ();
 FILLCELL_X32 FILLER_188_1432 ();
 FILLCELL_X32 FILLER_188_1464 ();
 FILLCELL_X32 FILLER_188_1496 ();
 FILLCELL_X32 FILLER_188_1528 ();
 FILLCELL_X32 FILLER_188_1560 ();
 FILLCELL_X32 FILLER_188_1592 ();
 FILLCELL_X32 FILLER_188_1624 ();
 FILLCELL_X32 FILLER_188_1656 ();
 FILLCELL_X32 FILLER_188_1688 ();
 FILLCELL_X32 FILLER_188_1720 ();
 FILLCELL_X32 FILLER_188_1752 ();
 FILLCELL_X32 FILLER_188_1784 ();
 FILLCELL_X32 FILLER_188_1816 ();
 FILLCELL_X32 FILLER_188_1848 ();
 FILLCELL_X8 FILLER_188_1880 ();
 FILLCELL_X4 FILLER_188_1888 ();
 FILLCELL_X2 FILLER_188_1892 ();
 FILLCELL_X32 FILLER_188_1895 ();
 FILLCELL_X32 FILLER_188_1927 ();
 FILLCELL_X32 FILLER_188_1959 ();
 FILLCELL_X32 FILLER_188_1991 ();
 FILLCELL_X32 FILLER_188_2023 ();
 FILLCELL_X32 FILLER_188_2055 ();
 FILLCELL_X16 FILLER_188_2087 ();
 FILLCELL_X8 FILLER_188_2103 ();
 FILLCELL_X4 FILLER_188_2111 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X8 FILLER_189_1249 ();
 FILLCELL_X4 FILLER_189_1257 ();
 FILLCELL_X2 FILLER_189_1261 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X32 FILLER_189_1584 ();
 FILLCELL_X32 FILLER_189_1616 ();
 FILLCELL_X32 FILLER_189_1648 ();
 FILLCELL_X32 FILLER_189_1680 ();
 FILLCELL_X32 FILLER_189_1712 ();
 FILLCELL_X32 FILLER_189_1744 ();
 FILLCELL_X32 FILLER_189_1776 ();
 FILLCELL_X32 FILLER_189_1808 ();
 FILLCELL_X32 FILLER_189_1840 ();
 FILLCELL_X32 FILLER_189_1872 ();
 FILLCELL_X32 FILLER_189_1904 ();
 FILLCELL_X32 FILLER_189_1936 ();
 FILLCELL_X32 FILLER_189_1968 ();
 FILLCELL_X32 FILLER_189_2000 ();
 FILLCELL_X32 FILLER_189_2032 ();
 FILLCELL_X32 FILLER_189_2064 ();
 FILLCELL_X16 FILLER_189_2096 ();
 FILLCELL_X2 FILLER_189_2112 ();
 FILLCELL_X1 FILLER_189_2114 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X32 FILLER_190_1240 ();
 FILLCELL_X32 FILLER_190_1272 ();
 FILLCELL_X32 FILLER_190_1304 ();
 FILLCELL_X32 FILLER_190_1336 ();
 FILLCELL_X32 FILLER_190_1368 ();
 FILLCELL_X32 FILLER_190_1400 ();
 FILLCELL_X32 FILLER_190_1432 ();
 FILLCELL_X32 FILLER_190_1464 ();
 FILLCELL_X32 FILLER_190_1496 ();
 FILLCELL_X32 FILLER_190_1528 ();
 FILLCELL_X32 FILLER_190_1560 ();
 FILLCELL_X32 FILLER_190_1592 ();
 FILLCELL_X32 FILLER_190_1624 ();
 FILLCELL_X32 FILLER_190_1656 ();
 FILLCELL_X32 FILLER_190_1688 ();
 FILLCELL_X32 FILLER_190_1720 ();
 FILLCELL_X32 FILLER_190_1752 ();
 FILLCELL_X32 FILLER_190_1784 ();
 FILLCELL_X32 FILLER_190_1816 ();
 FILLCELL_X32 FILLER_190_1848 ();
 FILLCELL_X8 FILLER_190_1880 ();
 FILLCELL_X4 FILLER_190_1888 ();
 FILLCELL_X2 FILLER_190_1892 ();
 FILLCELL_X32 FILLER_190_1895 ();
 FILLCELL_X32 FILLER_190_1927 ();
 FILLCELL_X32 FILLER_190_1959 ();
 FILLCELL_X32 FILLER_190_1991 ();
 FILLCELL_X32 FILLER_190_2023 ();
 FILLCELL_X32 FILLER_190_2055 ();
 FILLCELL_X16 FILLER_190_2087 ();
 FILLCELL_X8 FILLER_190_2103 ();
 FILLCELL_X4 FILLER_190_2111 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X32 FILLER_191_1217 ();
 FILLCELL_X8 FILLER_191_1249 ();
 FILLCELL_X4 FILLER_191_1257 ();
 FILLCELL_X2 FILLER_191_1261 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X32 FILLER_191_1584 ();
 FILLCELL_X32 FILLER_191_1616 ();
 FILLCELL_X32 FILLER_191_1648 ();
 FILLCELL_X32 FILLER_191_1680 ();
 FILLCELL_X32 FILLER_191_1712 ();
 FILLCELL_X32 FILLER_191_1744 ();
 FILLCELL_X32 FILLER_191_1776 ();
 FILLCELL_X32 FILLER_191_1808 ();
 FILLCELL_X32 FILLER_191_1840 ();
 FILLCELL_X32 FILLER_191_1872 ();
 FILLCELL_X32 FILLER_191_1904 ();
 FILLCELL_X32 FILLER_191_1936 ();
 FILLCELL_X32 FILLER_191_1968 ();
 FILLCELL_X32 FILLER_191_2000 ();
 FILLCELL_X32 FILLER_191_2032 ();
 FILLCELL_X32 FILLER_191_2064 ();
 FILLCELL_X16 FILLER_191_2096 ();
 FILLCELL_X2 FILLER_191_2112 ();
 FILLCELL_X1 FILLER_191_2114 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X32 FILLER_192_1208 ();
 FILLCELL_X32 FILLER_192_1240 ();
 FILLCELL_X32 FILLER_192_1272 ();
 FILLCELL_X32 FILLER_192_1304 ();
 FILLCELL_X32 FILLER_192_1336 ();
 FILLCELL_X32 FILLER_192_1368 ();
 FILLCELL_X32 FILLER_192_1400 ();
 FILLCELL_X32 FILLER_192_1432 ();
 FILLCELL_X32 FILLER_192_1464 ();
 FILLCELL_X32 FILLER_192_1496 ();
 FILLCELL_X32 FILLER_192_1528 ();
 FILLCELL_X32 FILLER_192_1560 ();
 FILLCELL_X32 FILLER_192_1592 ();
 FILLCELL_X32 FILLER_192_1624 ();
 FILLCELL_X32 FILLER_192_1656 ();
 FILLCELL_X32 FILLER_192_1688 ();
 FILLCELL_X32 FILLER_192_1720 ();
 FILLCELL_X32 FILLER_192_1752 ();
 FILLCELL_X32 FILLER_192_1784 ();
 FILLCELL_X32 FILLER_192_1816 ();
 FILLCELL_X32 FILLER_192_1848 ();
 FILLCELL_X8 FILLER_192_1880 ();
 FILLCELL_X4 FILLER_192_1888 ();
 FILLCELL_X2 FILLER_192_1892 ();
 FILLCELL_X32 FILLER_192_1895 ();
 FILLCELL_X32 FILLER_192_1927 ();
 FILLCELL_X32 FILLER_192_1959 ();
 FILLCELL_X32 FILLER_192_1991 ();
 FILLCELL_X32 FILLER_192_2023 ();
 FILLCELL_X32 FILLER_192_2055 ();
 FILLCELL_X16 FILLER_192_2087 ();
 FILLCELL_X8 FILLER_192_2103 ();
 FILLCELL_X4 FILLER_192_2111 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X32 FILLER_193_1584 ();
 FILLCELL_X32 FILLER_193_1616 ();
 FILLCELL_X32 FILLER_193_1648 ();
 FILLCELL_X32 FILLER_193_1680 ();
 FILLCELL_X32 FILLER_193_1712 ();
 FILLCELL_X32 FILLER_193_1744 ();
 FILLCELL_X32 FILLER_193_1776 ();
 FILLCELL_X32 FILLER_193_1808 ();
 FILLCELL_X32 FILLER_193_1840 ();
 FILLCELL_X32 FILLER_193_1872 ();
 FILLCELL_X32 FILLER_193_1904 ();
 FILLCELL_X32 FILLER_193_1936 ();
 FILLCELL_X32 FILLER_193_1968 ();
 FILLCELL_X32 FILLER_193_2000 ();
 FILLCELL_X32 FILLER_193_2032 ();
 FILLCELL_X32 FILLER_193_2064 ();
 FILLCELL_X16 FILLER_193_2096 ();
 FILLCELL_X2 FILLER_193_2112 ();
 FILLCELL_X1 FILLER_193_2114 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X32 FILLER_194_1208 ();
 FILLCELL_X32 FILLER_194_1240 ();
 FILLCELL_X32 FILLER_194_1272 ();
 FILLCELL_X32 FILLER_194_1304 ();
 FILLCELL_X32 FILLER_194_1336 ();
 FILLCELL_X32 FILLER_194_1368 ();
 FILLCELL_X32 FILLER_194_1400 ();
 FILLCELL_X32 FILLER_194_1432 ();
 FILLCELL_X32 FILLER_194_1464 ();
 FILLCELL_X32 FILLER_194_1496 ();
 FILLCELL_X32 FILLER_194_1528 ();
 FILLCELL_X32 FILLER_194_1560 ();
 FILLCELL_X32 FILLER_194_1592 ();
 FILLCELL_X32 FILLER_194_1624 ();
 FILLCELL_X32 FILLER_194_1656 ();
 FILLCELL_X32 FILLER_194_1688 ();
 FILLCELL_X32 FILLER_194_1720 ();
 FILLCELL_X32 FILLER_194_1752 ();
 FILLCELL_X32 FILLER_194_1784 ();
 FILLCELL_X32 FILLER_194_1816 ();
 FILLCELL_X32 FILLER_194_1848 ();
 FILLCELL_X8 FILLER_194_1880 ();
 FILLCELL_X4 FILLER_194_1888 ();
 FILLCELL_X2 FILLER_194_1892 ();
 FILLCELL_X32 FILLER_194_1895 ();
 FILLCELL_X32 FILLER_194_1927 ();
 FILLCELL_X32 FILLER_194_1959 ();
 FILLCELL_X32 FILLER_194_1991 ();
 FILLCELL_X32 FILLER_194_2023 ();
 FILLCELL_X32 FILLER_194_2055 ();
 FILLCELL_X16 FILLER_194_2087 ();
 FILLCELL_X8 FILLER_194_2103 ();
 FILLCELL_X4 FILLER_194_2111 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X32 FILLER_195_1217 ();
 FILLCELL_X8 FILLER_195_1249 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X32 FILLER_195_1584 ();
 FILLCELL_X32 FILLER_195_1616 ();
 FILLCELL_X32 FILLER_195_1648 ();
 FILLCELL_X32 FILLER_195_1680 ();
 FILLCELL_X32 FILLER_195_1712 ();
 FILLCELL_X32 FILLER_195_1744 ();
 FILLCELL_X32 FILLER_195_1776 ();
 FILLCELL_X32 FILLER_195_1808 ();
 FILLCELL_X32 FILLER_195_1840 ();
 FILLCELL_X32 FILLER_195_1872 ();
 FILLCELL_X32 FILLER_195_1904 ();
 FILLCELL_X32 FILLER_195_1936 ();
 FILLCELL_X32 FILLER_195_1968 ();
 FILLCELL_X32 FILLER_195_2000 ();
 FILLCELL_X32 FILLER_195_2032 ();
 FILLCELL_X32 FILLER_195_2064 ();
 FILLCELL_X16 FILLER_195_2096 ();
 FILLCELL_X2 FILLER_195_2112 ();
 FILLCELL_X1 FILLER_195_2114 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X32 FILLER_196_1272 ();
 FILLCELL_X32 FILLER_196_1304 ();
 FILLCELL_X32 FILLER_196_1336 ();
 FILLCELL_X32 FILLER_196_1368 ();
 FILLCELL_X32 FILLER_196_1400 ();
 FILLCELL_X32 FILLER_196_1432 ();
 FILLCELL_X32 FILLER_196_1464 ();
 FILLCELL_X32 FILLER_196_1496 ();
 FILLCELL_X32 FILLER_196_1528 ();
 FILLCELL_X32 FILLER_196_1560 ();
 FILLCELL_X32 FILLER_196_1592 ();
 FILLCELL_X32 FILLER_196_1624 ();
 FILLCELL_X32 FILLER_196_1656 ();
 FILLCELL_X32 FILLER_196_1688 ();
 FILLCELL_X32 FILLER_196_1720 ();
 FILLCELL_X32 FILLER_196_1752 ();
 FILLCELL_X32 FILLER_196_1784 ();
 FILLCELL_X32 FILLER_196_1816 ();
 FILLCELL_X32 FILLER_196_1848 ();
 FILLCELL_X8 FILLER_196_1880 ();
 FILLCELL_X4 FILLER_196_1888 ();
 FILLCELL_X2 FILLER_196_1892 ();
 FILLCELL_X32 FILLER_196_1895 ();
 FILLCELL_X32 FILLER_196_1927 ();
 FILLCELL_X32 FILLER_196_1959 ();
 FILLCELL_X32 FILLER_196_1991 ();
 FILLCELL_X32 FILLER_196_2023 ();
 FILLCELL_X32 FILLER_196_2055 ();
 FILLCELL_X16 FILLER_196_2087 ();
 FILLCELL_X8 FILLER_196_2103 ();
 FILLCELL_X4 FILLER_196_2111 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X32 FILLER_197_1584 ();
 FILLCELL_X32 FILLER_197_1616 ();
 FILLCELL_X32 FILLER_197_1648 ();
 FILLCELL_X32 FILLER_197_1680 ();
 FILLCELL_X32 FILLER_197_1712 ();
 FILLCELL_X32 FILLER_197_1744 ();
 FILLCELL_X32 FILLER_197_1776 ();
 FILLCELL_X32 FILLER_197_1808 ();
 FILLCELL_X32 FILLER_197_1840 ();
 FILLCELL_X32 FILLER_197_1872 ();
 FILLCELL_X32 FILLER_197_1904 ();
 FILLCELL_X32 FILLER_197_1936 ();
 FILLCELL_X32 FILLER_197_1968 ();
 FILLCELL_X32 FILLER_197_2000 ();
 FILLCELL_X32 FILLER_197_2032 ();
 FILLCELL_X32 FILLER_197_2064 ();
 FILLCELL_X16 FILLER_197_2096 ();
 FILLCELL_X2 FILLER_197_2112 ();
 FILLCELL_X1 FILLER_197_2114 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X32 FILLER_198_1208 ();
 FILLCELL_X32 FILLER_198_1240 ();
 FILLCELL_X32 FILLER_198_1272 ();
 FILLCELL_X32 FILLER_198_1304 ();
 FILLCELL_X32 FILLER_198_1336 ();
 FILLCELL_X32 FILLER_198_1368 ();
 FILLCELL_X32 FILLER_198_1400 ();
 FILLCELL_X32 FILLER_198_1432 ();
 FILLCELL_X32 FILLER_198_1464 ();
 FILLCELL_X32 FILLER_198_1496 ();
 FILLCELL_X32 FILLER_198_1528 ();
 FILLCELL_X32 FILLER_198_1560 ();
 FILLCELL_X32 FILLER_198_1592 ();
 FILLCELL_X32 FILLER_198_1624 ();
 FILLCELL_X32 FILLER_198_1656 ();
 FILLCELL_X32 FILLER_198_1688 ();
 FILLCELL_X32 FILLER_198_1720 ();
 FILLCELL_X32 FILLER_198_1752 ();
 FILLCELL_X32 FILLER_198_1784 ();
 FILLCELL_X32 FILLER_198_1816 ();
 FILLCELL_X32 FILLER_198_1848 ();
 FILLCELL_X8 FILLER_198_1880 ();
 FILLCELL_X4 FILLER_198_1888 ();
 FILLCELL_X2 FILLER_198_1892 ();
 FILLCELL_X32 FILLER_198_1895 ();
 FILLCELL_X32 FILLER_198_1927 ();
 FILLCELL_X32 FILLER_198_1959 ();
 FILLCELL_X32 FILLER_198_1991 ();
 FILLCELL_X32 FILLER_198_2023 ();
 FILLCELL_X32 FILLER_198_2055 ();
 FILLCELL_X16 FILLER_198_2087 ();
 FILLCELL_X8 FILLER_198_2103 ();
 FILLCELL_X4 FILLER_198_2111 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X32 FILLER_199_1584 ();
 FILLCELL_X32 FILLER_199_1616 ();
 FILLCELL_X32 FILLER_199_1648 ();
 FILLCELL_X32 FILLER_199_1680 ();
 FILLCELL_X32 FILLER_199_1712 ();
 FILLCELL_X32 FILLER_199_1744 ();
 FILLCELL_X32 FILLER_199_1776 ();
 FILLCELL_X32 FILLER_199_1808 ();
 FILLCELL_X32 FILLER_199_1840 ();
 FILLCELL_X32 FILLER_199_1872 ();
 FILLCELL_X32 FILLER_199_1904 ();
 FILLCELL_X32 FILLER_199_1936 ();
 FILLCELL_X32 FILLER_199_1968 ();
 FILLCELL_X32 FILLER_199_2000 ();
 FILLCELL_X32 FILLER_199_2032 ();
 FILLCELL_X32 FILLER_199_2064 ();
 FILLCELL_X16 FILLER_199_2096 ();
 FILLCELL_X2 FILLER_199_2112 ();
 FILLCELL_X1 FILLER_199_2114 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X32 FILLER_200_1304 ();
 FILLCELL_X32 FILLER_200_1336 ();
 FILLCELL_X32 FILLER_200_1368 ();
 FILLCELL_X32 FILLER_200_1400 ();
 FILLCELL_X32 FILLER_200_1432 ();
 FILLCELL_X32 FILLER_200_1464 ();
 FILLCELL_X32 FILLER_200_1496 ();
 FILLCELL_X32 FILLER_200_1528 ();
 FILLCELL_X32 FILLER_200_1560 ();
 FILLCELL_X32 FILLER_200_1592 ();
 FILLCELL_X32 FILLER_200_1624 ();
 FILLCELL_X32 FILLER_200_1656 ();
 FILLCELL_X32 FILLER_200_1688 ();
 FILLCELL_X32 FILLER_200_1720 ();
 FILLCELL_X32 FILLER_200_1752 ();
 FILLCELL_X32 FILLER_200_1784 ();
 FILLCELL_X32 FILLER_200_1816 ();
 FILLCELL_X32 FILLER_200_1848 ();
 FILLCELL_X8 FILLER_200_1880 ();
 FILLCELL_X4 FILLER_200_1888 ();
 FILLCELL_X2 FILLER_200_1892 ();
 FILLCELL_X32 FILLER_200_1895 ();
 FILLCELL_X32 FILLER_200_1927 ();
 FILLCELL_X32 FILLER_200_1959 ();
 FILLCELL_X32 FILLER_200_1991 ();
 FILLCELL_X32 FILLER_200_2023 ();
 FILLCELL_X32 FILLER_200_2055 ();
 FILLCELL_X16 FILLER_200_2087 ();
 FILLCELL_X8 FILLER_200_2103 ();
 FILLCELL_X4 FILLER_200_2111 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X32 FILLER_201_1648 ();
 FILLCELL_X32 FILLER_201_1680 ();
 FILLCELL_X32 FILLER_201_1712 ();
 FILLCELL_X32 FILLER_201_1744 ();
 FILLCELL_X32 FILLER_201_1776 ();
 FILLCELL_X32 FILLER_201_1808 ();
 FILLCELL_X32 FILLER_201_1840 ();
 FILLCELL_X32 FILLER_201_1872 ();
 FILLCELL_X32 FILLER_201_1904 ();
 FILLCELL_X32 FILLER_201_1936 ();
 FILLCELL_X32 FILLER_201_1968 ();
 FILLCELL_X32 FILLER_201_2000 ();
 FILLCELL_X32 FILLER_201_2032 ();
 FILLCELL_X32 FILLER_201_2064 ();
 FILLCELL_X16 FILLER_201_2096 ();
 FILLCELL_X2 FILLER_201_2112 ();
 FILLCELL_X1 FILLER_201_2114 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X32 FILLER_202_1592 ();
 FILLCELL_X32 FILLER_202_1624 ();
 FILLCELL_X32 FILLER_202_1656 ();
 FILLCELL_X32 FILLER_202_1688 ();
 FILLCELL_X32 FILLER_202_1720 ();
 FILLCELL_X32 FILLER_202_1752 ();
 FILLCELL_X32 FILLER_202_1784 ();
 FILLCELL_X32 FILLER_202_1816 ();
 FILLCELL_X32 FILLER_202_1848 ();
 FILLCELL_X8 FILLER_202_1880 ();
 FILLCELL_X4 FILLER_202_1888 ();
 FILLCELL_X2 FILLER_202_1892 ();
 FILLCELL_X32 FILLER_202_1895 ();
 FILLCELL_X32 FILLER_202_1927 ();
 FILLCELL_X32 FILLER_202_1959 ();
 FILLCELL_X32 FILLER_202_1991 ();
 FILLCELL_X32 FILLER_202_2023 ();
 FILLCELL_X32 FILLER_202_2055 ();
 FILLCELL_X16 FILLER_202_2087 ();
 FILLCELL_X8 FILLER_202_2103 ();
 FILLCELL_X4 FILLER_202_2111 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X32 FILLER_203_1648 ();
 FILLCELL_X32 FILLER_203_1680 ();
 FILLCELL_X32 FILLER_203_1712 ();
 FILLCELL_X32 FILLER_203_1744 ();
 FILLCELL_X32 FILLER_203_1776 ();
 FILLCELL_X32 FILLER_203_1808 ();
 FILLCELL_X32 FILLER_203_1840 ();
 FILLCELL_X32 FILLER_203_1872 ();
 FILLCELL_X32 FILLER_203_1904 ();
 FILLCELL_X32 FILLER_203_1936 ();
 FILLCELL_X32 FILLER_203_1968 ();
 FILLCELL_X32 FILLER_203_2000 ();
 FILLCELL_X32 FILLER_203_2032 ();
 FILLCELL_X32 FILLER_203_2064 ();
 FILLCELL_X16 FILLER_203_2096 ();
 FILLCELL_X2 FILLER_203_2112 ();
 FILLCELL_X1 FILLER_203_2114 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X32 FILLER_204_1592 ();
 FILLCELL_X32 FILLER_204_1624 ();
 FILLCELL_X32 FILLER_204_1656 ();
 FILLCELL_X32 FILLER_204_1688 ();
 FILLCELL_X32 FILLER_204_1720 ();
 FILLCELL_X32 FILLER_204_1752 ();
 FILLCELL_X32 FILLER_204_1784 ();
 FILLCELL_X32 FILLER_204_1816 ();
 FILLCELL_X32 FILLER_204_1848 ();
 FILLCELL_X8 FILLER_204_1880 ();
 FILLCELL_X4 FILLER_204_1888 ();
 FILLCELL_X2 FILLER_204_1892 ();
 FILLCELL_X32 FILLER_204_1895 ();
 FILLCELL_X32 FILLER_204_1927 ();
 FILLCELL_X32 FILLER_204_1959 ();
 FILLCELL_X32 FILLER_204_1991 ();
 FILLCELL_X32 FILLER_204_2023 ();
 FILLCELL_X32 FILLER_204_2055 ();
 FILLCELL_X16 FILLER_204_2087 ();
 FILLCELL_X8 FILLER_204_2103 ();
 FILLCELL_X4 FILLER_204_2111 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X32 FILLER_205_1648 ();
 FILLCELL_X32 FILLER_205_1680 ();
 FILLCELL_X32 FILLER_205_1712 ();
 FILLCELL_X32 FILLER_205_1744 ();
 FILLCELL_X32 FILLER_205_1776 ();
 FILLCELL_X32 FILLER_205_1808 ();
 FILLCELL_X32 FILLER_205_1840 ();
 FILLCELL_X32 FILLER_205_1872 ();
 FILLCELL_X32 FILLER_205_1904 ();
 FILLCELL_X32 FILLER_205_1936 ();
 FILLCELL_X32 FILLER_205_1968 ();
 FILLCELL_X32 FILLER_205_2000 ();
 FILLCELL_X32 FILLER_205_2032 ();
 FILLCELL_X32 FILLER_205_2064 ();
 FILLCELL_X16 FILLER_205_2096 ();
 FILLCELL_X2 FILLER_205_2112 ();
 FILLCELL_X1 FILLER_205_2114 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X32 FILLER_206_1592 ();
 FILLCELL_X32 FILLER_206_1624 ();
 FILLCELL_X32 FILLER_206_1656 ();
 FILLCELL_X32 FILLER_206_1688 ();
 FILLCELL_X32 FILLER_206_1720 ();
 FILLCELL_X32 FILLER_206_1752 ();
 FILLCELL_X32 FILLER_206_1784 ();
 FILLCELL_X32 FILLER_206_1816 ();
 FILLCELL_X32 FILLER_206_1848 ();
 FILLCELL_X8 FILLER_206_1880 ();
 FILLCELL_X4 FILLER_206_1888 ();
 FILLCELL_X2 FILLER_206_1892 ();
 FILLCELL_X32 FILLER_206_1895 ();
 FILLCELL_X32 FILLER_206_1927 ();
 FILLCELL_X32 FILLER_206_1959 ();
 FILLCELL_X32 FILLER_206_1991 ();
 FILLCELL_X32 FILLER_206_2023 ();
 FILLCELL_X32 FILLER_206_2055 ();
 FILLCELL_X16 FILLER_206_2087 ();
 FILLCELL_X8 FILLER_206_2103 ();
 FILLCELL_X4 FILLER_206_2111 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X32 FILLER_207_1648 ();
 FILLCELL_X32 FILLER_207_1680 ();
 FILLCELL_X32 FILLER_207_1712 ();
 FILLCELL_X32 FILLER_207_1744 ();
 FILLCELL_X32 FILLER_207_1776 ();
 FILLCELL_X32 FILLER_207_1808 ();
 FILLCELL_X32 FILLER_207_1840 ();
 FILLCELL_X32 FILLER_207_1872 ();
 FILLCELL_X32 FILLER_207_1904 ();
 FILLCELL_X32 FILLER_207_1936 ();
 FILLCELL_X32 FILLER_207_1968 ();
 FILLCELL_X32 FILLER_207_2000 ();
 FILLCELL_X32 FILLER_207_2032 ();
 FILLCELL_X32 FILLER_207_2064 ();
 FILLCELL_X16 FILLER_207_2096 ();
 FILLCELL_X2 FILLER_207_2112 ();
 FILLCELL_X1 FILLER_207_2114 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X32 FILLER_208_1592 ();
 FILLCELL_X32 FILLER_208_1624 ();
 FILLCELL_X32 FILLER_208_1656 ();
 FILLCELL_X32 FILLER_208_1688 ();
 FILLCELL_X32 FILLER_208_1720 ();
 FILLCELL_X32 FILLER_208_1752 ();
 FILLCELL_X32 FILLER_208_1784 ();
 FILLCELL_X32 FILLER_208_1816 ();
 FILLCELL_X32 FILLER_208_1848 ();
 FILLCELL_X8 FILLER_208_1880 ();
 FILLCELL_X4 FILLER_208_1888 ();
 FILLCELL_X2 FILLER_208_1892 ();
 FILLCELL_X32 FILLER_208_1895 ();
 FILLCELL_X32 FILLER_208_1927 ();
 FILLCELL_X32 FILLER_208_1959 ();
 FILLCELL_X32 FILLER_208_1991 ();
 FILLCELL_X32 FILLER_208_2023 ();
 FILLCELL_X32 FILLER_208_2055 ();
 FILLCELL_X16 FILLER_208_2087 ();
 FILLCELL_X8 FILLER_208_2103 ();
 FILLCELL_X4 FILLER_208_2111 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X32 FILLER_209_1744 ();
 FILLCELL_X32 FILLER_209_1776 ();
 FILLCELL_X32 FILLER_209_1808 ();
 FILLCELL_X32 FILLER_209_1840 ();
 FILLCELL_X32 FILLER_209_1872 ();
 FILLCELL_X32 FILLER_209_1904 ();
 FILLCELL_X32 FILLER_209_1936 ();
 FILLCELL_X32 FILLER_209_1968 ();
 FILLCELL_X32 FILLER_209_2000 ();
 FILLCELL_X32 FILLER_209_2032 ();
 FILLCELL_X32 FILLER_209_2064 ();
 FILLCELL_X16 FILLER_209_2096 ();
 FILLCELL_X2 FILLER_209_2112 ();
 FILLCELL_X1 FILLER_209_2114 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X32 FILLER_210_1752 ();
 FILLCELL_X32 FILLER_210_1784 ();
 FILLCELL_X32 FILLER_210_1816 ();
 FILLCELL_X32 FILLER_210_1848 ();
 FILLCELL_X8 FILLER_210_1880 ();
 FILLCELL_X4 FILLER_210_1888 ();
 FILLCELL_X2 FILLER_210_1892 ();
 FILLCELL_X32 FILLER_210_1895 ();
 FILLCELL_X32 FILLER_210_1927 ();
 FILLCELL_X32 FILLER_210_1959 ();
 FILLCELL_X32 FILLER_210_1991 ();
 FILLCELL_X32 FILLER_210_2023 ();
 FILLCELL_X32 FILLER_210_2055 ();
 FILLCELL_X16 FILLER_210_2087 ();
 FILLCELL_X8 FILLER_210_2103 ();
 FILLCELL_X4 FILLER_210_2111 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X32 FILLER_211_1744 ();
 FILLCELL_X32 FILLER_211_1776 ();
 FILLCELL_X32 FILLER_211_1808 ();
 FILLCELL_X32 FILLER_211_1840 ();
 FILLCELL_X32 FILLER_211_1872 ();
 FILLCELL_X32 FILLER_211_1904 ();
 FILLCELL_X32 FILLER_211_1936 ();
 FILLCELL_X32 FILLER_211_1968 ();
 FILLCELL_X32 FILLER_211_2000 ();
 FILLCELL_X32 FILLER_211_2032 ();
 FILLCELL_X32 FILLER_211_2064 ();
 FILLCELL_X16 FILLER_211_2096 ();
 FILLCELL_X2 FILLER_211_2112 ();
 FILLCELL_X1 FILLER_211_2114 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X32 FILLER_212_1752 ();
 FILLCELL_X32 FILLER_212_1784 ();
 FILLCELL_X32 FILLER_212_1816 ();
 FILLCELL_X32 FILLER_212_1848 ();
 FILLCELL_X8 FILLER_212_1880 ();
 FILLCELL_X4 FILLER_212_1888 ();
 FILLCELL_X2 FILLER_212_1892 ();
 FILLCELL_X32 FILLER_212_1895 ();
 FILLCELL_X32 FILLER_212_1927 ();
 FILLCELL_X32 FILLER_212_1959 ();
 FILLCELL_X32 FILLER_212_1991 ();
 FILLCELL_X32 FILLER_212_2023 ();
 FILLCELL_X32 FILLER_212_2055 ();
 FILLCELL_X16 FILLER_212_2087 ();
 FILLCELL_X8 FILLER_212_2103 ();
 FILLCELL_X4 FILLER_212_2111 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X32 FILLER_213_1744 ();
 FILLCELL_X32 FILLER_213_1776 ();
 FILLCELL_X32 FILLER_213_1808 ();
 FILLCELL_X32 FILLER_213_1840 ();
 FILLCELL_X32 FILLER_213_1872 ();
 FILLCELL_X32 FILLER_213_1904 ();
 FILLCELL_X32 FILLER_213_1936 ();
 FILLCELL_X32 FILLER_213_1968 ();
 FILLCELL_X32 FILLER_213_2000 ();
 FILLCELL_X32 FILLER_213_2032 ();
 FILLCELL_X32 FILLER_213_2064 ();
 FILLCELL_X16 FILLER_213_2096 ();
 FILLCELL_X2 FILLER_213_2112 ();
 FILLCELL_X1 FILLER_213_2114 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X32 FILLER_214_1752 ();
 FILLCELL_X32 FILLER_214_1784 ();
 FILLCELL_X32 FILLER_214_1816 ();
 FILLCELL_X32 FILLER_214_1848 ();
 FILLCELL_X8 FILLER_214_1880 ();
 FILLCELL_X4 FILLER_214_1888 ();
 FILLCELL_X2 FILLER_214_1892 ();
 FILLCELL_X32 FILLER_214_1895 ();
 FILLCELL_X32 FILLER_214_1927 ();
 FILLCELL_X32 FILLER_214_1959 ();
 FILLCELL_X32 FILLER_214_1991 ();
 FILLCELL_X32 FILLER_214_2023 ();
 FILLCELL_X32 FILLER_214_2055 ();
 FILLCELL_X16 FILLER_214_2087 ();
 FILLCELL_X8 FILLER_214_2103 ();
 FILLCELL_X4 FILLER_214_2111 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X32 FILLER_215_1744 ();
 FILLCELL_X32 FILLER_215_1776 ();
 FILLCELL_X32 FILLER_215_1808 ();
 FILLCELL_X32 FILLER_215_1840 ();
 FILLCELL_X32 FILLER_215_1872 ();
 FILLCELL_X32 FILLER_215_1904 ();
 FILLCELL_X32 FILLER_215_1936 ();
 FILLCELL_X32 FILLER_215_1968 ();
 FILLCELL_X32 FILLER_215_2000 ();
 FILLCELL_X32 FILLER_215_2032 ();
 FILLCELL_X32 FILLER_215_2064 ();
 FILLCELL_X16 FILLER_215_2096 ();
 FILLCELL_X2 FILLER_215_2112 ();
 FILLCELL_X1 FILLER_215_2114 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X32 FILLER_216_1752 ();
 FILLCELL_X32 FILLER_216_1784 ();
 FILLCELL_X32 FILLER_216_1816 ();
 FILLCELL_X32 FILLER_216_1848 ();
 FILLCELL_X8 FILLER_216_1880 ();
 FILLCELL_X4 FILLER_216_1888 ();
 FILLCELL_X2 FILLER_216_1892 ();
 FILLCELL_X32 FILLER_216_1895 ();
 FILLCELL_X32 FILLER_216_1927 ();
 FILLCELL_X32 FILLER_216_1959 ();
 FILLCELL_X32 FILLER_216_1991 ();
 FILLCELL_X32 FILLER_216_2023 ();
 FILLCELL_X32 FILLER_216_2055 ();
 FILLCELL_X16 FILLER_216_2087 ();
 FILLCELL_X8 FILLER_216_2103 ();
 FILLCELL_X4 FILLER_216_2111 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X32 FILLER_217_1744 ();
 FILLCELL_X32 FILLER_217_1776 ();
 FILLCELL_X32 FILLER_217_1808 ();
 FILLCELL_X32 FILLER_217_1840 ();
 FILLCELL_X32 FILLER_217_1872 ();
 FILLCELL_X32 FILLER_217_1904 ();
 FILLCELL_X32 FILLER_217_1936 ();
 FILLCELL_X32 FILLER_217_1968 ();
 FILLCELL_X32 FILLER_217_2000 ();
 FILLCELL_X32 FILLER_217_2032 ();
 FILLCELL_X32 FILLER_217_2064 ();
 FILLCELL_X16 FILLER_217_2096 ();
 FILLCELL_X2 FILLER_217_2112 ();
 FILLCELL_X1 FILLER_217_2114 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X32 FILLER_218_1752 ();
 FILLCELL_X32 FILLER_218_1784 ();
 FILLCELL_X32 FILLER_218_1816 ();
 FILLCELL_X32 FILLER_218_1848 ();
 FILLCELL_X8 FILLER_218_1880 ();
 FILLCELL_X4 FILLER_218_1888 ();
 FILLCELL_X2 FILLER_218_1892 ();
 FILLCELL_X32 FILLER_218_1895 ();
 FILLCELL_X32 FILLER_218_1927 ();
 FILLCELL_X32 FILLER_218_1959 ();
 FILLCELL_X32 FILLER_218_1991 ();
 FILLCELL_X32 FILLER_218_2023 ();
 FILLCELL_X32 FILLER_218_2055 ();
 FILLCELL_X16 FILLER_218_2087 ();
 FILLCELL_X8 FILLER_218_2103 ();
 FILLCELL_X4 FILLER_218_2111 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X32 FILLER_219_1744 ();
 FILLCELL_X32 FILLER_219_1776 ();
 FILLCELL_X32 FILLER_219_1808 ();
 FILLCELL_X32 FILLER_219_1840 ();
 FILLCELL_X32 FILLER_219_1872 ();
 FILLCELL_X32 FILLER_219_1904 ();
 FILLCELL_X32 FILLER_219_1936 ();
 FILLCELL_X32 FILLER_219_1968 ();
 FILLCELL_X32 FILLER_219_2000 ();
 FILLCELL_X32 FILLER_219_2032 ();
 FILLCELL_X32 FILLER_219_2064 ();
 FILLCELL_X16 FILLER_219_2096 ();
 FILLCELL_X2 FILLER_219_2112 ();
 FILLCELL_X1 FILLER_219_2114 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X32 FILLER_220_1752 ();
 FILLCELL_X32 FILLER_220_1784 ();
 FILLCELL_X32 FILLER_220_1816 ();
 FILLCELL_X32 FILLER_220_1848 ();
 FILLCELL_X8 FILLER_220_1880 ();
 FILLCELL_X4 FILLER_220_1888 ();
 FILLCELL_X2 FILLER_220_1892 ();
 FILLCELL_X32 FILLER_220_1895 ();
 FILLCELL_X32 FILLER_220_1927 ();
 FILLCELL_X32 FILLER_220_1959 ();
 FILLCELL_X32 FILLER_220_1991 ();
 FILLCELL_X32 FILLER_220_2023 ();
 FILLCELL_X32 FILLER_220_2055 ();
 FILLCELL_X16 FILLER_220_2087 ();
 FILLCELL_X8 FILLER_220_2103 ();
 FILLCELL_X4 FILLER_220_2111 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X32 FILLER_221_1744 ();
 FILLCELL_X32 FILLER_221_1776 ();
 FILLCELL_X32 FILLER_221_1808 ();
 FILLCELL_X32 FILLER_221_1840 ();
 FILLCELL_X32 FILLER_221_1872 ();
 FILLCELL_X32 FILLER_221_1904 ();
 FILLCELL_X32 FILLER_221_1936 ();
 FILLCELL_X32 FILLER_221_1968 ();
 FILLCELL_X32 FILLER_221_2000 ();
 FILLCELL_X32 FILLER_221_2032 ();
 FILLCELL_X32 FILLER_221_2064 ();
 FILLCELL_X16 FILLER_221_2096 ();
 FILLCELL_X2 FILLER_221_2112 ();
 FILLCELL_X1 FILLER_221_2114 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X32 FILLER_222_1720 ();
 FILLCELL_X32 FILLER_222_1752 ();
 FILLCELL_X32 FILLER_222_1784 ();
 FILLCELL_X32 FILLER_222_1816 ();
 FILLCELL_X32 FILLER_222_1848 ();
 FILLCELL_X8 FILLER_222_1880 ();
 FILLCELL_X4 FILLER_222_1888 ();
 FILLCELL_X2 FILLER_222_1892 ();
 FILLCELL_X32 FILLER_222_1895 ();
 FILLCELL_X32 FILLER_222_1927 ();
 FILLCELL_X32 FILLER_222_1959 ();
 FILLCELL_X32 FILLER_222_1991 ();
 FILLCELL_X32 FILLER_222_2023 ();
 FILLCELL_X32 FILLER_222_2055 ();
 FILLCELL_X16 FILLER_222_2087 ();
 FILLCELL_X8 FILLER_222_2103 ();
 FILLCELL_X4 FILLER_222_2111 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X32 FILLER_223_1744 ();
 FILLCELL_X32 FILLER_223_1776 ();
 FILLCELL_X32 FILLER_223_1808 ();
 FILLCELL_X32 FILLER_223_1840 ();
 FILLCELL_X32 FILLER_223_1872 ();
 FILLCELL_X32 FILLER_223_1904 ();
 FILLCELL_X32 FILLER_223_1936 ();
 FILLCELL_X32 FILLER_223_1968 ();
 FILLCELL_X32 FILLER_223_2000 ();
 FILLCELL_X32 FILLER_223_2032 ();
 FILLCELL_X32 FILLER_223_2064 ();
 FILLCELL_X16 FILLER_223_2096 ();
 FILLCELL_X2 FILLER_223_2112 ();
 FILLCELL_X1 FILLER_223_2114 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X32 FILLER_224_1752 ();
 FILLCELL_X32 FILLER_224_1784 ();
 FILLCELL_X32 FILLER_224_1816 ();
 FILLCELL_X32 FILLER_224_1848 ();
 FILLCELL_X8 FILLER_224_1880 ();
 FILLCELL_X4 FILLER_224_1888 ();
 FILLCELL_X2 FILLER_224_1892 ();
 FILLCELL_X32 FILLER_224_1895 ();
 FILLCELL_X32 FILLER_224_1927 ();
 FILLCELL_X32 FILLER_224_1959 ();
 FILLCELL_X32 FILLER_224_1991 ();
 FILLCELL_X32 FILLER_224_2023 ();
 FILLCELL_X32 FILLER_224_2055 ();
 FILLCELL_X16 FILLER_224_2087 ();
 FILLCELL_X8 FILLER_224_2103 ();
 FILLCELL_X4 FILLER_224_2111 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X32 FILLER_225_1744 ();
 FILLCELL_X32 FILLER_225_1776 ();
 FILLCELL_X32 FILLER_225_1808 ();
 FILLCELL_X32 FILLER_225_1840 ();
 FILLCELL_X32 FILLER_225_1872 ();
 FILLCELL_X32 FILLER_225_1904 ();
 FILLCELL_X32 FILLER_225_1936 ();
 FILLCELL_X32 FILLER_225_1968 ();
 FILLCELL_X32 FILLER_225_2000 ();
 FILLCELL_X32 FILLER_225_2032 ();
 FILLCELL_X32 FILLER_225_2064 ();
 FILLCELL_X16 FILLER_225_2096 ();
 FILLCELL_X2 FILLER_225_2112 ();
 FILLCELL_X1 FILLER_225_2114 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X32 FILLER_226_1752 ();
 FILLCELL_X32 FILLER_226_1784 ();
 FILLCELL_X32 FILLER_226_1816 ();
 FILLCELL_X32 FILLER_226_1848 ();
 FILLCELL_X8 FILLER_226_1880 ();
 FILLCELL_X4 FILLER_226_1888 ();
 FILLCELL_X2 FILLER_226_1892 ();
 FILLCELL_X32 FILLER_226_1895 ();
 FILLCELL_X32 FILLER_226_1927 ();
 FILLCELL_X32 FILLER_226_1959 ();
 FILLCELL_X32 FILLER_226_1991 ();
 FILLCELL_X32 FILLER_226_2023 ();
 FILLCELL_X32 FILLER_226_2055 ();
 FILLCELL_X16 FILLER_226_2087 ();
 FILLCELL_X8 FILLER_226_2103 ();
 FILLCELL_X4 FILLER_226_2111 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X32 FILLER_227_1744 ();
 FILLCELL_X32 FILLER_227_1776 ();
 FILLCELL_X32 FILLER_227_1808 ();
 FILLCELL_X32 FILLER_227_1840 ();
 FILLCELL_X32 FILLER_227_1872 ();
 FILLCELL_X32 FILLER_227_1904 ();
 FILLCELL_X32 FILLER_227_1936 ();
 FILLCELL_X32 FILLER_227_1968 ();
 FILLCELL_X32 FILLER_227_2000 ();
 FILLCELL_X32 FILLER_227_2032 ();
 FILLCELL_X32 FILLER_227_2064 ();
 FILLCELL_X16 FILLER_227_2096 ();
 FILLCELL_X2 FILLER_227_2112 ();
 FILLCELL_X1 FILLER_227_2114 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X32 FILLER_228_1752 ();
 FILLCELL_X32 FILLER_228_1784 ();
 FILLCELL_X32 FILLER_228_1816 ();
 FILLCELL_X32 FILLER_228_1848 ();
 FILLCELL_X8 FILLER_228_1880 ();
 FILLCELL_X4 FILLER_228_1888 ();
 FILLCELL_X2 FILLER_228_1892 ();
 FILLCELL_X32 FILLER_228_1895 ();
 FILLCELL_X32 FILLER_228_1927 ();
 FILLCELL_X32 FILLER_228_1959 ();
 FILLCELL_X32 FILLER_228_1991 ();
 FILLCELL_X32 FILLER_228_2023 ();
 FILLCELL_X32 FILLER_228_2055 ();
 FILLCELL_X16 FILLER_228_2087 ();
 FILLCELL_X8 FILLER_228_2103 ();
 FILLCELL_X4 FILLER_228_2111 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X32 FILLER_229_1744 ();
 FILLCELL_X32 FILLER_229_1776 ();
 FILLCELL_X32 FILLER_229_1808 ();
 FILLCELL_X32 FILLER_229_1840 ();
 FILLCELL_X32 FILLER_229_1872 ();
 FILLCELL_X32 FILLER_229_1904 ();
 FILLCELL_X32 FILLER_229_1936 ();
 FILLCELL_X32 FILLER_229_1968 ();
 FILLCELL_X32 FILLER_229_2000 ();
 FILLCELL_X32 FILLER_229_2032 ();
 FILLCELL_X32 FILLER_229_2064 ();
 FILLCELL_X16 FILLER_229_2096 ();
 FILLCELL_X2 FILLER_229_2112 ();
 FILLCELL_X1 FILLER_229_2114 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X32 FILLER_230_1752 ();
 FILLCELL_X32 FILLER_230_1784 ();
 FILLCELL_X32 FILLER_230_1816 ();
 FILLCELL_X32 FILLER_230_1848 ();
 FILLCELL_X8 FILLER_230_1880 ();
 FILLCELL_X4 FILLER_230_1888 ();
 FILLCELL_X2 FILLER_230_1892 ();
 FILLCELL_X32 FILLER_230_1895 ();
 FILLCELL_X32 FILLER_230_1927 ();
 FILLCELL_X32 FILLER_230_1959 ();
 FILLCELL_X32 FILLER_230_1991 ();
 FILLCELL_X32 FILLER_230_2023 ();
 FILLCELL_X32 FILLER_230_2055 ();
 FILLCELL_X16 FILLER_230_2087 ();
 FILLCELL_X8 FILLER_230_2103 ();
 FILLCELL_X4 FILLER_230_2111 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X32 FILLER_231_1744 ();
 FILLCELL_X32 FILLER_231_1776 ();
 FILLCELL_X32 FILLER_231_1808 ();
 FILLCELL_X32 FILLER_231_1840 ();
 FILLCELL_X32 FILLER_231_1872 ();
 FILLCELL_X32 FILLER_231_1904 ();
 FILLCELL_X32 FILLER_231_1936 ();
 FILLCELL_X32 FILLER_231_1968 ();
 FILLCELL_X32 FILLER_231_2000 ();
 FILLCELL_X32 FILLER_231_2032 ();
 FILLCELL_X32 FILLER_231_2064 ();
 FILLCELL_X16 FILLER_231_2096 ();
 FILLCELL_X2 FILLER_231_2112 ();
 FILLCELL_X1 FILLER_231_2114 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X32 FILLER_232_1720 ();
 FILLCELL_X32 FILLER_232_1752 ();
 FILLCELL_X32 FILLER_232_1784 ();
 FILLCELL_X32 FILLER_232_1816 ();
 FILLCELL_X32 FILLER_232_1848 ();
 FILLCELL_X8 FILLER_232_1880 ();
 FILLCELL_X4 FILLER_232_1888 ();
 FILLCELL_X2 FILLER_232_1892 ();
 FILLCELL_X32 FILLER_232_1895 ();
 FILLCELL_X32 FILLER_232_1927 ();
 FILLCELL_X32 FILLER_232_1959 ();
 FILLCELL_X32 FILLER_232_1991 ();
 FILLCELL_X32 FILLER_232_2023 ();
 FILLCELL_X32 FILLER_232_2055 ();
 FILLCELL_X16 FILLER_232_2087 ();
 FILLCELL_X8 FILLER_232_2103 ();
 FILLCELL_X4 FILLER_232_2111 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X32 FILLER_233_1744 ();
 FILLCELL_X32 FILLER_233_1776 ();
 FILLCELL_X32 FILLER_233_1808 ();
 FILLCELL_X32 FILLER_233_1840 ();
 FILLCELL_X32 FILLER_233_1872 ();
 FILLCELL_X32 FILLER_233_1904 ();
 FILLCELL_X32 FILLER_233_1936 ();
 FILLCELL_X32 FILLER_233_1968 ();
 FILLCELL_X32 FILLER_233_2000 ();
 FILLCELL_X32 FILLER_233_2032 ();
 FILLCELL_X32 FILLER_233_2064 ();
 FILLCELL_X16 FILLER_233_2096 ();
 FILLCELL_X2 FILLER_233_2112 ();
 FILLCELL_X1 FILLER_233_2114 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X32 FILLER_234_1752 ();
 FILLCELL_X32 FILLER_234_1784 ();
 FILLCELL_X32 FILLER_234_1816 ();
 FILLCELL_X32 FILLER_234_1848 ();
 FILLCELL_X8 FILLER_234_1880 ();
 FILLCELL_X4 FILLER_234_1888 ();
 FILLCELL_X2 FILLER_234_1892 ();
 FILLCELL_X32 FILLER_234_1895 ();
 FILLCELL_X32 FILLER_234_1927 ();
 FILLCELL_X32 FILLER_234_1959 ();
 FILLCELL_X32 FILLER_234_1991 ();
 FILLCELL_X32 FILLER_234_2023 ();
 FILLCELL_X32 FILLER_234_2055 ();
 FILLCELL_X16 FILLER_234_2087 ();
 FILLCELL_X8 FILLER_234_2103 ();
 FILLCELL_X4 FILLER_234_2111 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X32 FILLER_235_1744 ();
 FILLCELL_X32 FILLER_235_1776 ();
 FILLCELL_X32 FILLER_235_1808 ();
 FILLCELL_X32 FILLER_235_1840 ();
 FILLCELL_X32 FILLER_235_1872 ();
 FILLCELL_X32 FILLER_235_1904 ();
 FILLCELL_X32 FILLER_235_1936 ();
 FILLCELL_X32 FILLER_235_1968 ();
 FILLCELL_X32 FILLER_235_2000 ();
 FILLCELL_X32 FILLER_235_2032 ();
 FILLCELL_X32 FILLER_235_2064 ();
 FILLCELL_X16 FILLER_235_2096 ();
 FILLCELL_X2 FILLER_235_2112 ();
 FILLCELL_X1 FILLER_235_2114 ();
 FILLCELL_X32 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_33 ();
 FILLCELL_X32 FILLER_236_65 ();
 FILLCELL_X32 FILLER_236_97 ();
 FILLCELL_X32 FILLER_236_129 ();
 FILLCELL_X32 FILLER_236_161 ();
 FILLCELL_X32 FILLER_236_193 ();
 FILLCELL_X32 FILLER_236_225 ();
 FILLCELL_X32 FILLER_236_257 ();
 FILLCELL_X32 FILLER_236_289 ();
 FILLCELL_X32 FILLER_236_321 ();
 FILLCELL_X32 FILLER_236_353 ();
 FILLCELL_X32 FILLER_236_385 ();
 FILLCELL_X32 FILLER_236_417 ();
 FILLCELL_X32 FILLER_236_449 ();
 FILLCELL_X32 FILLER_236_481 ();
 FILLCELL_X32 FILLER_236_513 ();
 FILLCELL_X32 FILLER_236_545 ();
 FILLCELL_X32 FILLER_236_577 ();
 FILLCELL_X16 FILLER_236_609 ();
 FILLCELL_X4 FILLER_236_625 ();
 FILLCELL_X2 FILLER_236_629 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X32 FILLER_236_1752 ();
 FILLCELL_X32 FILLER_236_1784 ();
 FILLCELL_X32 FILLER_236_1816 ();
 FILLCELL_X32 FILLER_236_1848 ();
 FILLCELL_X8 FILLER_236_1880 ();
 FILLCELL_X4 FILLER_236_1888 ();
 FILLCELL_X2 FILLER_236_1892 ();
 FILLCELL_X32 FILLER_236_1895 ();
 FILLCELL_X32 FILLER_236_1927 ();
 FILLCELL_X32 FILLER_236_1959 ();
 FILLCELL_X32 FILLER_236_1991 ();
 FILLCELL_X32 FILLER_236_2023 ();
 FILLCELL_X32 FILLER_236_2055 ();
 FILLCELL_X16 FILLER_236_2087 ();
 FILLCELL_X8 FILLER_236_2103 ();
 FILLCELL_X4 FILLER_236_2111 ();
 FILLCELL_X32 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_33 ();
 FILLCELL_X32 FILLER_237_65 ();
 FILLCELL_X32 FILLER_237_97 ();
 FILLCELL_X32 FILLER_237_129 ();
 FILLCELL_X32 FILLER_237_161 ();
 FILLCELL_X32 FILLER_237_193 ();
 FILLCELL_X32 FILLER_237_225 ();
 FILLCELL_X32 FILLER_237_257 ();
 FILLCELL_X32 FILLER_237_289 ();
 FILLCELL_X32 FILLER_237_321 ();
 FILLCELL_X32 FILLER_237_353 ();
 FILLCELL_X32 FILLER_237_385 ();
 FILLCELL_X32 FILLER_237_417 ();
 FILLCELL_X32 FILLER_237_449 ();
 FILLCELL_X32 FILLER_237_481 ();
 FILLCELL_X32 FILLER_237_513 ();
 FILLCELL_X32 FILLER_237_545 ();
 FILLCELL_X32 FILLER_237_577 ();
 FILLCELL_X32 FILLER_237_609 ();
 FILLCELL_X32 FILLER_237_641 ();
 FILLCELL_X32 FILLER_237_673 ();
 FILLCELL_X32 FILLER_237_705 ();
 FILLCELL_X32 FILLER_237_737 ();
 FILLCELL_X32 FILLER_237_769 ();
 FILLCELL_X32 FILLER_237_801 ();
 FILLCELL_X32 FILLER_237_833 ();
 FILLCELL_X32 FILLER_237_865 ();
 FILLCELL_X32 FILLER_237_897 ();
 FILLCELL_X32 FILLER_237_929 ();
 FILLCELL_X32 FILLER_237_961 ();
 FILLCELL_X32 FILLER_237_993 ();
 FILLCELL_X32 FILLER_237_1025 ();
 FILLCELL_X32 FILLER_237_1057 ();
 FILLCELL_X32 FILLER_237_1089 ();
 FILLCELL_X32 FILLER_237_1121 ();
 FILLCELL_X32 FILLER_237_1153 ();
 FILLCELL_X32 FILLER_237_1185 ();
 FILLCELL_X32 FILLER_237_1217 ();
 FILLCELL_X8 FILLER_237_1249 ();
 FILLCELL_X4 FILLER_237_1257 ();
 FILLCELL_X2 FILLER_237_1261 ();
 FILLCELL_X32 FILLER_237_1264 ();
 FILLCELL_X32 FILLER_237_1296 ();
 FILLCELL_X32 FILLER_237_1328 ();
 FILLCELL_X32 FILLER_237_1360 ();
 FILLCELL_X32 FILLER_237_1392 ();
 FILLCELL_X32 FILLER_237_1424 ();
 FILLCELL_X32 FILLER_237_1456 ();
 FILLCELL_X32 FILLER_237_1488 ();
 FILLCELL_X32 FILLER_237_1520 ();
 FILLCELL_X32 FILLER_237_1552 ();
 FILLCELL_X32 FILLER_237_1584 ();
 FILLCELL_X32 FILLER_237_1616 ();
 FILLCELL_X32 FILLER_237_1648 ();
 FILLCELL_X32 FILLER_237_1680 ();
 FILLCELL_X32 FILLER_237_1712 ();
 FILLCELL_X32 FILLER_237_1744 ();
 FILLCELL_X32 FILLER_237_1776 ();
 FILLCELL_X32 FILLER_237_1808 ();
 FILLCELL_X32 FILLER_237_1840 ();
 FILLCELL_X32 FILLER_237_1872 ();
 FILLCELL_X32 FILLER_237_1904 ();
 FILLCELL_X32 FILLER_237_1936 ();
 FILLCELL_X32 FILLER_237_1968 ();
 FILLCELL_X32 FILLER_237_2000 ();
 FILLCELL_X32 FILLER_237_2032 ();
 FILLCELL_X32 FILLER_237_2064 ();
 FILLCELL_X16 FILLER_237_2096 ();
 FILLCELL_X2 FILLER_237_2112 ();
 FILLCELL_X1 FILLER_237_2114 ();
 FILLCELL_X32 FILLER_238_1 ();
 FILLCELL_X32 FILLER_238_33 ();
 FILLCELL_X32 FILLER_238_65 ();
 FILLCELL_X32 FILLER_238_97 ();
 FILLCELL_X32 FILLER_238_129 ();
 FILLCELL_X32 FILLER_238_161 ();
 FILLCELL_X32 FILLER_238_193 ();
 FILLCELL_X32 FILLER_238_225 ();
 FILLCELL_X32 FILLER_238_257 ();
 FILLCELL_X32 FILLER_238_289 ();
 FILLCELL_X32 FILLER_238_321 ();
 FILLCELL_X32 FILLER_238_353 ();
 FILLCELL_X32 FILLER_238_385 ();
 FILLCELL_X32 FILLER_238_417 ();
 FILLCELL_X32 FILLER_238_449 ();
 FILLCELL_X32 FILLER_238_481 ();
 FILLCELL_X32 FILLER_238_513 ();
 FILLCELL_X32 FILLER_238_545 ();
 FILLCELL_X32 FILLER_238_577 ();
 FILLCELL_X16 FILLER_238_609 ();
 FILLCELL_X4 FILLER_238_625 ();
 FILLCELL_X2 FILLER_238_629 ();
 FILLCELL_X32 FILLER_238_632 ();
 FILLCELL_X32 FILLER_238_664 ();
 FILLCELL_X32 FILLER_238_696 ();
 FILLCELL_X32 FILLER_238_728 ();
 FILLCELL_X32 FILLER_238_760 ();
 FILLCELL_X32 FILLER_238_792 ();
 FILLCELL_X32 FILLER_238_824 ();
 FILLCELL_X32 FILLER_238_856 ();
 FILLCELL_X32 FILLER_238_888 ();
 FILLCELL_X32 FILLER_238_920 ();
 FILLCELL_X32 FILLER_238_952 ();
 FILLCELL_X32 FILLER_238_984 ();
 FILLCELL_X32 FILLER_238_1016 ();
 FILLCELL_X32 FILLER_238_1048 ();
 FILLCELL_X32 FILLER_238_1080 ();
 FILLCELL_X32 FILLER_238_1112 ();
 FILLCELL_X32 FILLER_238_1144 ();
 FILLCELL_X32 FILLER_238_1176 ();
 FILLCELL_X32 FILLER_238_1208 ();
 FILLCELL_X32 FILLER_238_1240 ();
 FILLCELL_X32 FILLER_238_1272 ();
 FILLCELL_X32 FILLER_238_1304 ();
 FILLCELL_X32 FILLER_238_1336 ();
 FILLCELL_X32 FILLER_238_1368 ();
 FILLCELL_X32 FILLER_238_1400 ();
 FILLCELL_X32 FILLER_238_1432 ();
 FILLCELL_X32 FILLER_238_1464 ();
 FILLCELL_X32 FILLER_238_1496 ();
 FILLCELL_X32 FILLER_238_1528 ();
 FILLCELL_X32 FILLER_238_1560 ();
 FILLCELL_X32 FILLER_238_1592 ();
 FILLCELL_X32 FILLER_238_1624 ();
 FILLCELL_X32 FILLER_238_1656 ();
 FILLCELL_X32 FILLER_238_1688 ();
 FILLCELL_X32 FILLER_238_1720 ();
 FILLCELL_X32 FILLER_238_1752 ();
 FILLCELL_X32 FILLER_238_1784 ();
 FILLCELL_X32 FILLER_238_1816 ();
 FILLCELL_X32 FILLER_238_1848 ();
 FILLCELL_X8 FILLER_238_1880 ();
 FILLCELL_X4 FILLER_238_1888 ();
 FILLCELL_X2 FILLER_238_1892 ();
 FILLCELL_X32 FILLER_238_1895 ();
 FILLCELL_X32 FILLER_238_1927 ();
 FILLCELL_X32 FILLER_238_1959 ();
 FILLCELL_X32 FILLER_238_1991 ();
 FILLCELL_X32 FILLER_238_2023 ();
 FILLCELL_X32 FILLER_238_2055 ();
 FILLCELL_X16 FILLER_238_2087 ();
 FILLCELL_X8 FILLER_238_2103 ();
 FILLCELL_X4 FILLER_238_2111 ();
 FILLCELL_X32 FILLER_239_1 ();
 FILLCELL_X32 FILLER_239_33 ();
 FILLCELL_X32 FILLER_239_65 ();
 FILLCELL_X32 FILLER_239_97 ();
 FILLCELL_X32 FILLER_239_129 ();
 FILLCELL_X32 FILLER_239_161 ();
 FILLCELL_X32 FILLER_239_193 ();
 FILLCELL_X32 FILLER_239_225 ();
 FILLCELL_X32 FILLER_239_257 ();
 FILLCELL_X32 FILLER_239_289 ();
 FILLCELL_X32 FILLER_239_321 ();
 FILLCELL_X32 FILLER_239_353 ();
 FILLCELL_X32 FILLER_239_385 ();
 FILLCELL_X32 FILLER_239_417 ();
 FILLCELL_X32 FILLER_239_449 ();
 FILLCELL_X32 FILLER_239_481 ();
 FILLCELL_X32 FILLER_239_513 ();
 FILLCELL_X32 FILLER_239_545 ();
 FILLCELL_X32 FILLER_239_577 ();
 FILLCELL_X32 FILLER_239_609 ();
 FILLCELL_X32 FILLER_239_641 ();
 FILLCELL_X32 FILLER_239_673 ();
 FILLCELL_X32 FILLER_239_705 ();
 FILLCELL_X32 FILLER_239_737 ();
 FILLCELL_X32 FILLER_239_769 ();
 FILLCELL_X32 FILLER_239_801 ();
 FILLCELL_X32 FILLER_239_833 ();
 FILLCELL_X32 FILLER_239_865 ();
 FILLCELL_X32 FILLER_239_897 ();
 FILLCELL_X32 FILLER_239_929 ();
 FILLCELL_X32 FILLER_239_961 ();
 FILLCELL_X32 FILLER_239_993 ();
 FILLCELL_X32 FILLER_239_1025 ();
 FILLCELL_X32 FILLER_239_1057 ();
 FILLCELL_X32 FILLER_239_1089 ();
 FILLCELL_X32 FILLER_239_1121 ();
 FILLCELL_X32 FILLER_239_1153 ();
 FILLCELL_X32 FILLER_239_1185 ();
 FILLCELL_X32 FILLER_239_1217 ();
 FILLCELL_X8 FILLER_239_1249 ();
 FILLCELL_X4 FILLER_239_1257 ();
 FILLCELL_X2 FILLER_239_1261 ();
 FILLCELL_X32 FILLER_239_1264 ();
 FILLCELL_X32 FILLER_239_1296 ();
 FILLCELL_X32 FILLER_239_1328 ();
 FILLCELL_X32 FILLER_239_1360 ();
 FILLCELL_X32 FILLER_239_1392 ();
 FILLCELL_X32 FILLER_239_1424 ();
 FILLCELL_X32 FILLER_239_1456 ();
 FILLCELL_X32 FILLER_239_1488 ();
 FILLCELL_X32 FILLER_239_1520 ();
 FILLCELL_X32 FILLER_239_1552 ();
 FILLCELL_X32 FILLER_239_1584 ();
 FILLCELL_X32 FILLER_239_1616 ();
 FILLCELL_X32 FILLER_239_1648 ();
 FILLCELL_X32 FILLER_239_1680 ();
 FILLCELL_X32 FILLER_239_1712 ();
 FILLCELL_X32 FILLER_239_1744 ();
 FILLCELL_X32 FILLER_239_1776 ();
 FILLCELL_X32 FILLER_239_1808 ();
 FILLCELL_X32 FILLER_239_1840 ();
 FILLCELL_X32 FILLER_239_1872 ();
 FILLCELL_X32 FILLER_239_1904 ();
 FILLCELL_X32 FILLER_239_1936 ();
 FILLCELL_X32 FILLER_239_1968 ();
 FILLCELL_X32 FILLER_239_2000 ();
 FILLCELL_X32 FILLER_239_2032 ();
 FILLCELL_X32 FILLER_239_2064 ();
 FILLCELL_X16 FILLER_239_2096 ();
 FILLCELL_X2 FILLER_239_2112 ();
 FILLCELL_X1 FILLER_239_2114 ();
 FILLCELL_X32 FILLER_240_1 ();
 FILLCELL_X32 FILLER_240_33 ();
 FILLCELL_X32 FILLER_240_65 ();
 FILLCELL_X32 FILLER_240_97 ();
 FILLCELL_X32 FILLER_240_129 ();
 FILLCELL_X32 FILLER_240_161 ();
 FILLCELL_X32 FILLER_240_193 ();
 FILLCELL_X32 FILLER_240_225 ();
 FILLCELL_X32 FILLER_240_257 ();
 FILLCELL_X32 FILLER_240_289 ();
 FILLCELL_X32 FILLER_240_321 ();
 FILLCELL_X32 FILLER_240_353 ();
 FILLCELL_X32 FILLER_240_385 ();
 FILLCELL_X32 FILLER_240_417 ();
 FILLCELL_X32 FILLER_240_449 ();
 FILLCELL_X32 FILLER_240_481 ();
 FILLCELL_X32 FILLER_240_513 ();
 FILLCELL_X32 FILLER_240_545 ();
 FILLCELL_X32 FILLER_240_577 ();
 FILLCELL_X16 FILLER_240_609 ();
 FILLCELL_X4 FILLER_240_625 ();
 FILLCELL_X2 FILLER_240_629 ();
 FILLCELL_X32 FILLER_240_632 ();
 FILLCELL_X32 FILLER_240_664 ();
 FILLCELL_X32 FILLER_240_696 ();
 FILLCELL_X32 FILLER_240_728 ();
 FILLCELL_X32 FILLER_240_760 ();
 FILLCELL_X32 FILLER_240_792 ();
 FILLCELL_X32 FILLER_240_824 ();
 FILLCELL_X32 FILLER_240_856 ();
 FILLCELL_X32 FILLER_240_888 ();
 FILLCELL_X32 FILLER_240_920 ();
 FILLCELL_X32 FILLER_240_952 ();
 FILLCELL_X32 FILLER_240_984 ();
 FILLCELL_X32 FILLER_240_1016 ();
 FILLCELL_X32 FILLER_240_1048 ();
 FILLCELL_X32 FILLER_240_1080 ();
 FILLCELL_X32 FILLER_240_1112 ();
 FILLCELL_X32 FILLER_240_1144 ();
 FILLCELL_X32 FILLER_240_1176 ();
 FILLCELL_X32 FILLER_240_1208 ();
 FILLCELL_X32 FILLER_240_1240 ();
 FILLCELL_X32 FILLER_240_1272 ();
 FILLCELL_X32 FILLER_240_1304 ();
 FILLCELL_X32 FILLER_240_1336 ();
 FILLCELL_X32 FILLER_240_1368 ();
 FILLCELL_X32 FILLER_240_1400 ();
 FILLCELL_X32 FILLER_240_1432 ();
 FILLCELL_X32 FILLER_240_1464 ();
 FILLCELL_X32 FILLER_240_1496 ();
 FILLCELL_X32 FILLER_240_1528 ();
 FILLCELL_X32 FILLER_240_1560 ();
 FILLCELL_X32 FILLER_240_1592 ();
 FILLCELL_X32 FILLER_240_1624 ();
 FILLCELL_X32 FILLER_240_1656 ();
 FILLCELL_X32 FILLER_240_1688 ();
 FILLCELL_X32 FILLER_240_1720 ();
 FILLCELL_X32 FILLER_240_1752 ();
 FILLCELL_X32 FILLER_240_1784 ();
 FILLCELL_X32 FILLER_240_1816 ();
 FILLCELL_X32 FILLER_240_1848 ();
 FILLCELL_X8 FILLER_240_1880 ();
 FILLCELL_X4 FILLER_240_1888 ();
 FILLCELL_X2 FILLER_240_1892 ();
 FILLCELL_X32 FILLER_240_1895 ();
 FILLCELL_X32 FILLER_240_1927 ();
 FILLCELL_X32 FILLER_240_1959 ();
 FILLCELL_X32 FILLER_240_1991 ();
 FILLCELL_X32 FILLER_240_2023 ();
 FILLCELL_X32 FILLER_240_2055 ();
 FILLCELL_X16 FILLER_240_2087 ();
 FILLCELL_X8 FILLER_240_2103 ();
 FILLCELL_X4 FILLER_240_2111 ();
 FILLCELL_X32 FILLER_241_1 ();
 FILLCELL_X32 FILLER_241_33 ();
 FILLCELL_X32 FILLER_241_65 ();
 FILLCELL_X32 FILLER_241_97 ();
 FILLCELL_X32 FILLER_241_129 ();
 FILLCELL_X32 FILLER_241_161 ();
 FILLCELL_X32 FILLER_241_193 ();
 FILLCELL_X32 FILLER_241_225 ();
 FILLCELL_X32 FILLER_241_257 ();
 FILLCELL_X32 FILLER_241_289 ();
 FILLCELL_X32 FILLER_241_321 ();
 FILLCELL_X32 FILLER_241_353 ();
 FILLCELL_X32 FILLER_241_385 ();
 FILLCELL_X32 FILLER_241_417 ();
 FILLCELL_X32 FILLER_241_449 ();
 FILLCELL_X32 FILLER_241_481 ();
 FILLCELL_X32 FILLER_241_513 ();
 FILLCELL_X32 FILLER_241_545 ();
 FILLCELL_X32 FILLER_241_577 ();
 FILLCELL_X32 FILLER_241_609 ();
 FILLCELL_X32 FILLER_241_641 ();
 FILLCELL_X32 FILLER_241_673 ();
 FILLCELL_X32 FILLER_241_705 ();
 FILLCELL_X32 FILLER_241_737 ();
 FILLCELL_X32 FILLER_241_769 ();
 FILLCELL_X32 FILLER_241_801 ();
 FILLCELL_X32 FILLER_241_833 ();
 FILLCELL_X32 FILLER_241_865 ();
 FILLCELL_X32 FILLER_241_897 ();
 FILLCELL_X32 FILLER_241_929 ();
 FILLCELL_X32 FILLER_241_961 ();
 FILLCELL_X32 FILLER_241_993 ();
 FILLCELL_X32 FILLER_241_1025 ();
 FILLCELL_X32 FILLER_241_1057 ();
 FILLCELL_X32 FILLER_241_1089 ();
 FILLCELL_X32 FILLER_241_1121 ();
 FILLCELL_X32 FILLER_241_1153 ();
 FILLCELL_X32 FILLER_241_1185 ();
 FILLCELL_X32 FILLER_241_1217 ();
 FILLCELL_X8 FILLER_241_1249 ();
 FILLCELL_X4 FILLER_241_1257 ();
 FILLCELL_X2 FILLER_241_1261 ();
 FILLCELL_X32 FILLER_241_1264 ();
 FILLCELL_X32 FILLER_241_1296 ();
 FILLCELL_X32 FILLER_241_1328 ();
 FILLCELL_X32 FILLER_241_1360 ();
 FILLCELL_X32 FILLER_241_1392 ();
 FILLCELL_X32 FILLER_241_1424 ();
 FILLCELL_X32 FILLER_241_1456 ();
 FILLCELL_X32 FILLER_241_1488 ();
 FILLCELL_X32 FILLER_241_1520 ();
 FILLCELL_X32 FILLER_241_1552 ();
 FILLCELL_X32 FILLER_241_1584 ();
 FILLCELL_X32 FILLER_241_1616 ();
 FILLCELL_X32 FILLER_241_1648 ();
 FILLCELL_X32 FILLER_241_1680 ();
 FILLCELL_X32 FILLER_241_1712 ();
 FILLCELL_X32 FILLER_241_1744 ();
 FILLCELL_X32 FILLER_241_1776 ();
 FILLCELL_X32 FILLER_241_1808 ();
 FILLCELL_X32 FILLER_241_1840 ();
 FILLCELL_X32 FILLER_241_1872 ();
 FILLCELL_X32 FILLER_241_1904 ();
 FILLCELL_X32 FILLER_241_1936 ();
 FILLCELL_X32 FILLER_241_1968 ();
 FILLCELL_X32 FILLER_241_2000 ();
 FILLCELL_X32 FILLER_241_2032 ();
 FILLCELL_X32 FILLER_241_2064 ();
 FILLCELL_X16 FILLER_241_2096 ();
 FILLCELL_X2 FILLER_241_2112 ();
 FILLCELL_X1 FILLER_241_2114 ();
 FILLCELL_X32 FILLER_242_1 ();
 FILLCELL_X32 FILLER_242_33 ();
 FILLCELL_X32 FILLER_242_65 ();
 FILLCELL_X32 FILLER_242_97 ();
 FILLCELL_X32 FILLER_242_129 ();
 FILLCELL_X32 FILLER_242_161 ();
 FILLCELL_X32 FILLER_242_193 ();
 FILLCELL_X32 FILLER_242_225 ();
 FILLCELL_X32 FILLER_242_257 ();
 FILLCELL_X32 FILLER_242_289 ();
 FILLCELL_X32 FILLER_242_321 ();
 FILLCELL_X32 FILLER_242_353 ();
 FILLCELL_X32 FILLER_242_385 ();
 FILLCELL_X32 FILLER_242_417 ();
 FILLCELL_X32 FILLER_242_449 ();
 FILLCELL_X32 FILLER_242_481 ();
 FILLCELL_X32 FILLER_242_513 ();
 FILLCELL_X32 FILLER_242_545 ();
 FILLCELL_X32 FILLER_242_577 ();
 FILLCELL_X16 FILLER_242_609 ();
 FILLCELL_X4 FILLER_242_625 ();
 FILLCELL_X2 FILLER_242_629 ();
 FILLCELL_X32 FILLER_242_632 ();
 FILLCELL_X32 FILLER_242_664 ();
 FILLCELL_X32 FILLER_242_696 ();
 FILLCELL_X32 FILLER_242_728 ();
 FILLCELL_X32 FILLER_242_760 ();
 FILLCELL_X32 FILLER_242_792 ();
 FILLCELL_X32 FILLER_242_824 ();
 FILLCELL_X32 FILLER_242_856 ();
 FILLCELL_X32 FILLER_242_888 ();
 FILLCELL_X32 FILLER_242_920 ();
 FILLCELL_X32 FILLER_242_952 ();
 FILLCELL_X32 FILLER_242_984 ();
 FILLCELL_X32 FILLER_242_1016 ();
 FILLCELL_X32 FILLER_242_1048 ();
 FILLCELL_X32 FILLER_242_1080 ();
 FILLCELL_X32 FILLER_242_1112 ();
 FILLCELL_X32 FILLER_242_1144 ();
 FILLCELL_X32 FILLER_242_1176 ();
 FILLCELL_X32 FILLER_242_1208 ();
 FILLCELL_X32 FILLER_242_1240 ();
 FILLCELL_X32 FILLER_242_1272 ();
 FILLCELL_X32 FILLER_242_1304 ();
 FILLCELL_X32 FILLER_242_1336 ();
 FILLCELL_X32 FILLER_242_1368 ();
 FILLCELL_X32 FILLER_242_1400 ();
 FILLCELL_X32 FILLER_242_1432 ();
 FILLCELL_X32 FILLER_242_1464 ();
 FILLCELL_X32 FILLER_242_1496 ();
 FILLCELL_X32 FILLER_242_1528 ();
 FILLCELL_X32 FILLER_242_1560 ();
 FILLCELL_X32 FILLER_242_1592 ();
 FILLCELL_X32 FILLER_242_1624 ();
 FILLCELL_X32 FILLER_242_1656 ();
 FILLCELL_X32 FILLER_242_1688 ();
 FILLCELL_X32 FILLER_242_1720 ();
 FILLCELL_X32 FILLER_242_1752 ();
 FILLCELL_X32 FILLER_242_1784 ();
 FILLCELL_X32 FILLER_242_1816 ();
 FILLCELL_X32 FILLER_242_1848 ();
 FILLCELL_X8 FILLER_242_1880 ();
 FILLCELL_X4 FILLER_242_1888 ();
 FILLCELL_X2 FILLER_242_1892 ();
 FILLCELL_X32 FILLER_242_1895 ();
 FILLCELL_X32 FILLER_242_1927 ();
 FILLCELL_X32 FILLER_242_1959 ();
 FILLCELL_X32 FILLER_242_1991 ();
 FILLCELL_X32 FILLER_242_2023 ();
 FILLCELL_X32 FILLER_242_2055 ();
 FILLCELL_X16 FILLER_242_2087 ();
 FILLCELL_X8 FILLER_242_2103 ();
 FILLCELL_X4 FILLER_242_2111 ();
 FILLCELL_X32 FILLER_243_1 ();
 FILLCELL_X32 FILLER_243_33 ();
 FILLCELL_X32 FILLER_243_65 ();
 FILLCELL_X32 FILLER_243_97 ();
 FILLCELL_X32 FILLER_243_129 ();
 FILLCELL_X32 FILLER_243_161 ();
 FILLCELL_X32 FILLER_243_193 ();
 FILLCELL_X32 FILLER_243_225 ();
 FILLCELL_X32 FILLER_243_257 ();
 FILLCELL_X32 FILLER_243_289 ();
 FILLCELL_X32 FILLER_243_321 ();
 FILLCELL_X32 FILLER_243_353 ();
 FILLCELL_X32 FILLER_243_385 ();
 FILLCELL_X32 FILLER_243_417 ();
 FILLCELL_X32 FILLER_243_449 ();
 FILLCELL_X32 FILLER_243_481 ();
 FILLCELL_X32 FILLER_243_513 ();
 FILLCELL_X32 FILLER_243_545 ();
 FILLCELL_X32 FILLER_243_577 ();
 FILLCELL_X32 FILLER_243_609 ();
 FILLCELL_X32 FILLER_243_641 ();
 FILLCELL_X32 FILLER_243_673 ();
 FILLCELL_X32 FILLER_243_705 ();
 FILLCELL_X32 FILLER_243_737 ();
 FILLCELL_X32 FILLER_243_769 ();
 FILLCELL_X32 FILLER_243_801 ();
 FILLCELL_X32 FILLER_243_833 ();
 FILLCELL_X32 FILLER_243_865 ();
 FILLCELL_X32 FILLER_243_897 ();
 FILLCELL_X32 FILLER_243_929 ();
 FILLCELL_X32 FILLER_243_961 ();
 FILLCELL_X32 FILLER_243_993 ();
 FILLCELL_X32 FILLER_243_1025 ();
 FILLCELL_X32 FILLER_243_1057 ();
 FILLCELL_X32 FILLER_243_1089 ();
 FILLCELL_X32 FILLER_243_1121 ();
 FILLCELL_X32 FILLER_243_1153 ();
 FILLCELL_X32 FILLER_243_1185 ();
 FILLCELL_X32 FILLER_243_1217 ();
 FILLCELL_X8 FILLER_243_1249 ();
 FILLCELL_X4 FILLER_243_1257 ();
 FILLCELL_X2 FILLER_243_1261 ();
 FILLCELL_X32 FILLER_243_1264 ();
 FILLCELL_X32 FILLER_243_1296 ();
 FILLCELL_X32 FILLER_243_1328 ();
 FILLCELL_X32 FILLER_243_1360 ();
 FILLCELL_X32 FILLER_243_1392 ();
 FILLCELL_X32 FILLER_243_1424 ();
 FILLCELL_X32 FILLER_243_1456 ();
 FILLCELL_X32 FILLER_243_1488 ();
 FILLCELL_X32 FILLER_243_1520 ();
 FILLCELL_X32 FILLER_243_1552 ();
 FILLCELL_X32 FILLER_243_1584 ();
 FILLCELL_X32 FILLER_243_1616 ();
 FILLCELL_X32 FILLER_243_1648 ();
 FILLCELL_X32 FILLER_243_1680 ();
 FILLCELL_X32 FILLER_243_1712 ();
 FILLCELL_X32 FILLER_243_1744 ();
 FILLCELL_X32 FILLER_243_1776 ();
 FILLCELL_X32 FILLER_243_1808 ();
 FILLCELL_X32 FILLER_243_1840 ();
 FILLCELL_X32 FILLER_243_1872 ();
 FILLCELL_X32 FILLER_243_1904 ();
 FILLCELL_X32 FILLER_243_1936 ();
 FILLCELL_X32 FILLER_243_1968 ();
 FILLCELL_X32 FILLER_243_2000 ();
 FILLCELL_X32 FILLER_243_2032 ();
 FILLCELL_X32 FILLER_243_2064 ();
 FILLCELL_X16 FILLER_243_2096 ();
 FILLCELL_X2 FILLER_243_2112 ();
 FILLCELL_X1 FILLER_243_2114 ();
 FILLCELL_X32 FILLER_244_1 ();
 FILLCELL_X32 FILLER_244_33 ();
 FILLCELL_X32 FILLER_244_65 ();
 FILLCELL_X32 FILLER_244_97 ();
 FILLCELL_X32 FILLER_244_129 ();
 FILLCELL_X32 FILLER_244_161 ();
 FILLCELL_X32 FILLER_244_193 ();
 FILLCELL_X32 FILLER_244_225 ();
 FILLCELL_X32 FILLER_244_257 ();
 FILLCELL_X32 FILLER_244_289 ();
 FILLCELL_X32 FILLER_244_321 ();
 FILLCELL_X32 FILLER_244_353 ();
 FILLCELL_X32 FILLER_244_385 ();
 FILLCELL_X32 FILLER_244_417 ();
 FILLCELL_X32 FILLER_244_449 ();
 FILLCELL_X32 FILLER_244_481 ();
 FILLCELL_X32 FILLER_244_513 ();
 FILLCELL_X32 FILLER_244_545 ();
 FILLCELL_X32 FILLER_244_577 ();
 FILLCELL_X16 FILLER_244_609 ();
 FILLCELL_X4 FILLER_244_625 ();
 FILLCELL_X2 FILLER_244_629 ();
 FILLCELL_X32 FILLER_244_632 ();
 FILLCELL_X32 FILLER_244_664 ();
 FILLCELL_X32 FILLER_244_696 ();
 FILLCELL_X32 FILLER_244_728 ();
 FILLCELL_X32 FILLER_244_760 ();
 FILLCELL_X32 FILLER_244_792 ();
 FILLCELL_X32 FILLER_244_824 ();
 FILLCELL_X32 FILLER_244_856 ();
 FILLCELL_X32 FILLER_244_888 ();
 FILLCELL_X32 FILLER_244_920 ();
 FILLCELL_X32 FILLER_244_952 ();
 FILLCELL_X32 FILLER_244_984 ();
 FILLCELL_X32 FILLER_244_1016 ();
 FILLCELL_X32 FILLER_244_1048 ();
 FILLCELL_X32 FILLER_244_1080 ();
 FILLCELL_X32 FILLER_244_1112 ();
 FILLCELL_X32 FILLER_244_1144 ();
 FILLCELL_X32 FILLER_244_1176 ();
 FILLCELL_X32 FILLER_244_1208 ();
 FILLCELL_X32 FILLER_244_1240 ();
 FILLCELL_X32 FILLER_244_1272 ();
 FILLCELL_X32 FILLER_244_1304 ();
 FILLCELL_X32 FILLER_244_1336 ();
 FILLCELL_X32 FILLER_244_1368 ();
 FILLCELL_X32 FILLER_244_1400 ();
 FILLCELL_X32 FILLER_244_1432 ();
 FILLCELL_X32 FILLER_244_1464 ();
 FILLCELL_X32 FILLER_244_1496 ();
 FILLCELL_X32 FILLER_244_1528 ();
 FILLCELL_X32 FILLER_244_1560 ();
 FILLCELL_X32 FILLER_244_1592 ();
 FILLCELL_X32 FILLER_244_1624 ();
 FILLCELL_X32 FILLER_244_1656 ();
 FILLCELL_X32 FILLER_244_1688 ();
 FILLCELL_X32 FILLER_244_1720 ();
 FILLCELL_X32 FILLER_244_1752 ();
 FILLCELL_X32 FILLER_244_1784 ();
 FILLCELL_X32 FILLER_244_1816 ();
 FILLCELL_X32 FILLER_244_1848 ();
 FILLCELL_X8 FILLER_244_1880 ();
 FILLCELL_X4 FILLER_244_1888 ();
 FILLCELL_X2 FILLER_244_1892 ();
 FILLCELL_X32 FILLER_244_1895 ();
 FILLCELL_X32 FILLER_244_1927 ();
 FILLCELL_X32 FILLER_244_1959 ();
 FILLCELL_X32 FILLER_244_1991 ();
 FILLCELL_X32 FILLER_244_2023 ();
 FILLCELL_X32 FILLER_244_2055 ();
 FILLCELL_X16 FILLER_244_2087 ();
 FILLCELL_X8 FILLER_244_2103 ();
 FILLCELL_X4 FILLER_244_2111 ();
 FILLCELL_X32 FILLER_245_1 ();
 FILLCELL_X32 FILLER_245_33 ();
 FILLCELL_X32 FILLER_245_65 ();
 FILLCELL_X32 FILLER_245_97 ();
 FILLCELL_X32 FILLER_245_129 ();
 FILLCELL_X32 FILLER_245_161 ();
 FILLCELL_X32 FILLER_245_193 ();
 FILLCELL_X32 FILLER_245_225 ();
 FILLCELL_X32 FILLER_245_257 ();
 FILLCELL_X32 FILLER_245_289 ();
 FILLCELL_X32 FILLER_245_321 ();
 FILLCELL_X32 FILLER_245_353 ();
 FILLCELL_X32 FILLER_245_385 ();
 FILLCELL_X32 FILLER_245_417 ();
 FILLCELL_X32 FILLER_245_449 ();
 FILLCELL_X32 FILLER_245_481 ();
 FILLCELL_X32 FILLER_245_513 ();
 FILLCELL_X32 FILLER_245_545 ();
 FILLCELL_X32 FILLER_245_577 ();
 FILLCELL_X32 FILLER_245_609 ();
 FILLCELL_X32 FILLER_245_641 ();
 FILLCELL_X32 FILLER_245_673 ();
 FILLCELL_X32 FILLER_245_705 ();
 FILLCELL_X32 FILLER_245_737 ();
 FILLCELL_X32 FILLER_245_769 ();
 FILLCELL_X32 FILLER_245_801 ();
 FILLCELL_X32 FILLER_245_833 ();
 FILLCELL_X32 FILLER_245_865 ();
 FILLCELL_X32 FILLER_245_897 ();
 FILLCELL_X32 FILLER_245_929 ();
 FILLCELL_X32 FILLER_245_961 ();
 FILLCELL_X32 FILLER_245_993 ();
 FILLCELL_X32 FILLER_245_1025 ();
 FILLCELL_X32 FILLER_245_1057 ();
 FILLCELL_X32 FILLER_245_1089 ();
 FILLCELL_X32 FILLER_245_1121 ();
 FILLCELL_X32 FILLER_245_1153 ();
 FILLCELL_X32 FILLER_245_1185 ();
 FILLCELL_X32 FILLER_245_1217 ();
 FILLCELL_X8 FILLER_245_1249 ();
 FILLCELL_X4 FILLER_245_1257 ();
 FILLCELL_X2 FILLER_245_1261 ();
 FILLCELL_X32 FILLER_245_1264 ();
 FILLCELL_X32 FILLER_245_1296 ();
 FILLCELL_X32 FILLER_245_1328 ();
 FILLCELL_X32 FILLER_245_1360 ();
 FILLCELL_X32 FILLER_245_1392 ();
 FILLCELL_X32 FILLER_245_1424 ();
 FILLCELL_X32 FILLER_245_1456 ();
 FILLCELL_X32 FILLER_245_1488 ();
 FILLCELL_X32 FILLER_245_1520 ();
 FILLCELL_X32 FILLER_245_1552 ();
 FILLCELL_X32 FILLER_245_1584 ();
 FILLCELL_X32 FILLER_245_1616 ();
 FILLCELL_X32 FILLER_245_1648 ();
 FILLCELL_X32 FILLER_245_1680 ();
 FILLCELL_X32 FILLER_245_1712 ();
 FILLCELL_X32 FILLER_245_1744 ();
 FILLCELL_X32 FILLER_245_1776 ();
 FILLCELL_X32 FILLER_245_1808 ();
 FILLCELL_X32 FILLER_245_1840 ();
 FILLCELL_X32 FILLER_245_1872 ();
 FILLCELL_X32 FILLER_245_1904 ();
 FILLCELL_X32 FILLER_245_1936 ();
 FILLCELL_X32 FILLER_245_1968 ();
 FILLCELL_X32 FILLER_245_2000 ();
 FILLCELL_X32 FILLER_245_2032 ();
 FILLCELL_X32 FILLER_245_2064 ();
 FILLCELL_X16 FILLER_245_2096 ();
 FILLCELL_X2 FILLER_245_2112 ();
 FILLCELL_X1 FILLER_245_2114 ();
 FILLCELL_X32 FILLER_246_1 ();
 FILLCELL_X32 FILLER_246_33 ();
 FILLCELL_X32 FILLER_246_65 ();
 FILLCELL_X32 FILLER_246_97 ();
 FILLCELL_X32 FILLER_246_129 ();
 FILLCELL_X32 FILLER_246_161 ();
 FILLCELL_X32 FILLER_246_193 ();
 FILLCELL_X32 FILLER_246_225 ();
 FILLCELL_X32 FILLER_246_257 ();
 FILLCELL_X32 FILLER_246_289 ();
 FILLCELL_X32 FILLER_246_321 ();
 FILLCELL_X32 FILLER_246_353 ();
 FILLCELL_X32 FILLER_246_385 ();
 FILLCELL_X32 FILLER_246_417 ();
 FILLCELL_X32 FILLER_246_449 ();
 FILLCELL_X32 FILLER_246_481 ();
 FILLCELL_X32 FILLER_246_513 ();
 FILLCELL_X32 FILLER_246_545 ();
 FILLCELL_X32 FILLER_246_577 ();
 FILLCELL_X16 FILLER_246_609 ();
 FILLCELL_X4 FILLER_246_625 ();
 FILLCELL_X2 FILLER_246_629 ();
 FILLCELL_X32 FILLER_246_632 ();
 FILLCELL_X32 FILLER_246_664 ();
 FILLCELL_X32 FILLER_246_696 ();
 FILLCELL_X32 FILLER_246_728 ();
 FILLCELL_X32 FILLER_246_760 ();
 FILLCELL_X32 FILLER_246_792 ();
 FILLCELL_X32 FILLER_246_824 ();
 FILLCELL_X32 FILLER_246_856 ();
 FILLCELL_X32 FILLER_246_888 ();
 FILLCELL_X32 FILLER_246_920 ();
 FILLCELL_X32 FILLER_246_952 ();
 FILLCELL_X32 FILLER_246_984 ();
 FILLCELL_X32 FILLER_246_1016 ();
 FILLCELL_X32 FILLER_246_1048 ();
 FILLCELL_X32 FILLER_246_1080 ();
 FILLCELL_X32 FILLER_246_1112 ();
 FILLCELL_X32 FILLER_246_1144 ();
 FILLCELL_X32 FILLER_246_1176 ();
 FILLCELL_X32 FILLER_246_1208 ();
 FILLCELL_X32 FILLER_246_1240 ();
 FILLCELL_X32 FILLER_246_1272 ();
 FILLCELL_X32 FILLER_246_1304 ();
 FILLCELL_X32 FILLER_246_1336 ();
 FILLCELL_X32 FILLER_246_1368 ();
 FILLCELL_X32 FILLER_246_1400 ();
 FILLCELL_X32 FILLER_246_1432 ();
 FILLCELL_X32 FILLER_246_1464 ();
 FILLCELL_X32 FILLER_246_1496 ();
 FILLCELL_X32 FILLER_246_1528 ();
 FILLCELL_X32 FILLER_246_1560 ();
 FILLCELL_X32 FILLER_246_1592 ();
 FILLCELL_X32 FILLER_246_1624 ();
 FILLCELL_X32 FILLER_246_1656 ();
 FILLCELL_X32 FILLER_246_1688 ();
 FILLCELL_X32 FILLER_246_1720 ();
 FILLCELL_X32 FILLER_246_1752 ();
 FILLCELL_X32 FILLER_246_1784 ();
 FILLCELL_X32 FILLER_246_1816 ();
 FILLCELL_X32 FILLER_246_1848 ();
 FILLCELL_X8 FILLER_246_1880 ();
 FILLCELL_X4 FILLER_246_1888 ();
 FILLCELL_X2 FILLER_246_1892 ();
 FILLCELL_X32 FILLER_246_1895 ();
 FILLCELL_X32 FILLER_246_1927 ();
 FILLCELL_X32 FILLER_246_1959 ();
 FILLCELL_X32 FILLER_246_1991 ();
 FILLCELL_X32 FILLER_246_2023 ();
 FILLCELL_X32 FILLER_246_2055 ();
 FILLCELL_X16 FILLER_246_2087 ();
 FILLCELL_X8 FILLER_246_2103 ();
 FILLCELL_X4 FILLER_246_2111 ();
 FILLCELL_X32 FILLER_247_1 ();
 FILLCELL_X32 FILLER_247_33 ();
 FILLCELL_X32 FILLER_247_65 ();
 FILLCELL_X32 FILLER_247_97 ();
 FILLCELL_X32 FILLER_247_129 ();
 FILLCELL_X32 FILLER_247_161 ();
 FILLCELL_X32 FILLER_247_193 ();
 FILLCELL_X32 FILLER_247_225 ();
 FILLCELL_X32 FILLER_247_257 ();
 FILLCELL_X32 FILLER_247_289 ();
 FILLCELL_X32 FILLER_247_321 ();
 FILLCELL_X32 FILLER_247_353 ();
 FILLCELL_X32 FILLER_247_385 ();
 FILLCELL_X32 FILLER_247_417 ();
 FILLCELL_X32 FILLER_247_449 ();
 FILLCELL_X32 FILLER_247_481 ();
 FILLCELL_X32 FILLER_247_513 ();
 FILLCELL_X32 FILLER_247_545 ();
 FILLCELL_X32 FILLER_247_577 ();
 FILLCELL_X32 FILLER_247_609 ();
 FILLCELL_X32 FILLER_247_641 ();
 FILLCELL_X32 FILLER_247_673 ();
 FILLCELL_X32 FILLER_247_705 ();
 FILLCELL_X32 FILLER_247_737 ();
 FILLCELL_X32 FILLER_247_769 ();
 FILLCELL_X32 FILLER_247_801 ();
 FILLCELL_X32 FILLER_247_833 ();
 FILLCELL_X32 FILLER_247_865 ();
 FILLCELL_X32 FILLER_247_897 ();
 FILLCELL_X32 FILLER_247_929 ();
 FILLCELL_X32 FILLER_247_961 ();
 FILLCELL_X32 FILLER_247_993 ();
 FILLCELL_X32 FILLER_247_1025 ();
 FILLCELL_X32 FILLER_247_1057 ();
 FILLCELL_X32 FILLER_247_1089 ();
 FILLCELL_X32 FILLER_247_1121 ();
 FILLCELL_X32 FILLER_247_1153 ();
 FILLCELL_X32 FILLER_247_1185 ();
 FILLCELL_X32 FILLER_247_1217 ();
 FILLCELL_X8 FILLER_247_1249 ();
 FILLCELL_X4 FILLER_247_1257 ();
 FILLCELL_X2 FILLER_247_1261 ();
 FILLCELL_X32 FILLER_247_1264 ();
 FILLCELL_X32 FILLER_247_1296 ();
 FILLCELL_X32 FILLER_247_1328 ();
 FILLCELL_X32 FILLER_247_1360 ();
 FILLCELL_X32 FILLER_247_1392 ();
 FILLCELL_X32 FILLER_247_1424 ();
 FILLCELL_X32 FILLER_247_1456 ();
 FILLCELL_X32 FILLER_247_1488 ();
 FILLCELL_X32 FILLER_247_1520 ();
 FILLCELL_X32 FILLER_247_1552 ();
 FILLCELL_X32 FILLER_247_1584 ();
 FILLCELL_X32 FILLER_247_1616 ();
 FILLCELL_X32 FILLER_247_1648 ();
 FILLCELL_X32 FILLER_247_1680 ();
 FILLCELL_X32 FILLER_247_1712 ();
 FILLCELL_X32 FILLER_247_1744 ();
 FILLCELL_X32 FILLER_247_1776 ();
 FILLCELL_X32 FILLER_247_1808 ();
 FILLCELL_X32 FILLER_247_1840 ();
 FILLCELL_X32 FILLER_247_1872 ();
 FILLCELL_X32 FILLER_247_1904 ();
 FILLCELL_X32 FILLER_247_1936 ();
 FILLCELL_X32 FILLER_247_1968 ();
 FILLCELL_X32 FILLER_247_2000 ();
 FILLCELL_X32 FILLER_247_2032 ();
 FILLCELL_X32 FILLER_247_2064 ();
 FILLCELL_X16 FILLER_247_2096 ();
 FILLCELL_X2 FILLER_247_2112 ();
 FILLCELL_X1 FILLER_247_2114 ();
 FILLCELL_X32 FILLER_248_1 ();
 FILLCELL_X32 FILLER_248_33 ();
 FILLCELL_X32 FILLER_248_65 ();
 FILLCELL_X32 FILLER_248_97 ();
 FILLCELL_X32 FILLER_248_129 ();
 FILLCELL_X32 FILLER_248_161 ();
 FILLCELL_X32 FILLER_248_193 ();
 FILLCELL_X32 FILLER_248_225 ();
 FILLCELL_X32 FILLER_248_257 ();
 FILLCELL_X32 FILLER_248_289 ();
 FILLCELL_X32 FILLER_248_321 ();
 FILLCELL_X32 FILLER_248_353 ();
 FILLCELL_X32 FILLER_248_385 ();
 FILLCELL_X32 FILLER_248_417 ();
 FILLCELL_X32 FILLER_248_449 ();
 FILLCELL_X32 FILLER_248_481 ();
 FILLCELL_X32 FILLER_248_513 ();
 FILLCELL_X32 FILLER_248_545 ();
 FILLCELL_X32 FILLER_248_577 ();
 FILLCELL_X16 FILLER_248_609 ();
 FILLCELL_X4 FILLER_248_625 ();
 FILLCELL_X2 FILLER_248_629 ();
 FILLCELL_X32 FILLER_248_632 ();
 FILLCELL_X32 FILLER_248_664 ();
 FILLCELL_X32 FILLER_248_696 ();
 FILLCELL_X32 FILLER_248_728 ();
 FILLCELL_X32 FILLER_248_760 ();
 FILLCELL_X32 FILLER_248_792 ();
 FILLCELL_X32 FILLER_248_824 ();
 FILLCELL_X32 FILLER_248_856 ();
 FILLCELL_X32 FILLER_248_888 ();
 FILLCELL_X32 FILLER_248_920 ();
 FILLCELL_X32 FILLER_248_952 ();
 FILLCELL_X32 FILLER_248_984 ();
 FILLCELL_X32 FILLER_248_1016 ();
 FILLCELL_X32 FILLER_248_1048 ();
 FILLCELL_X32 FILLER_248_1080 ();
 FILLCELL_X32 FILLER_248_1112 ();
 FILLCELL_X32 FILLER_248_1144 ();
 FILLCELL_X32 FILLER_248_1176 ();
 FILLCELL_X32 FILLER_248_1208 ();
 FILLCELL_X32 FILLER_248_1240 ();
 FILLCELL_X32 FILLER_248_1272 ();
 FILLCELL_X32 FILLER_248_1304 ();
 FILLCELL_X32 FILLER_248_1336 ();
 FILLCELL_X32 FILLER_248_1368 ();
 FILLCELL_X32 FILLER_248_1400 ();
 FILLCELL_X32 FILLER_248_1432 ();
 FILLCELL_X32 FILLER_248_1464 ();
 FILLCELL_X32 FILLER_248_1496 ();
 FILLCELL_X32 FILLER_248_1528 ();
 FILLCELL_X32 FILLER_248_1560 ();
 FILLCELL_X32 FILLER_248_1592 ();
 FILLCELL_X32 FILLER_248_1624 ();
 FILLCELL_X32 FILLER_248_1656 ();
 FILLCELL_X32 FILLER_248_1688 ();
 FILLCELL_X32 FILLER_248_1720 ();
 FILLCELL_X32 FILLER_248_1752 ();
 FILLCELL_X32 FILLER_248_1784 ();
 FILLCELL_X32 FILLER_248_1816 ();
 FILLCELL_X32 FILLER_248_1848 ();
 FILLCELL_X8 FILLER_248_1880 ();
 FILLCELL_X4 FILLER_248_1888 ();
 FILLCELL_X2 FILLER_248_1892 ();
 FILLCELL_X32 FILLER_248_1895 ();
 FILLCELL_X32 FILLER_248_1927 ();
 FILLCELL_X32 FILLER_248_1959 ();
 FILLCELL_X32 FILLER_248_1991 ();
 FILLCELL_X32 FILLER_248_2023 ();
 FILLCELL_X32 FILLER_248_2055 ();
 FILLCELL_X16 FILLER_248_2087 ();
 FILLCELL_X8 FILLER_248_2103 ();
 FILLCELL_X4 FILLER_248_2111 ();
 FILLCELL_X32 FILLER_249_1 ();
 FILLCELL_X32 FILLER_249_33 ();
 FILLCELL_X32 FILLER_249_65 ();
 FILLCELL_X32 FILLER_249_97 ();
 FILLCELL_X32 FILLER_249_129 ();
 FILLCELL_X32 FILLER_249_161 ();
 FILLCELL_X32 FILLER_249_193 ();
 FILLCELL_X32 FILLER_249_225 ();
 FILLCELL_X32 FILLER_249_257 ();
 FILLCELL_X32 FILLER_249_289 ();
 FILLCELL_X32 FILLER_249_321 ();
 FILLCELL_X32 FILLER_249_353 ();
 FILLCELL_X32 FILLER_249_385 ();
 FILLCELL_X32 FILLER_249_417 ();
 FILLCELL_X32 FILLER_249_449 ();
 FILLCELL_X32 FILLER_249_481 ();
 FILLCELL_X32 FILLER_249_513 ();
 FILLCELL_X32 FILLER_249_545 ();
 FILLCELL_X32 FILLER_249_577 ();
 FILLCELL_X32 FILLER_249_609 ();
 FILLCELL_X32 FILLER_249_641 ();
 FILLCELL_X32 FILLER_249_673 ();
 FILLCELL_X32 FILLER_249_705 ();
 FILLCELL_X32 FILLER_249_737 ();
 FILLCELL_X32 FILLER_249_769 ();
 FILLCELL_X32 FILLER_249_801 ();
 FILLCELL_X32 FILLER_249_833 ();
 FILLCELL_X32 FILLER_249_865 ();
 FILLCELL_X32 FILLER_249_897 ();
 FILLCELL_X32 FILLER_249_929 ();
 FILLCELL_X32 FILLER_249_961 ();
 FILLCELL_X32 FILLER_249_993 ();
 FILLCELL_X32 FILLER_249_1025 ();
 FILLCELL_X32 FILLER_249_1057 ();
 FILLCELL_X32 FILLER_249_1089 ();
 FILLCELL_X32 FILLER_249_1121 ();
 FILLCELL_X32 FILLER_249_1153 ();
 FILLCELL_X32 FILLER_249_1185 ();
 FILLCELL_X32 FILLER_249_1217 ();
 FILLCELL_X8 FILLER_249_1249 ();
 FILLCELL_X4 FILLER_249_1257 ();
 FILLCELL_X2 FILLER_249_1261 ();
 FILLCELL_X32 FILLER_249_1264 ();
 FILLCELL_X32 FILLER_249_1296 ();
 FILLCELL_X32 FILLER_249_1328 ();
 FILLCELL_X32 FILLER_249_1360 ();
 FILLCELL_X32 FILLER_249_1392 ();
 FILLCELL_X32 FILLER_249_1424 ();
 FILLCELL_X32 FILLER_249_1456 ();
 FILLCELL_X32 FILLER_249_1488 ();
 FILLCELL_X32 FILLER_249_1520 ();
 FILLCELL_X32 FILLER_249_1552 ();
 FILLCELL_X32 FILLER_249_1584 ();
 FILLCELL_X32 FILLER_249_1616 ();
 FILLCELL_X32 FILLER_249_1648 ();
 FILLCELL_X32 FILLER_249_1680 ();
 FILLCELL_X32 FILLER_249_1712 ();
 FILLCELL_X32 FILLER_249_1744 ();
 FILLCELL_X32 FILLER_249_1776 ();
 FILLCELL_X32 FILLER_249_1808 ();
 FILLCELL_X32 FILLER_249_1840 ();
 FILLCELL_X32 FILLER_249_1872 ();
 FILLCELL_X32 FILLER_249_1904 ();
 FILLCELL_X32 FILLER_249_1936 ();
 FILLCELL_X32 FILLER_249_1968 ();
 FILLCELL_X32 FILLER_249_2000 ();
 FILLCELL_X32 FILLER_249_2032 ();
 FILLCELL_X32 FILLER_249_2064 ();
 FILLCELL_X16 FILLER_249_2096 ();
 FILLCELL_X2 FILLER_249_2112 ();
 FILLCELL_X1 FILLER_249_2114 ();
 FILLCELL_X32 FILLER_250_1 ();
 FILLCELL_X32 FILLER_250_33 ();
 FILLCELL_X32 FILLER_250_65 ();
 FILLCELL_X32 FILLER_250_97 ();
 FILLCELL_X32 FILLER_250_129 ();
 FILLCELL_X32 FILLER_250_161 ();
 FILLCELL_X32 FILLER_250_193 ();
 FILLCELL_X32 FILLER_250_225 ();
 FILLCELL_X32 FILLER_250_257 ();
 FILLCELL_X32 FILLER_250_289 ();
 FILLCELL_X32 FILLER_250_321 ();
 FILLCELL_X32 FILLER_250_353 ();
 FILLCELL_X32 FILLER_250_385 ();
 FILLCELL_X32 FILLER_250_417 ();
 FILLCELL_X32 FILLER_250_449 ();
 FILLCELL_X32 FILLER_250_481 ();
 FILLCELL_X32 FILLER_250_513 ();
 FILLCELL_X32 FILLER_250_545 ();
 FILLCELL_X32 FILLER_250_577 ();
 FILLCELL_X16 FILLER_250_609 ();
 FILLCELL_X4 FILLER_250_625 ();
 FILLCELL_X2 FILLER_250_629 ();
 FILLCELL_X32 FILLER_250_632 ();
 FILLCELL_X32 FILLER_250_664 ();
 FILLCELL_X32 FILLER_250_696 ();
 FILLCELL_X32 FILLER_250_728 ();
 FILLCELL_X32 FILLER_250_760 ();
 FILLCELL_X32 FILLER_250_792 ();
 FILLCELL_X32 FILLER_250_824 ();
 FILLCELL_X32 FILLER_250_856 ();
 FILLCELL_X32 FILLER_250_888 ();
 FILLCELL_X32 FILLER_250_920 ();
 FILLCELL_X32 FILLER_250_952 ();
 FILLCELL_X32 FILLER_250_984 ();
 FILLCELL_X32 FILLER_250_1016 ();
 FILLCELL_X32 FILLER_250_1048 ();
 FILLCELL_X32 FILLER_250_1080 ();
 FILLCELL_X32 FILLER_250_1112 ();
 FILLCELL_X32 FILLER_250_1144 ();
 FILLCELL_X32 FILLER_250_1176 ();
 FILLCELL_X32 FILLER_250_1208 ();
 FILLCELL_X32 FILLER_250_1240 ();
 FILLCELL_X32 FILLER_250_1272 ();
 FILLCELL_X32 FILLER_250_1304 ();
 FILLCELL_X32 FILLER_250_1336 ();
 FILLCELL_X32 FILLER_250_1368 ();
 FILLCELL_X32 FILLER_250_1400 ();
 FILLCELL_X32 FILLER_250_1432 ();
 FILLCELL_X32 FILLER_250_1464 ();
 FILLCELL_X32 FILLER_250_1496 ();
 FILLCELL_X32 FILLER_250_1528 ();
 FILLCELL_X32 FILLER_250_1560 ();
 FILLCELL_X32 FILLER_250_1592 ();
 FILLCELL_X32 FILLER_250_1624 ();
 FILLCELL_X32 FILLER_250_1656 ();
 FILLCELL_X32 FILLER_250_1688 ();
 FILLCELL_X32 FILLER_250_1720 ();
 FILLCELL_X32 FILLER_250_1752 ();
 FILLCELL_X32 FILLER_250_1784 ();
 FILLCELL_X32 FILLER_250_1816 ();
 FILLCELL_X32 FILLER_250_1848 ();
 FILLCELL_X8 FILLER_250_1880 ();
 FILLCELL_X4 FILLER_250_1888 ();
 FILLCELL_X2 FILLER_250_1892 ();
 FILLCELL_X32 FILLER_250_1895 ();
 FILLCELL_X32 FILLER_250_1927 ();
 FILLCELL_X32 FILLER_250_1959 ();
 FILLCELL_X32 FILLER_250_1991 ();
 FILLCELL_X32 FILLER_250_2023 ();
 FILLCELL_X32 FILLER_250_2055 ();
 FILLCELL_X16 FILLER_250_2087 ();
 FILLCELL_X8 FILLER_250_2103 ();
 FILLCELL_X4 FILLER_250_2111 ();
 FILLCELL_X32 FILLER_251_1 ();
 FILLCELL_X32 FILLER_251_33 ();
 FILLCELL_X32 FILLER_251_65 ();
 FILLCELL_X32 FILLER_251_97 ();
 FILLCELL_X32 FILLER_251_129 ();
 FILLCELL_X32 FILLER_251_161 ();
 FILLCELL_X32 FILLER_251_193 ();
 FILLCELL_X32 FILLER_251_225 ();
 FILLCELL_X32 FILLER_251_257 ();
 FILLCELL_X32 FILLER_251_289 ();
 FILLCELL_X32 FILLER_251_321 ();
 FILLCELL_X32 FILLER_251_353 ();
 FILLCELL_X32 FILLER_251_385 ();
 FILLCELL_X32 FILLER_251_417 ();
 FILLCELL_X32 FILLER_251_449 ();
 FILLCELL_X32 FILLER_251_481 ();
 FILLCELL_X32 FILLER_251_513 ();
 FILLCELL_X32 FILLER_251_545 ();
 FILLCELL_X32 FILLER_251_577 ();
 FILLCELL_X32 FILLER_251_609 ();
 FILLCELL_X32 FILLER_251_641 ();
 FILLCELL_X32 FILLER_251_673 ();
 FILLCELL_X32 FILLER_251_705 ();
 FILLCELL_X32 FILLER_251_737 ();
 FILLCELL_X32 FILLER_251_769 ();
 FILLCELL_X32 FILLER_251_801 ();
 FILLCELL_X32 FILLER_251_833 ();
 FILLCELL_X32 FILLER_251_865 ();
 FILLCELL_X32 FILLER_251_897 ();
 FILLCELL_X32 FILLER_251_929 ();
 FILLCELL_X32 FILLER_251_961 ();
 FILLCELL_X32 FILLER_251_993 ();
 FILLCELL_X32 FILLER_251_1025 ();
 FILLCELL_X32 FILLER_251_1057 ();
 FILLCELL_X32 FILLER_251_1089 ();
 FILLCELL_X32 FILLER_251_1121 ();
 FILLCELL_X32 FILLER_251_1153 ();
 FILLCELL_X32 FILLER_251_1185 ();
 FILLCELL_X32 FILLER_251_1217 ();
 FILLCELL_X8 FILLER_251_1249 ();
 FILLCELL_X4 FILLER_251_1257 ();
 FILLCELL_X2 FILLER_251_1261 ();
 FILLCELL_X32 FILLER_251_1264 ();
 FILLCELL_X32 FILLER_251_1296 ();
 FILLCELL_X32 FILLER_251_1328 ();
 FILLCELL_X32 FILLER_251_1360 ();
 FILLCELL_X32 FILLER_251_1392 ();
 FILLCELL_X32 FILLER_251_1424 ();
 FILLCELL_X32 FILLER_251_1456 ();
 FILLCELL_X32 FILLER_251_1488 ();
 FILLCELL_X32 FILLER_251_1520 ();
 FILLCELL_X32 FILLER_251_1552 ();
 FILLCELL_X32 FILLER_251_1584 ();
 FILLCELL_X32 FILLER_251_1616 ();
 FILLCELL_X32 FILLER_251_1648 ();
 FILLCELL_X32 FILLER_251_1680 ();
 FILLCELL_X32 FILLER_251_1712 ();
 FILLCELL_X32 FILLER_251_1744 ();
 FILLCELL_X32 FILLER_251_1776 ();
 FILLCELL_X32 FILLER_251_1808 ();
 FILLCELL_X32 FILLER_251_1840 ();
 FILLCELL_X32 FILLER_251_1872 ();
 FILLCELL_X32 FILLER_251_1904 ();
 FILLCELL_X32 FILLER_251_1936 ();
 FILLCELL_X32 FILLER_251_1968 ();
 FILLCELL_X32 FILLER_251_2000 ();
 FILLCELL_X32 FILLER_251_2032 ();
 FILLCELL_X32 FILLER_251_2064 ();
 FILLCELL_X16 FILLER_251_2096 ();
 FILLCELL_X2 FILLER_251_2112 ();
 FILLCELL_X1 FILLER_251_2114 ();
 FILLCELL_X32 FILLER_252_1 ();
 FILLCELL_X32 FILLER_252_33 ();
 FILLCELL_X32 FILLER_252_65 ();
 FILLCELL_X32 FILLER_252_97 ();
 FILLCELL_X32 FILLER_252_129 ();
 FILLCELL_X32 FILLER_252_161 ();
 FILLCELL_X32 FILLER_252_193 ();
 FILLCELL_X32 FILLER_252_225 ();
 FILLCELL_X32 FILLER_252_257 ();
 FILLCELL_X32 FILLER_252_289 ();
 FILLCELL_X32 FILLER_252_321 ();
 FILLCELL_X32 FILLER_252_353 ();
 FILLCELL_X32 FILLER_252_385 ();
 FILLCELL_X32 FILLER_252_417 ();
 FILLCELL_X32 FILLER_252_449 ();
 FILLCELL_X32 FILLER_252_481 ();
 FILLCELL_X32 FILLER_252_513 ();
 FILLCELL_X32 FILLER_252_545 ();
 FILLCELL_X32 FILLER_252_577 ();
 FILLCELL_X16 FILLER_252_609 ();
 FILLCELL_X4 FILLER_252_625 ();
 FILLCELL_X2 FILLER_252_629 ();
 FILLCELL_X32 FILLER_252_632 ();
 FILLCELL_X32 FILLER_252_664 ();
 FILLCELL_X32 FILLER_252_696 ();
 FILLCELL_X32 FILLER_252_728 ();
 FILLCELL_X32 FILLER_252_760 ();
 FILLCELL_X32 FILLER_252_792 ();
 FILLCELL_X32 FILLER_252_824 ();
 FILLCELL_X32 FILLER_252_856 ();
 FILLCELL_X32 FILLER_252_888 ();
 FILLCELL_X32 FILLER_252_920 ();
 FILLCELL_X32 FILLER_252_952 ();
 FILLCELL_X32 FILLER_252_984 ();
 FILLCELL_X32 FILLER_252_1016 ();
 FILLCELL_X32 FILLER_252_1048 ();
 FILLCELL_X32 FILLER_252_1080 ();
 FILLCELL_X32 FILLER_252_1112 ();
 FILLCELL_X32 FILLER_252_1144 ();
 FILLCELL_X32 FILLER_252_1176 ();
 FILLCELL_X32 FILLER_252_1208 ();
 FILLCELL_X32 FILLER_252_1240 ();
 FILLCELL_X32 FILLER_252_1272 ();
 FILLCELL_X32 FILLER_252_1304 ();
 FILLCELL_X32 FILLER_252_1336 ();
 FILLCELL_X32 FILLER_252_1368 ();
 FILLCELL_X32 FILLER_252_1400 ();
 FILLCELL_X32 FILLER_252_1432 ();
 FILLCELL_X32 FILLER_252_1464 ();
 FILLCELL_X32 FILLER_252_1496 ();
 FILLCELL_X32 FILLER_252_1528 ();
 FILLCELL_X32 FILLER_252_1560 ();
 FILLCELL_X32 FILLER_252_1592 ();
 FILLCELL_X32 FILLER_252_1624 ();
 FILLCELL_X32 FILLER_252_1656 ();
 FILLCELL_X32 FILLER_252_1688 ();
 FILLCELL_X32 FILLER_252_1720 ();
 FILLCELL_X32 FILLER_252_1752 ();
 FILLCELL_X32 FILLER_252_1784 ();
 FILLCELL_X32 FILLER_252_1816 ();
 FILLCELL_X32 FILLER_252_1848 ();
 FILLCELL_X8 FILLER_252_1880 ();
 FILLCELL_X4 FILLER_252_1888 ();
 FILLCELL_X2 FILLER_252_1892 ();
 FILLCELL_X32 FILLER_252_1895 ();
 FILLCELL_X32 FILLER_252_1927 ();
 FILLCELL_X32 FILLER_252_1959 ();
 FILLCELL_X32 FILLER_252_1991 ();
 FILLCELL_X32 FILLER_252_2023 ();
 FILLCELL_X32 FILLER_252_2055 ();
 FILLCELL_X16 FILLER_252_2087 ();
 FILLCELL_X8 FILLER_252_2103 ();
 FILLCELL_X4 FILLER_252_2111 ();
 FILLCELL_X32 FILLER_253_1 ();
 FILLCELL_X32 FILLER_253_33 ();
 FILLCELL_X32 FILLER_253_65 ();
 FILLCELL_X32 FILLER_253_97 ();
 FILLCELL_X32 FILLER_253_129 ();
 FILLCELL_X32 FILLER_253_161 ();
 FILLCELL_X32 FILLER_253_193 ();
 FILLCELL_X32 FILLER_253_225 ();
 FILLCELL_X32 FILLER_253_257 ();
 FILLCELL_X32 FILLER_253_289 ();
 FILLCELL_X32 FILLER_253_321 ();
 FILLCELL_X32 FILLER_253_353 ();
 FILLCELL_X32 FILLER_253_385 ();
 FILLCELL_X32 FILLER_253_417 ();
 FILLCELL_X32 FILLER_253_449 ();
 FILLCELL_X32 FILLER_253_481 ();
 FILLCELL_X32 FILLER_253_513 ();
 FILLCELL_X32 FILLER_253_545 ();
 FILLCELL_X32 FILLER_253_577 ();
 FILLCELL_X32 FILLER_253_609 ();
 FILLCELL_X32 FILLER_253_641 ();
 FILLCELL_X32 FILLER_253_673 ();
 FILLCELL_X32 FILLER_253_705 ();
 FILLCELL_X32 FILLER_253_737 ();
 FILLCELL_X32 FILLER_253_769 ();
 FILLCELL_X32 FILLER_253_801 ();
 FILLCELL_X32 FILLER_253_833 ();
 FILLCELL_X32 FILLER_253_865 ();
 FILLCELL_X32 FILLER_253_897 ();
 FILLCELL_X32 FILLER_253_929 ();
 FILLCELL_X32 FILLER_253_961 ();
 FILLCELL_X32 FILLER_253_993 ();
 FILLCELL_X32 FILLER_253_1025 ();
 FILLCELL_X32 FILLER_253_1057 ();
 FILLCELL_X32 FILLER_253_1089 ();
 FILLCELL_X32 FILLER_253_1121 ();
 FILLCELL_X32 FILLER_253_1153 ();
 FILLCELL_X32 FILLER_253_1185 ();
 FILLCELL_X32 FILLER_253_1217 ();
 FILLCELL_X8 FILLER_253_1249 ();
 FILLCELL_X4 FILLER_253_1257 ();
 FILLCELL_X2 FILLER_253_1261 ();
 FILLCELL_X32 FILLER_253_1264 ();
 FILLCELL_X32 FILLER_253_1296 ();
 FILLCELL_X32 FILLER_253_1328 ();
 FILLCELL_X32 FILLER_253_1360 ();
 FILLCELL_X32 FILLER_253_1392 ();
 FILLCELL_X32 FILLER_253_1424 ();
 FILLCELL_X32 FILLER_253_1456 ();
 FILLCELL_X32 FILLER_253_1488 ();
 FILLCELL_X32 FILLER_253_1520 ();
 FILLCELL_X32 FILLER_253_1552 ();
 FILLCELL_X32 FILLER_253_1584 ();
 FILLCELL_X32 FILLER_253_1616 ();
 FILLCELL_X32 FILLER_253_1648 ();
 FILLCELL_X32 FILLER_253_1680 ();
 FILLCELL_X32 FILLER_253_1712 ();
 FILLCELL_X32 FILLER_253_1744 ();
 FILLCELL_X32 FILLER_253_1776 ();
 FILLCELL_X32 FILLER_253_1808 ();
 FILLCELL_X32 FILLER_253_1840 ();
 FILLCELL_X32 FILLER_253_1872 ();
 FILLCELL_X32 FILLER_253_1904 ();
 FILLCELL_X32 FILLER_253_1936 ();
 FILLCELL_X32 FILLER_253_1968 ();
 FILLCELL_X32 FILLER_253_2000 ();
 FILLCELL_X32 FILLER_253_2032 ();
 FILLCELL_X32 FILLER_253_2064 ();
 FILLCELL_X16 FILLER_253_2096 ();
 FILLCELL_X2 FILLER_253_2112 ();
 FILLCELL_X1 FILLER_253_2114 ();
 FILLCELL_X32 FILLER_254_1 ();
 FILLCELL_X32 FILLER_254_33 ();
 FILLCELL_X32 FILLER_254_65 ();
 FILLCELL_X32 FILLER_254_97 ();
 FILLCELL_X32 FILLER_254_129 ();
 FILLCELL_X32 FILLER_254_161 ();
 FILLCELL_X32 FILLER_254_193 ();
 FILLCELL_X32 FILLER_254_225 ();
 FILLCELL_X32 FILLER_254_257 ();
 FILLCELL_X32 FILLER_254_289 ();
 FILLCELL_X32 FILLER_254_321 ();
 FILLCELL_X32 FILLER_254_353 ();
 FILLCELL_X32 FILLER_254_385 ();
 FILLCELL_X32 FILLER_254_417 ();
 FILLCELL_X32 FILLER_254_449 ();
 FILLCELL_X32 FILLER_254_481 ();
 FILLCELL_X32 FILLER_254_513 ();
 FILLCELL_X32 FILLER_254_545 ();
 FILLCELL_X32 FILLER_254_577 ();
 FILLCELL_X16 FILLER_254_609 ();
 FILLCELL_X4 FILLER_254_625 ();
 FILLCELL_X2 FILLER_254_629 ();
 FILLCELL_X32 FILLER_254_632 ();
 FILLCELL_X32 FILLER_254_664 ();
 FILLCELL_X32 FILLER_254_696 ();
 FILLCELL_X32 FILLER_254_728 ();
 FILLCELL_X32 FILLER_254_760 ();
 FILLCELL_X32 FILLER_254_792 ();
 FILLCELL_X32 FILLER_254_824 ();
 FILLCELL_X32 FILLER_254_856 ();
 FILLCELL_X32 FILLER_254_888 ();
 FILLCELL_X32 FILLER_254_920 ();
 FILLCELL_X32 FILLER_254_952 ();
 FILLCELL_X32 FILLER_254_984 ();
 FILLCELL_X32 FILLER_254_1016 ();
 FILLCELL_X32 FILLER_254_1048 ();
 FILLCELL_X32 FILLER_254_1080 ();
 FILLCELL_X32 FILLER_254_1112 ();
 FILLCELL_X32 FILLER_254_1144 ();
 FILLCELL_X32 FILLER_254_1176 ();
 FILLCELL_X32 FILLER_254_1208 ();
 FILLCELL_X32 FILLER_254_1240 ();
 FILLCELL_X32 FILLER_254_1272 ();
 FILLCELL_X32 FILLER_254_1304 ();
 FILLCELL_X32 FILLER_254_1336 ();
 FILLCELL_X32 FILLER_254_1368 ();
 FILLCELL_X32 FILLER_254_1400 ();
 FILLCELL_X32 FILLER_254_1432 ();
 FILLCELL_X32 FILLER_254_1464 ();
 FILLCELL_X32 FILLER_254_1496 ();
 FILLCELL_X32 FILLER_254_1528 ();
 FILLCELL_X32 FILLER_254_1560 ();
 FILLCELL_X32 FILLER_254_1592 ();
 FILLCELL_X32 FILLER_254_1624 ();
 FILLCELL_X32 FILLER_254_1656 ();
 FILLCELL_X32 FILLER_254_1688 ();
 FILLCELL_X32 FILLER_254_1720 ();
 FILLCELL_X32 FILLER_254_1752 ();
 FILLCELL_X32 FILLER_254_1784 ();
 FILLCELL_X32 FILLER_254_1816 ();
 FILLCELL_X32 FILLER_254_1848 ();
 FILLCELL_X8 FILLER_254_1880 ();
 FILLCELL_X4 FILLER_254_1888 ();
 FILLCELL_X2 FILLER_254_1892 ();
 FILLCELL_X32 FILLER_254_1895 ();
 FILLCELL_X32 FILLER_254_1927 ();
 FILLCELL_X32 FILLER_254_1959 ();
 FILLCELL_X32 FILLER_254_1991 ();
 FILLCELL_X32 FILLER_254_2023 ();
 FILLCELL_X32 FILLER_254_2055 ();
 FILLCELL_X16 FILLER_254_2087 ();
 FILLCELL_X8 FILLER_254_2103 ();
 FILLCELL_X4 FILLER_254_2111 ();
 FILLCELL_X32 FILLER_255_1 ();
 FILLCELL_X32 FILLER_255_33 ();
 FILLCELL_X32 FILLER_255_65 ();
 FILLCELL_X32 FILLER_255_97 ();
 FILLCELL_X32 FILLER_255_129 ();
 FILLCELL_X32 FILLER_255_161 ();
 FILLCELL_X32 FILLER_255_193 ();
 FILLCELL_X32 FILLER_255_225 ();
 FILLCELL_X32 FILLER_255_257 ();
 FILLCELL_X32 FILLER_255_289 ();
 FILLCELL_X32 FILLER_255_321 ();
 FILLCELL_X32 FILLER_255_353 ();
 FILLCELL_X32 FILLER_255_385 ();
 FILLCELL_X32 FILLER_255_417 ();
 FILLCELL_X32 FILLER_255_449 ();
 FILLCELL_X32 FILLER_255_481 ();
 FILLCELL_X32 FILLER_255_513 ();
 FILLCELL_X32 FILLER_255_545 ();
 FILLCELL_X32 FILLER_255_577 ();
 FILLCELL_X32 FILLER_255_609 ();
 FILLCELL_X32 FILLER_255_641 ();
 FILLCELL_X32 FILLER_255_673 ();
 FILLCELL_X32 FILLER_255_705 ();
 FILLCELL_X32 FILLER_255_737 ();
 FILLCELL_X32 FILLER_255_769 ();
 FILLCELL_X32 FILLER_255_801 ();
 FILLCELL_X32 FILLER_255_833 ();
 FILLCELL_X32 FILLER_255_865 ();
 FILLCELL_X32 FILLER_255_897 ();
 FILLCELL_X32 FILLER_255_929 ();
 FILLCELL_X32 FILLER_255_961 ();
 FILLCELL_X32 FILLER_255_993 ();
 FILLCELL_X32 FILLER_255_1025 ();
 FILLCELL_X32 FILLER_255_1057 ();
 FILLCELL_X32 FILLER_255_1089 ();
 FILLCELL_X32 FILLER_255_1121 ();
 FILLCELL_X32 FILLER_255_1153 ();
 FILLCELL_X32 FILLER_255_1185 ();
 FILLCELL_X32 FILLER_255_1217 ();
 FILLCELL_X8 FILLER_255_1249 ();
 FILLCELL_X4 FILLER_255_1257 ();
 FILLCELL_X2 FILLER_255_1261 ();
 FILLCELL_X32 FILLER_255_1264 ();
 FILLCELL_X32 FILLER_255_1296 ();
 FILLCELL_X32 FILLER_255_1328 ();
 FILLCELL_X32 FILLER_255_1360 ();
 FILLCELL_X32 FILLER_255_1392 ();
 FILLCELL_X32 FILLER_255_1424 ();
 FILLCELL_X32 FILLER_255_1456 ();
 FILLCELL_X32 FILLER_255_1488 ();
 FILLCELL_X32 FILLER_255_1520 ();
 FILLCELL_X32 FILLER_255_1552 ();
 FILLCELL_X32 FILLER_255_1584 ();
 FILLCELL_X32 FILLER_255_1616 ();
 FILLCELL_X32 FILLER_255_1648 ();
 FILLCELL_X32 FILLER_255_1680 ();
 FILLCELL_X32 FILLER_255_1712 ();
 FILLCELL_X32 FILLER_255_1744 ();
 FILLCELL_X32 FILLER_255_1776 ();
 FILLCELL_X32 FILLER_255_1808 ();
 FILLCELL_X32 FILLER_255_1840 ();
 FILLCELL_X32 FILLER_255_1872 ();
 FILLCELL_X32 FILLER_255_1904 ();
 FILLCELL_X32 FILLER_255_1936 ();
 FILLCELL_X32 FILLER_255_1968 ();
 FILLCELL_X32 FILLER_255_2000 ();
 FILLCELL_X32 FILLER_255_2032 ();
 FILLCELL_X32 FILLER_255_2064 ();
 FILLCELL_X16 FILLER_255_2096 ();
 FILLCELL_X2 FILLER_255_2112 ();
 FILLCELL_X1 FILLER_255_2114 ();
 FILLCELL_X32 FILLER_256_1 ();
 FILLCELL_X32 FILLER_256_33 ();
 FILLCELL_X32 FILLER_256_65 ();
 FILLCELL_X32 FILLER_256_97 ();
 FILLCELL_X32 FILLER_256_129 ();
 FILLCELL_X32 FILLER_256_161 ();
 FILLCELL_X32 FILLER_256_193 ();
 FILLCELL_X32 FILLER_256_225 ();
 FILLCELL_X32 FILLER_256_257 ();
 FILLCELL_X32 FILLER_256_289 ();
 FILLCELL_X32 FILLER_256_321 ();
 FILLCELL_X32 FILLER_256_353 ();
 FILLCELL_X32 FILLER_256_385 ();
 FILLCELL_X32 FILLER_256_417 ();
 FILLCELL_X32 FILLER_256_449 ();
 FILLCELL_X32 FILLER_256_481 ();
 FILLCELL_X32 FILLER_256_513 ();
 FILLCELL_X32 FILLER_256_545 ();
 FILLCELL_X32 FILLER_256_577 ();
 FILLCELL_X16 FILLER_256_609 ();
 FILLCELL_X4 FILLER_256_625 ();
 FILLCELL_X2 FILLER_256_629 ();
 FILLCELL_X32 FILLER_256_632 ();
 FILLCELL_X32 FILLER_256_664 ();
 FILLCELL_X32 FILLER_256_696 ();
 FILLCELL_X32 FILLER_256_728 ();
 FILLCELL_X32 FILLER_256_760 ();
 FILLCELL_X32 FILLER_256_792 ();
 FILLCELL_X32 FILLER_256_824 ();
 FILLCELL_X32 FILLER_256_856 ();
 FILLCELL_X32 FILLER_256_888 ();
 FILLCELL_X32 FILLER_256_920 ();
 FILLCELL_X32 FILLER_256_952 ();
 FILLCELL_X32 FILLER_256_984 ();
 FILLCELL_X32 FILLER_256_1016 ();
 FILLCELL_X32 FILLER_256_1048 ();
 FILLCELL_X32 FILLER_256_1080 ();
 FILLCELL_X32 FILLER_256_1112 ();
 FILLCELL_X32 FILLER_256_1144 ();
 FILLCELL_X32 FILLER_256_1176 ();
 FILLCELL_X32 FILLER_256_1208 ();
 FILLCELL_X32 FILLER_256_1240 ();
 FILLCELL_X32 FILLER_256_1272 ();
 FILLCELL_X32 FILLER_256_1304 ();
 FILLCELL_X32 FILLER_256_1336 ();
 FILLCELL_X32 FILLER_256_1368 ();
 FILLCELL_X32 FILLER_256_1400 ();
 FILLCELL_X32 FILLER_256_1432 ();
 FILLCELL_X32 FILLER_256_1464 ();
 FILLCELL_X32 FILLER_256_1496 ();
 FILLCELL_X32 FILLER_256_1528 ();
 FILLCELL_X32 FILLER_256_1560 ();
 FILLCELL_X32 FILLER_256_1592 ();
 FILLCELL_X32 FILLER_256_1624 ();
 FILLCELL_X32 FILLER_256_1656 ();
 FILLCELL_X32 FILLER_256_1688 ();
 FILLCELL_X32 FILLER_256_1720 ();
 FILLCELL_X32 FILLER_256_1752 ();
 FILLCELL_X32 FILLER_256_1784 ();
 FILLCELL_X32 FILLER_256_1816 ();
 FILLCELL_X32 FILLER_256_1848 ();
 FILLCELL_X8 FILLER_256_1880 ();
 FILLCELL_X4 FILLER_256_1888 ();
 FILLCELL_X2 FILLER_256_1892 ();
 FILLCELL_X32 FILLER_256_1895 ();
 FILLCELL_X32 FILLER_256_1927 ();
 FILLCELL_X32 FILLER_256_1959 ();
 FILLCELL_X32 FILLER_256_1991 ();
 FILLCELL_X32 FILLER_256_2023 ();
 FILLCELL_X32 FILLER_256_2055 ();
 FILLCELL_X16 FILLER_256_2087 ();
 FILLCELL_X8 FILLER_256_2103 ();
 FILLCELL_X4 FILLER_256_2111 ();
 FILLCELL_X32 FILLER_257_1 ();
 FILLCELL_X32 FILLER_257_33 ();
 FILLCELL_X32 FILLER_257_65 ();
 FILLCELL_X32 FILLER_257_97 ();
 FILLCELL_X32 FILLER_257_129 ();
 FILLCELL_X32 FILLER_257_161 ();
 FILLCELL_X32 FILLER_257_193 ();
 FILLCELL_X32 FILLER_257_225 ();
 FILLCELL_X32 FILLER_257_257 ();
 FILLCELL_X32 FILLER_257_289 ();
 FILLCELL_X32 FILLER_257_321 ();
 FILLCELL_X32 FILLER_257_353 ();
 FILLCELL_X32 FILLER_257_385 ();
 FILLCELL_X32 FILLER_257_417 ();
 FILLCELL_X32 FILLER_257_449 ();
 FILLCELL_X32 FILLER_257_481 ();
 FILLCELL_X32 FILLER_257_513 ();
 FILLCELL_X32 FILLER_257_545 ();
 FILLCELL_X32 FILLER_257_577 ();
 FILLCELL_X32 FILLER_257_609 ();
 FILLCELL_X32 FILLER_257_641 ();
 FILLCELL_X32 FILLER_257_673 ();
 FILLCELL_X32 FILLER_257_705 ();
 FILLCELL_X32 FILLER_257_737 ();
 FILLCELL_X32 FILLER_257_769 ();
 FILLCELL_X32 FILLER_257_801 ();
 FILLCELL_X32 FILLER_257_833 ();
 FILLCELL_X32 FILLER_257_865 ();
 FILLCELL_X32 FILLER_257_897 ();
 FILLCELL_X32 FILLER_257_929 ();
 FILLCELL_X32 FILLER_257_961 ();
 FILLCELL_X32 FILLER_257_993 ();
 FILLCELL_X32 FILLER_257_1025 ();
 FILLCELL_X32 FILLER_257_1057 ();
 FILLCELL_X32 FILLER_257_1089 ();
 FILLCELL_X32 FILLER_257_1121 ();
 FILLCELL_X32 FILLER_257_1153 ();
 FILLCELL_X32 FILLER_257_1185 ();
 FILLCELL_X32 FILLER_257_1217 ();
 FILLCELL_X8 FILLER_257_1249 ();
 FILLCELL_X4 FILLER_257_1257 ();
 FILLCELL_X2 FILLER_257_1261 ();
 FILLCELL_X32 FILLER_257_1264 ();
 FILLCELL_X32 FILLER_257_1296 ();
 FILLCELL_X32 FILLER_257_1328 ();
 FILLCELL_X32 FILLER_257_1360 ();
 FILLCELL_X32 FILLER_257_1392 ();
 FILLCELL_X32 FILLER_257_1424 ();
 FILLCELL_X32 FILLER_257_1456 ();
 FILLCELL_X32 FILLER_257_1488 ();
 FILLCELL_X32 FILLER_257_1520 ();
 FILLCELL_X32 FILLER_257_1552 ();
 FILLCELL_X32 FILLER_257_1584 ();
 FILLCELL_X32 FILLER_257_1616 ();
 FILLCELL_X32 FILLER_257_1648 ();
 FILLCELL_X32 FILLER_257_1680 ();
 FILLCELL_X32 FILLER_257_1712 ();
 FILLCELL_X32 FILLER_257_1744 ();
 FILLCELL_X32 FILLER_257_1776 ();
 FILLCELL_X32 FILLER_257_1808 ();
 FILLCELL_X32 FILLER_257_1840 ();
 FILLCELL_X32 FILLER_257_1872 ();
 FILLCELL_X32 FILLER_257_1904 ();
 FILLCELL_X32 FILLER_257_1936 ();
 FILLCELL_X32 FILLER_257_1968 ();
 FILLCELL_X32 FILLER_257_2000 ();
 FILLCELL_X32 FILLER_257_2032 ();
 FILLCELL_X32 FILLER_257_2064 ();
 FILLCELL_X16 FILLER_257_2096 ();
 FILLCELL_X2 FILLER_257_2112 ();
 FILLCELL_X1 FILLER_257_2114 ();
 FILLCELL_X32 FILLER_258_1 ();
 FILLCELL_X32 FILLER_258_33 ();
 FILLCELL_X32 FILLER_258_65 ();
 FILLCELL_X32 FILLER_258_97 ();
 FILLCELL_X32 FILLER_258_129 ();
 FILLCELL_X32 FILLER_258_161 ();
 FILLCELL_X32 FILLER_258_193 ();
 FILLCELL_X32 FILLER_258_225 ();
 FILLCELL_X32 FILLER_258_257 ();
 FILLCELL_X32 FILLER_258_289 ();
 FILLCELL_X32 FILLER_258_321 ();
 FILLCELL_X32 FILLER_258_353 ();
 FILLCELL_X32 FILLER_258_385 ();
 FILLCELL_X32 FILLER_258_417 ();
 FILLCELL_X32 FILLER_258_449 ();
 FILLCELL_X32 FILLER_258_481 ();
 FILLCELL_X32 FILLER_258_513 ();
 FILLCELL_X32 FILLER_258_545 ();
 FILLCELL_X32 FILLER_258_577 ();
 FILLCELL_X16 FILLER_258_609 ();
 FILLCELL_X4 FILLER_258_625 ();
 FILLCELL_X2 FILLER_258_629 ();
 FILLCELL_X32 FILLER_258_632 ();
 FILLCELL_X32 FILLER_258_664 ();
 FILLCELL_X32 FILLER_258_696 ();
 FILLCELL_X32 FILLER_258_728 ();
 FILLCELL_X32 FILLER_258_760 ();
 FILLCELL_X32 FILLER_258_792 ();
 FILLCELL_X32 FILLER_258_824 ();
 FILLCELL_X32 FILLER_258_856 ();
 FILLCELL_X32 FILLER_258_888 ();
 FILLCELL_X32 FILLER_258_920 ();
 FILLCELL_X32 FILLER_258_952 ();
 FILLCELL_X32 FILLER_258_984 ();
 FILLCELL_X32 FILLER_258_1016 ();
 FILLCELL_X32 FILLER_258_1048 ();
 FILLCELL_X32 FILLER_258_1080 ();
 FILLCELL_X32 FILLER_258_1112 ();
 FILLCELL_X32 FILLER_258_1144 ();
 FILLCELL_X32 FILLER_258_1176 ();
 FILLCELL_X32 FILLER_258_1208 ();
 FILLCELL_X32 FILLER_258_1240 ();
 FILLCELL_X32 FILLER_258_1272 ();
 FILLCELL_X32 FILLER_258_1304 ();
 FILLCELL_X32 FILLER_258_1336 ();
 FILLCELL_X32 FILLER_258_1368 ();
 FILLCELL_X32 FILLER_258_1400 ();
 FILLCELL_X32 FILLER_258_1432 ();
 FILLCELL_X32 FILLER_258_1464 ();
 FILLCELL_X32 FILLER_258_1496 ();
 FILLCELL_X32 FILLER_258_1528 ();
 FILLCELL_X32 FILLER_258_1560 ();
 FILLCELL_X32 FILLER_258_1592 ();
 FILLCELL_X32 FILLER_258_1624 ();
 FILLCELL_X32 FILLER_258_1656 ();
 FILLCELL_X32 FILLER_258_1688 ();
 FILLCELL_X32 FILLER_258_1720 ();
 FILLCELL_X32 FILLER_258_1752 ();
 FILLCELL_X32 FILLER_258_1784 ();
 FILLCELL_X32 FILLER_258_1816 ();
 FILLCELL_X32 FILLER_258_1848 ();
 FILLCELL_X8 FILLER_258_1880 ();
 FILLCELL_X4 FILLER_258_1888 ();
 FILLCELL_X2 FILLER_258_1892 ();
 FILLCELL_X32 FILLER_258_1895 ();
 FILLCELL_X32 FILLER_258_1927 ();
 FILLCELL_X32 FILLER_258_1959 ();
 FILLCELL_X32 FILLER_258_1991 ();
 FILLCELL_X32 FILLER_258_2023 ();
 FILLCELL_X32 FILLER_258_2055 ();
 FILLCELL_X16 FILLER_258_2087 ();
 FILLCELL_X8 FILLER_258_2103 ();
 FILLCELL_X4 FILLER_258_2111 ();
 FILLCELL_X32 FILLER_259_1 ();
 FILLCELL_X32 FILLER_259_33 ();
 FILLCELL_X32 FILLER_259_65 ();
 FILLCELL_X32 FILLER_259_97 ();
 FILLCELL_X32 FILLER_259_129 ();
 FILLCELL_X32 FILLER_259_161 ();
 FILLCELL_X32 FILLER_259_193 ();
 FILLCELL_X32 FILLER_259_225 ();
 FILLCELL_X32 FILLER_259_257 ();
 FILLCELL_X32 FILLER_259_289 ();
 FILLCELL_X32 FILLER_259_321 ();
 FILLCELL_X32 FILLER_259_353 ();
 FILLCELL_X32 FILLER_259_385 ();
 FILLCELL_X32 FILLER_259_417 ();
 FILLCELL_X32 FILLER_259_449 ();
 FILLCELL_X32 FILLER_259_481 ();
 FILLCELL_X32 FILLER_259_513 ();
 FILLCELL_X32 FILLER_259_545 ();
 FILLCELL_X32 FILLER_259_577 ();
 FILLCELL_X32 FILLER_259_609 ();
 FILLCELL_X32 FILLER_259_641 ();
 FILLCELL_X32 FILLER_259_673 ();
 FILLCELL_X32 FILLER_259_705 ();
 FILLCELL_X32 FILLER_259_737 ();
 FILLCELL_X32 FILLER_259_769 ();
 FILLCELL_X32 FILLER_259_801 ();
 FILLCELL_X32 FILLER_259_833 ();
 FILLCELL_X32 FILLER_259_865 ();
 FILLCELL_X32 FILLER_259_897 ();
 FILLCELL_X32 FILLER_259_929 ();
 FILLCELL_X32 FILLER_259_961 ();
 FILLCELL_X32 FILLER_259_993 ();
 FILLCELL_X32 FILLER_259_1025 ();
 FILLCELL_X32 FILLER_259_1057 ();
 FILLCELL_X32 FILLER_259_1089 ();
 FILLCELL_X32 FILLER_259_1121 ();
 FILLCELL_X32 FILLER_259_1153 ();
 FILLCELL_X32 FILLER_259_1185 ();
 FILLCELL_X32 FILLER_259_1217 ();
 FILLCELL_X8 FILLER_259_1249 ();
 FILLCELL_X4 FILLER_259_1257 ();
 FILLCELL_X2 FILLER_259_1261 ();
 FILLCELL_X32 FILLER_259_1264 ();
 FILLCELL_X32 FILLER_259_1296 ();
 FILLCELL_X32 FILLER_259_1328 ();
 FILLCELL_X32 FILLER_259_1360 ();
 FILLCELL_X32 FILLER_259_1392 ();
 FILLCELL_X32 FILLER_259_1424 ();
 FILLCELL_X32 FILLER_259_1456 ();
 FILLCELL_X32 FILLER_259_1488 ();
 FILLCELL_X32 FILLER_259_1520 ();
 FILLCELL_X32 FILLER_259_1552 ();
 FILLCELL_X32 FILLER_259_1584 ();
 FILLCELL_X32 FILLER_259_1616 ();
 FILLCELL_X32 FILLER_259_1648 ();
 FILLCELL_X32 FILLER_259_1680 ();
 FILLCELL_X32 FILLER_259_1712 ();
 FILLCELL_X32 FILLER_259_1744 ();
 FILLCELL_X32 FILLER_259_1776 ();
 FILLCELL_X32 FILLER_259_1808 ();
 FILLCELL_X32 FILLER_259_1840 ();
 FILLCELL_X32 FILLER_259_1872 ();
 FILLCELL_X32 FILLER_259_1904 ();
 FILLCELL_X32 FILLER_259_1936 ();
 FILLCELL_X32 FILLER_259_1968 ();
 FILLCELL_X32 FILLER_259_2000 ();
 FILLCELL_X32 FILLER_259_2032 ();
 FILLCELL_X32 FILLER_259_2064 ();
 FILLCELL_X16 FILLER_259_2096 ();
 FILLCELL_X2 FILLER_259_2112 ();
 FILLCELL_X1 FILLER_259_2114 ();
 FILLCELL_X32 FILLER_260_1 ();
 FILLCELL_X32 FILLER_260_33 ();
 FILLCELL_X32 FILLER_260_65 ();
 FILLCELL_X32 FILLER_260_97 ();
 FILLCELL_X32 FILLER_260_129 ();
 FILLCELL_X32 FILLER_260_161 ();
 FILLCELL_X32 FILLER_260_193 ();
 FILLCELL_X32 FILLER_260_225 ();
 FILLCELL_X32 FILLER_260_257 ();
 FILLCELL_X32 FILLER_260_289 ();
 FILLCELL_X32 FILLER_260_321 ();
 FILLCELL_X32 FILLER_260_353 ();
 FILLCELL_X32 FILLER_260_385 ();
 FILLCELL_X32 FILLER_260_417 ();
 FILLCELL_X32 FILLER_260_449 ();
 FILLCELL_X32 FILLER_260_481 ();
 FILLCELL_X32 FILLER_260_513 ();
 FILLCELL_X32 FILLER_260_545 ();
 FILLCELL_X32 FILLER_260_577 ();
 FILLCELL_X16 FILLER_260_609 ();
 FILLCELL_X4 FILLER_260_625 ();
 FILLCELL_X2 FILLER_260_629 ();
 FILLCELL_X32 FILLER_260_632 ();
 FILLCELL_X32 FILLER_260_664 ();
 FILLCELL_X32 FILLER_260_696 ();
 FILLCELL_X32 FILLER_260_728 ();
 FILLCELL_X32 FILLER_260_760 ();
 FILLCELL_X32 FILLER_260_792 ();
 FILLCELL_X32 FILLER_260_824 ();
 FILLCELL_X32 FILLER_260_856 ();
 FILLCELL_X32 FILLER_260_888 ();
 FILLCELL_X32 FILLER_260_920 ();
 FILLCELL_X32 FILLER_260_952 ();
 FILLCELL_X32 FILLER_260_984 ();
 FILLCELL_X32 FILLER_260_1016 ();
 FILLCELL_X32 FILLER_260_1048 ();
 FILLCELL_X32 FILLER_260_1080 ();
 FILLCELL_X32 FILLER_260_1112 ();
 FILLCELL_X32 FILLER_260_1144 ();
 FILLCELL_X32 FILLER_260_1176 ();
 FILLCELL_X32 FILLER_260_1208 ();
 FILLCELL_X32 FILLER_260_1240 ();
 FILLCELL_X32 FILLER_260_1272 ();
 FILLCELL_X32 FILLER_260_1304 ();
 FILLCELL_X32 FILLER_260_1336 ();
 FILLCELL_X32 FILLER_260_1368 ();
 FILLCELL_X32 FILLER_260_1400 ();
 FILLCELL_X32 FILLER_260_1432 ();
 FILLCELL_X32 FILLER_260_1464 ();
 FILLCELL_X32 FILLER_260_1496 ();
 FILLCELL_X32 FILLER_260_1528 ();
 FILLCELL_X32 FILLER_260_1560 ();
 FILLCELL_X32 FILLER_260_1592 ();
 FILLCELL_X32 FILLER_260_1624 ();
 FILLCELL_X32 FILLER_260_1656 ();
 FILLCELL_X32 FILLER_260_1688 ();
 FILLCELL_X32 FILLER_260_1720 ();
 FILLCELL_X32 FILLER_260_1752 ();
 FILLCELL_X32 FILLER_260_1784 ();
 FILLCELL_X32 FILLER_260_1816 ();
 FILLCELL_X32 FILLER_260_1848 ();
 FILLCELL_X8 FILLER_260_1880 ();
 FILLCELL_X4 FILLER_260_1888 ();
 FILLCELL_X2 FILLER_260_1892 ();
 FILLCELL_X32 FILLER_260_1895 ();
 FILLCELL_X32 FILLER_260_1927 ();
 FILLCELL_X32 FILLER_260_1959 ();
 FILLCELL_X32 FILLER_260_1991 ();
 FILLCELL_X32 FILLER_260_2023 ();
 FILLCELL_X32 FILLER_260_2055 ();
 FILLCELL_X16 FILLER_260_2087 ();
 FILLCELL_X8 FILLER_260_2103 ();
 FILLCELL_X4 FILLER_260_2111 ();
 FILLCELL_X32 FILLER_261_1 ();
 FILLCELL_X32 FILLER_261_33 ();
 FILLCELL_X32 FILLER_261_65 ();
 FILLCELL_X32 FILLER_261_97 ();
 FILLCELL_X32 FILLER_261_129 ();
 FILLCELL_X32 FILLER_261_161 ();
 FILLCELL_X32 FILLER_261_193 ();
 FILLCELL_X32 FILLER_261_225 ();
 FILLCELL_X32 FILLER_261_257 ();
 FILLCELL_X32 FILLER_261_289 ();
 FILLCELL_X32 FILLER_261_321 ();
 FILLCELL_X32 FILLER_261_353 ();
 FILLCELL_X32 FILLER_261_385 ();
 FILLCELL_X32 FILLER_261_417 ();
 FILLCELL_X32 FILLER_261_449 ();
 FILLCELL_X32 FILLER_261_481 ();
 FILLCELL_X32 FILLER_261_513 ();
 FILLCELL_X32 FILLER_261_545 ();
 FILLCELL_X32 FILLER_261_577 ();
 FILLCELL_X32 FILLER_261_609 ();
 FILLCELL_X32 FILLER_261_641 ();
 FILLCELL_X32 FILLER_261_673 ();
 FILLCELL_X32 FILLER_261_705 ();
 FILLCELL_X32 FILLER_261_737 ();
 FILLCELL_X32 FILLER_261_769 ();
 FILLCELL_X32 FILLER_261_801 ();
 FILLCELL_X32 FILLER_261_833 ();
 FILLCELL_X32 FILLER_261_865 ();
 FILLCELL_X32 FILLER_261_897 ();
 FILLCELL_X32 FILLER_261_929 ();
 FILLCELL_X32 FILLER_261_961 ();
 FILLCELL_X32 FILLER_261_993 ();
 FILLCELL_X32 FILLER_261_1025 ();
 FILLCELL_X32 FILLER_261_1057 ();
 FILLCELL_X32 FILLER_261_1089 ();
 FILLCELL_X32 FILLER_261_1121 ();
 FILLCELL_X32 FILLER_261_1153 ();
 FILLCELL_X32 FILLER_261_1185 ();
 FILLCELL_X32 FILLER_261_1217 ();
 FILLCELL_X8 FILLER_261_1249 ();
 FILLCELL_X4 FILLER_261_1257 ();
 FILLCELL_X2 FILLER_261_1261 ();
 FILLCELL_X32 FILLER_261_1264 ();
 FILLCELL_X32 FILLER_261_1296 ();
 FILLCELL_X32 FILLER_261_1328 ();
 FILLCELL_X32 FILLER_261_1360 ();
 FILLCELL_X32 FILLER_261_1392 ();
 FILLCELL_X32 FILLER_261_1424 ();
 FILLCELL_X32 FILLER_261_1456 ();
 FILLCELL_X32 FILLER_261_1488 ();
 FILLCELL_X32 FILLER_261_1520 ();
 FILLCELL_X32 FILLER_261_1552 ();
 FILLCELL_X32 FILLER_261_1584 ();
 FILLCELL_X32 FILLER_261_1616 ();
 FILLCELL_X32 FILLER_261_1648 ();
 FILLCELL_X32 FILLER_261_1680 ();
 FILLCELL_X32 FILLER_261_1712 ();
 FILLCELL_X32 FILLER_261_1744 ();
 FILLCELL_X32 FILLER_261_1776 ();
 FILLCELL_X32 FILLER_261_1808 ();
 FILLCELL_X32 FILLER_261_1840 ();
 FILLCELL_X32 FILLER_261_1872 ();
 FILLCELL_X32 FILLER_261_1904 ();
 FILLCELL_X32 FILLER_261_1936 ();
 FILLCELL_X32 FILLER_261_1968 ();
 FILLCELL_X32 FILLER_261_2000 ();
 FILLCELL_X32 FILLER_261_2032 ();
 FILLCELL_X32 FILLER_261_2064 ();
 FILLCELL_X16 FILLER_261_2096 ();
 FILLCELL_X2 FILLER_261_2112 ();
 FILLCELL_X1 FILLER_261_2114 ();
 FILLCELL_X32 FILLER_262_1 ();
 FILLCELL_X32 FILLER_262_33 ();
 FILLCELL_X32 FILLER_262_65 ();
 FILLCELL_X32 FILLER_262_97 ();
 FILLCELL_X32 FILLER_262_129 ();
 FILLCELL_X32 FILLER_262_161 ();
 FILLCELL_X32 FILLER_262_193 ();
 FILLCELL_X32 FILLER_262_225 ();
 FILLCELL_X32 FILLER_262_257 ();
 FILLCELL_X32 FILLER_262_289 ();
 FILLCELL_X32 FILLER_262_321 ();
 FILLCELL_X32 FILLER_262_353 ();
 FILLCELL_X32 FILLER_262_385 ();
 FILLCELL_X32 FILLER_262_417 ();
 FILLCELL_X32 FILLER_262_449 ();
 FILLCELL_X32 FILLER_262_481 ();
 FILLCELL_X32 FILLER_262_513 ();
 FILLCELL_X32 FILLER_262_545 ();
 FILLCELL_X32 FILLER_262_577 ();
 FILLCELL_X16 FILLER_262_609 ();
 FILLCELL_X4 FILLER_262_625 ();
 FILLCELL_X2 FILLER_262_629 ();
 FILLCELL_X32 FILLER_262_632 ();
 FILLCELL_X32 FILLER_262_664 ();
 FILLCELL_X32 FILLER_262_696 ();
 FILLCELL_X32 FILLER_262_728 ();
 FILLCELL_X32 FILLER_262_760 ();
 FILLCELL_X32 FILLER_262_792 ();
 FILLCELL_X32 FILLER_262_824 ();
 FILLCELL_X32 FILLER_262_856 ();
 FILLCELL_X32 FILLER_262_888 ();
 FILLCELL_X32 FILLER_262_920 ();
 FILLCELL_X32 FILLER_262_952 ();
 FILLCELL_X32 FILLER_262_984 ();
 FILLCELL_X32 FILLER_262_1016 ();
 FILLCELL_X32 FILLER_262_1048 ();
 FILLCELL_X32 FILLER_262_1080 ();
 FILLCELL_X32 FILLER_262_1112 ();
 FILLCELL_X32 FILLER_262_1144 ();
 FILLCELL_X32 FILLER_262_1176 ();
 FILLCELL_X32 FILLER_262_1208 ();
 FILLCELL_X32 FILLER_262_1240 ();
 FILLCELL_X32 FILLER_262_1272 ();
 FILLCELL_X32 FILLER_262_1304 ();
 FILLCELL_X32 FILLER_262_1336 ();
 FILLCELL_X32 FILLER_262_1368 ();
 FILLCELL_X32 FILLER_262_1400 ();
 FILLCELL_X32 FILLER_262_1432 ();
 FILLCELL_X32 FILLER_262_1464 ();
 FILLCELL_X32 FILLER_262_1496 ();
 FILLCELL_X32 FILLER_262_1528 ();
 FILLCELL_X32 FILLER_262_1560 ();
 FILLCELL_X32 FILLER_262_1592 ();
 FILLCELL_X32 FILLER_262_1624 ();
 FILLCELL_X32 FILLER_262_1656 ();
 FILLCELL_X32 FILLER_262_1688 ();
 FILLCELL_X32 FILLER_262_1720 ();
 FILLCELL_X32 FILLER_262_1752 ();
 FILLCELL_X32 FILLER_262_1784 ();
 FILLCELL_X32 FILLER_262_1816 ();
 FILLCELL_X32 FILLER_262_1848 ();
 FILLCELL_X8 FILLER_262_1880 ();
 FILLCELL_X4 FILLER_262_1888 ();
 FILLCELL_X2 FILLER_262_1892 ();
 FILLCELL_X32 FILLER_262_1895 ();
 FILLCELL_X32 FILLER_262_1927 ();
 FILLCELL_X32 FILLER_262_1959 ();
 FILLCELL_X32 FILLER_262_1991 ();
 FILLCELL_X32 FILLER_262_2023 ();
 FILLCELL_X32 FILLER_262_2055 ();
 FILLCELL_X16 FILLER_262_2087 ();
 FILLCELL_X8 FILLER_262_2103 ();
 FILLCELL_X4 FILLER_262_2111 ();
 FILLCELL_X32 FILLER_263_1 ();
 FILLCELL_X32 FILLER_263_33 ();
 FILLCELL_X32 FILLER_263_65 ();
 FILLCELL_X32 FILLER_263_97 ();
 FILLCELL_X32 FILLER_263_129 ();
 FILLCELL_X32 FILLER_263_161 ();
 FILLCELL_X32 FILLER_263_193 ();
 FILLCELL_X32 FILLER_263_225 ();
 FILLCELL_X32 FILLER_263_257 ();
 FILLCELL_X32 FILLER_263_289 ();
 FILLCELL_X32 FILLER_263_321 ();
 FILLCELL_X32 FILLER_263_353 ();
 FILLCELL_X32 FILLER_263_385 ();
 FILLCELL_X32 FILLER_263_417 ();
 FILLCELL_X32 FILLER_263_449 ();
 FILLCELL_X32 FILLER_263_481 ();
 FILLCELL_X32 FILLER_263_513 ();
 FILLCELL_X32 FILLER_263_545 ();
 FILLCELL_X32 FILLER_263_577 ();
 FILLCELL_X32 FILLER_263_609 ();
 FILLCELL_X32 FILLER_263_641 ();
 FILLCELL_X32 FILLER_263_673 ();
 FILLCELL_X32 FILLER_263_705 ();
 FILLCELL_X32 FILLER_263_737 ();
 FILLCELL_X32 FILLER_263_769 ();
 FILLCELL_X32 FILLER_263_801 ();
 FILLCELL_X32 FILLER_263_833 ();
 FILLCELL_X32 FILLER_263_865 ();
 FILLCELL_X32 FILLER_263_897 ();
 FILLCELL_X32 FILLER_263_929 ();
 FILLCELL_X32 FILLER_263_961 ();
 FILLCELL_X32 FILLER_263_993 ();
 FILLCELL_X32 FILLER_263_1025 ();
 FILLCELL_X32 FILLER_263_1057 ();
 FILLCELL_X32 FILLER_263_1089 ();
 FILLCELL_X32 FILLER_263_1121 ();
 FILLCELL_X32 FILLER_263_1153 ();
 FILLCELL_X32 FILLER_263_1185 ();
 FILLCELL_X32 FILLER_263_1217 ();
 FILLCELL_X8 FILLER_263_1249 ();
 FILLCELL_X4 FILLER_263_1257 ();
 FILLCELL_X2 FILLER_263_1261 ();
 FILLCELL_X32 FILLER_263_1264 ();
 FILLCELL_X32 FILLER_263_1296 ();
 FILLCELL_X32 FILLER_263_1328 ();
 FILLCELL_X32 FILLER_263_1360 ();
 FILLCELL_X32 FILLER_263_1392 ();
 FILLCELL_X32 FILLER_263_1424 ();
 FILLCELL_X32 FILLER_263_1456 ();
 FILLCELL_X32 FILLER_263_1488 ();
 FILLCELL_X32 FILLER_263_1520 ();
 FILLCELL_X32 FILLER_263_1552 ();
 FILLCELL_X32 FILLER_263_1584 ();
 FILLCELL_X32 FILLER_263_1616 ();
 FILLCELL_X32 FILLER_263_1648 ();
 FILLCELL_X32 FILLER_263_1680 ();
 FILLCELL_X32 FILLER_263_1712 ();
 FILLCELL_X32 FILLER_263_1744 ();
 FILLCELL_X32 FILLER_263_1776 ();
 FILLCELL_X32 FILLER_263_1808 ();
 FILLCELL_X32 FILLER_263_1840 ();
 FILLCELL_X32 FILLER_263_1872 ();
 FILLCELL_X32 FILLER_263_1904 ();
 FILLCELL_X32 FILLER_263_1936 ();
 FILLCELL_X32 FILLER_263_1968 ();
 FILLCELL_X32 FILLER_263_2000 ();
 FILLCELL_X32 FILLER_263_2032 ();
 FILLCELL_X32 FILLER_263_2064 ();
 FILLCELL_X16 FILLER_263_2096 ();
 FILLCELL_X2 FILLER_263_2112 ();
 FILLCELL_X1 FILLER_263_2114 ();
 FILLCELL_X32 FILLER_264_1 ();
 FILLCELL_X32 FILLER_264_33 ();
 FILLCELL_X32 FILLER_264_65 ();
 FILLCELL_X32 FILLER_264_97 ();
 FILLCELL_X32 FILLER_264_129 ();
 FILLCELL_X32 FILLER_264_161 ();
 FILLCELL_X32 FILLER_264_193 ();
 FILLCELL_X32 FILLER_264_225 ();
 FILLCELL_X32 FILLER_264_257 ();
 FILLCELL_X32 FILLER_264_289 ();
 FILLCELL_X32 FILLER_264_321 ();
 FILLCELL_X32 FILLER_264_353 ();
 FILLCELL_X32 FILLER_264_385 ();
 FILLCELL_X32 FILLER_264_417 ();
 FILLCELL_X32 FILLER_264_449 ();
 FILLCELL_X32 FILLER_264_481 ();
 FILLCELL_X32 FILLER_264_513 ();
 FILLCELL_X32 FILLER_264_545 ();
 FILLCELL_X32 FILLER_264_577 ();
 FILLCELL_X16 FILLER_264_609 ();
 FILLCELL_X4 FILLER_264_625 ();
 FILLCELL_X2 FILLER_264_629 ();
 FILLCELL_X32 FILLER_264_632 ();
 FILLCELL_X32 FILLER_264_664 ();
 FILLCELL_X32 FILLER_264_696 ();
 FILLCELL_X32 FILLER_264_728 ();
 FILLCELL_X32 FILLER_264_760 ();
 FILLCELL_X32 FILLER_264_792 ();
 FILLCELL_X32 FILLER_264_824 ();
 FILLCELL_X32 FILLER_264_856 ();
 FILLCELL_X32 FILLER_264_888 ();
 FILLCELL_X32 FILLER_264_920 ();
 FILLCELL_X32 FILLER_264_952 ();
 FILLCELL_X32 FILLER_264_984 ();
 FILLCELL_X32 FILLER_264_1016 ();
 FILLCELL_X32 FILLER_264_1048 ();
 FILLCELL_X32 FILLER_264_1080 ();
 FILLCELL_X32 FILLER_264_1112 ();
 FILLCELL_X32 FILLER_264_1144 ();
 FILLCELL_X32 FILLER_264_1176 ();
 FILLCELL_X32 FILLER_264_1208 ();
 FILLCELL_X32 FILLER_264_1240 ();
 FILLCELL_X32 FILLER_264_1272 ();
 FILLCELL_X32 FILLER_264_1304 ();
 FILLCELL_X32 FILLER_264_1336 ();
 FILLCELL_X32 FILLER_264_1368 ();
 FILLCELL_X32 FILLER_264_1400 ();
 FILLCELL_X32 FILLER_264_1432 ();
 FILLCELL_X32 FILLER_264_1464 ();
 FILLCELL_X32 FILLER_264_1496 ();
 FILLCELL_X32 FILLER_264_1528 ();
 FILLCELL_X32 FILLER_264_1560 ();
 FILLCELL_X32 FILLER_264_1592 ();
 FILLCELL_X32 FILLER_264_1624 ();
 FILLCELL_X32 FILLER_264_1656 ();
 FILLCELL_X32 FILLER_264_1688 ();
 FILLCELL_X32 FILLER_264_1720 ();
 FILLCELL_X32 FILLER_264_1752 ();
 FILLCELL_X32 FILLER_264_1784 ();
 FILLCELL_X32 FILLER_264_1816 ();
 FILLCELL_X32 FILLER_264_1848 ();
 FILLCELL_X8 FILLER_264_1880 ();
 FILLCELL_X4 FILLER_264_1888 ();
 FILLCELL_X2 FILLER_264_1892 ();
 FILLCELL_X32 FILLER_264_1895 ();
 FILLCELL_X32 FILLER_264_1927 ();
 FILLCELL_X32 FILLER_264_1959 ();
 FILLCELL_X32 FILLER_264_1991 ();
 FILLCELL_X32 FILLER_264_2023 ();
 FILLCELL_X32 FILLER_264_2055 ();
 FILLCELL_X16 FILLER_264_2087 ();
 FILLCELL_X8 FILLER_264_2103 ();
 FILLCELL_X4 FILLER_264_2111 ();
 FILLCELL_X32 FILLER_265_1 ();
 FILLCELL_X32 FILLER_265_33 ();
 FILLCELL_X32 FILLER_265_65 ();
 FILLCELL_X32 FILLER_265_97 ();
 FILLCELL_X32 FILLER_265_129 ();
 FILLCELL_X32 FILLER_265_161 ();
 FILLCELL_X32 FILLER_265_193 ();
 FILLCELL_X32 FILLER_265_225 ();
 FILLCELL_X32 FILLER_265_257 ();
 FILLCELL_X32 FILLER_265_289 ();
 FILLCELL_X32 FILLER_265_321 ();
 FILLCELL_X32 FILLER_265_353 ();
 FILLCELL_X32 FILLER_265_385 ();
 FILLCELL_X32 FILLER_265_417 ();
 FILLCELL_X32 FILLER_265_449 ();
 FILLCELL_X32 FILLER_265_481 ();
 FILLCELL_X32 FILLER_265_513 ();
 FILLCELL_X32 FILLER_265_545 ();
 FILLCELL_X32 FILLER_265_577 ();
 FILLCELL_X32 FILLER_265_609 ();
 FILLCELL_X32 FILLER_265_641 ();
 FILLCELL_X32 FILLER_265_673 ();
 FILLCELL_X32 FILLER_265_705 ();
 FILLCELL_X32 FILLER_265_737 ();
 FILLCELL_X32 FILLER_265_769 ();
 FILLCELL_X32 FILLER_265_801 ();
 FILLCELL_X32 FILLER_265_833 ();
 FILLCELL_X32 FILLER_265_865 ();
 FILLCELL_X32 FILLER_265_897 ();
 FILLCELL_X32 FILLER_265_929 ();
 FILLCELL_X32 FILLER_265_961 ();
 FILLCELL_X32 FILLER_265_993 ();
 FILLCELL_X32 FILLER_265_1025 ();
 FILLCELL_X32 FILLER_265_1057 ();
 FILLCELL_X32 FILLER_265_1089 ();
 FILLCELL_X32 FILLER_265_1121 ();
 FILLCELL_X32 FILLER_265_1153 ();
 FILLCELL_X32 FILLER_265_1185 ();
 FILLCELL_X32 FILLER_265_1217 ();
 FILLCELL_X8 FILLER_265_1249 ();
 FILLCELL_X4 FILLER_265_1257 ();
 FILLCELL_X2 FILLER_265_1261 ();
 FILLCELL_X32 FILLER_265_1264 ();
 FILLCELL_X32 FILLER_265_1296 ();
 FILLCELL_X32 FILLER_265_1328 ();
 FILLCELL_X32 FILLER_265_1360 ();
 FILLCELL_X32 FILLER_265_1392 ();
 FILLCELL_X32 FILLER_265_1424 ();
 FILLCELL_X32 FILLER_265_1456 ();
 FILLCELL_X32 FILLER_265_1488 ();
 FILLCELL_X32 FILLER_265_1520 ();
 FILLCELL_X32 FILLER_265_1552 ();
 FILLCELL_X32 FILLER_265_1584 ();
 FILLCELL_X32 FILLER_265_1616 ();
 FILLCELL_X32 FILLER_265_1648 ();
 FILLCELL_X32 FILLER_265_1680 ();
 FILLCELL_X32 FILLER_265_1712 ();
 FILLCELL_X32 FILLER_265_1744 ();
 FILLCELL_X32 FILLER_265_1776 ();
 FILLCELL_X32 FILLER_265_1808 ();
 FILLCELL_X32 FILLER_265_1840 ();
 FILLCELL_X32 FILLER_265_1872 ();
 FILLCELL_X32 FILLER_265_1904 ();
 FILLCELL_X32 FILLER_265_1936 ();
 FILLCELL_X32 FILLER_265_1968 ();
 FILLCELL_X32 FILLER_265_2000 ();
 FILLCELL_X32 FILLER_265_2032 ();
 FILLCELL_X32 FILLER_265_2064 ();
 FILLCELL_X16 FILLER_265_2096 ();
 FILLCELL_X2 FILLER_265_2112 ();
 FILLCELL_X1 FILLER_265_2114 ();
 FILLCELL_X32 FILLER_266_1 ();
 FILLCELL_X32 FILLER_266_33 ();
 FILLCELL_X32 FILLER_266_65 ();
 FILLCELL_X32 FILLER_266_97 ();
 FILLCELL_X32 FILLER_266_129 ();
 FILLCELL_X32 FILLER_266_161 ();
 FILLCELL_X32 FILLER_266_193 ();
 FILLCELL_X32 FILLER_266_225 ();
 FILLCELL_X32 FILLER_266_257 ();
 FILLCELL_X32 FILLER_266_289 ();
 FILLCELL_X32 FILLER_266_321 ();
 FILLCELL_X32 FILLER_266_353 ();
 FILLCELL_X32 FILLER_266_385 ();
 FILLCELL_X32 FILLER_266_417 ();
 FILLCELL_X32 FILLER_266_449 ();
 FILLCELL_X32 FILLER_266_481 ();
 FILLCELL_X32 FILLER_266_513 ();
 FILLCELL_X32 FILLER_266_545 ();
 FILLCELL_X32 FILLER_266_577 ();
 FILLCELL_X16 FILLER_266_609 ();
 FILLCELL_X4 FILLER_266_625 ();
 FILLCELL_X2 FILLER_266_629 ();
 FILLCELL_X32 FILLER_266_632 ();
 FILLCELL_X32 FILLER_266_664 ();
 FILLCELL_X32 FILLER_266_696 ();
 FILLCELL_X32 FILLER_266_728 ();
 FILLCELL_X32 FILLER_266_760 ();
 FILLCELL_X32 FILLER_266_792 ();
 FILLCELL_X32 FILLER_266_824 ();
 FILLCELL_X32 FILLER_266_856 ();
 FILLCELL_X32 FILLER_266_888 ();
 FILLCELL_X32 FILLER_266_920 ();
 FILLCELL_X32 FILLER_266_952 ();
 FILLCELL_X32 FILLER_266_984 ();
 FILLCELL_X32 FILLER_266_1016 ();
 FILLCELL_X32 FILLER_266_1048 ();
 FILLCELL_X32 FILLER_266_1080 ();
 FILLCELL_X32 FILLER_266_1112 ();
 FILLCELL_X32 FILLER_266_1144 ();
 FILLCELL_X32 FILLER_266_1176 ();
 FILLCELL_X32 FILLER_266_1208 ();
 FILLCELL_X32 FILLER_266_1240 ();
 FILLCELL_X32 FILLER_266_1272 ();
 FILLCELL_X32 FILLER_266_1304 ();
 FILLCELL_X32 FILLER_266_1336 ();
 FILLCELL_X32 FILLER_266_1368 ();
 FILLCELL_X32 FILLER_266_1400 ();
 FILLCELL_X32 FILLER_266_1432 ();
 FILLCELL_X32 FILLER_266_1464 ();
 FILLCELL_X32 FILLER_266_1496 ();
 FILLCELL_X32 FILLER_266_1528 ();
 FILLCELL_X32 FILLER_266_1560 ();
 FILLCELL_X32 FILLER_266_1592 ();
 FILLCELL_X32 FILLER_266_1624 ();
 FILLCELL_X32 FILLER_266_1656 ();
 FILLCELL_X32 FILLER_266_1688 ();
 FILLCELL_X32 FILLER_266_1720 ();
 FILLCELL_X32 FILLER_266_1752 ();
 FILLCELL_X32 FILLER_266_1784 ();
 FILLCELL_X32 FILLER_266_1816 ();
 FILLCELL_X32 FILLER_266_1848 ();
 FILLCELL_X8 FILLER_266_1880 ();
 FILLCELL_X4 FILLER_266_1888 ();
 FILLCELL_X2 FILLER_266_1892 ();
 FILLCELL_X32 FILLER_266_1895 ();
 FILLCELL_X32 FILLER_266_1927 ();
 FILLCELL_X32 FILLER_266_1959 ();
 FILLCELL_X32 FILLER_266_1991 ();
 FILLCELL_X32 FILLER_266_2023 ();
 FILLCELL_X32 FILLER_266_2055 ();
 FILLCELL_X16 FILLER_266_2087 ();
 FILLCELL_X8 FILLER_266_2103 ();
 FILLCELL_X4 FILLER_266_2111 ();
 FILLCELL_X32 FILLER_267_1 ();
 FILLCELL_X32 FILLER_267_33 ();
 FILLCELL_X32 FILLER_267_65 ();
 FILLCELL_X32 FILLER_267_97 ();
 FILLCELL_X32 FILLER_267_129 ();
 FILLCELL_X32 FILLER_267_161 ();
 FILLCELL_X32 FILLER_267_193 ();
 FILLCELL_X32 FILLER_267_225 ();
 FILLCELL_X32 FILLER_267_257 ();
 FILLCELL_X32 FILLER_267_289 ();
 FILLCELL_X32 FILLER_267_321 ();
 FILLCELL_X32 FILLER_267_353 ();
 FILLCELL_X32 FILLER_267_385 ();
 FILLCELL_X32 FILLER_267_417 ();
 FILLCELL_X32 FILLER_267_449 ();
 FILLCELL_X32 FILLER_267_481 ();
 FILLCELL_X32 FILLER_267_513 ();
 FILLCELL_X32 FILLER_267_545 ();
 FILLCELL_X32 FILLER_267_577 ();
 FILLCELL_X32 FILLER_267_609 ();
 FILLCELL_X32 FILLER_267_641 ();
 FILLCELL_X32 FILLER_267_673 ();
 FILLCELL_X32 FILLER_267_705 ();
 FILLCELL_X32 FILLER_267_737 ();
 FILLCELL_X32 FILLER_267_769 ();
 FILLCELL_X32 FILLER_267_801 ();
 FILLCELL_X32 FILLER_267_833 ();
 FILLCELL_X32 FILLER_267_865 ();
 FILLCELL_X32 FILLER_267_897 ();
 FILLCELL_X32 FILLER_267_929 ();
 FILLCELL_X32 FILLER_267_961 ();
 FILLCELL_X32 FILLER_267_993 ();
 FILLCELL_X32 FILLER_267_1025 ();
 FILLCELL_X32 FILLER_267_1057 ();
 FILLCELL_X32 FILLER_267_1089 ();
 FILLCELL_X32 FILLER_267_1121 ();
 FILLCELL_X32 FILLER_267_1153 ();
 FILLCELL_X32 FILLER_267_1185 ();
 FILLCELL_X32 FILLER_267_1217 ();
 FILLCELL_X8 FILLER_267_1249 ();
 FILLCELL_X4 FILLER_267_1257 ();
 FILLCELL_X2 FILLER_267_1261 ();
 FILLCELL_X32 FILLER_267_1264 ();
 FILLCELL_X32 FILLER_267_1296 ();
 FILLCELL_X32 FILLER_267_1328 ();
 FILLCELL_X32 FILLER_267_1360 ();
 FILLCELL_X32 FILLER_267_1392 ();
 FILLCELL_X32 FILLER_267_1424 ();
 FILLCELL_X32 FILLER_267_1456 ();
 FILLCELL_X32 FILLER_267_1488 ();
 FILLCELL_X32 FILLER_267_1520 ();
 FILLCELL_X32 FILLER_267_1552 ();
 FILLCELL_X32 FILLER_267_1584 ();
 FILLCELL_X32 FILLER_267_1616 ();
 FILLCELL_X32 FILLER_267_1648 ();
 FILLCELL_X32 FILLER_267_1680 ();
 FILLCELL_X32 FILLER_267_1712 ();
 FILLCELL_X32 FILLER_267_1744 ();
 FILLCELL_X32 FILLER_267_1776 ();
 FILLCELL_X32 FILLER_267_1808 ();
 FILLCELL_X32 FILLER_267_1840 ();
 FILLCELL_X32 FILLER_267_1872 ();
 FILLCELL_X32 FILLER_267_1904 ();
 FILLCELL_X32 FILLER_267_1936 ();
 FILLCELL_X32 FILLER_267_1968 ();
 FILLCELL_X32 FILLER_267_2000 ();
 FILLCELL_X32 FILLER_267_2032 ();
 FILLCELL_X32 FILLER_267_2064 ();
 FILLCELL_X16 FILLER_267_2096 ();
 FILLCELL_X2 FILLER_267_2112 ();
 FILLCELL_X1 FILLER_267_2114 ();
 FILLCELL_X32 FILLER_268_1 ();
 FILLCELL_X32 FILLER_268_33 ();
 FILLCELL_X32 FILLER_268_65 ();
 FILLCELL_X32 FILLER_268_97 ();
 FILLCELL_X32 FILLER_268_129 ();
 FILLCELL_X32 FILLER_268_161 ();
 FILLCELL_X32 FILLER_268_193 ();
 FILLCELL_X32 FILLER_268_225 ();
 FILLCELL_X32 FILLER_268_257 ();
 FILLCELL_X32 FILLER_268_289 ();
 FILLCELL_X32 FILLER_268_321 ();
 FILLCELL_X32 FILLER_268_353 ();
 FILLCELL_X32 FILLER_268_385 ();
 FILLCELL_X32 FILLER_268_417 ();
 FILLCELL_X32 FILLER_268_449 ();
 FILLCELL_X32 FILLER_268_481 ();
 FILLCELL_X32 FILLER_268_513 ();
 FILLCELL_X32 FILLER_268_545 ();
 FILLCELL_X32 FILLER_268_577 ();
 FILLCELL_X16 FILLER_268_609 ();
 FILLCELL_X4 FILLER_268_625 ();
 FILLCELL_X2 FILLER_268_629 ();
 FILLCELL_X32 FILLER_268_632 ();
 FILLCELL_X32 FILLER_268_664 ();
 FILLCELL_X32 FILLER_268_696 ();
 FILLCELL_X32 FILLER_268_728 ();
 FILLCELL_X32 FILLER_268_760 ();
 FILLCELL_X32 FILLER_268_792 ();
 FILLCELL_X32 FILLER_268_824 ();
 FILLCELL_X32 FILLER_268_856 ();
 FILLCELL_X32 FILLER_268_888 ();
 FILLCELL_X32 FILLER_268_920 ();
 FILLCELL_X32 FILLER_268_952 ();
 FILLCELL_X32 FILLER_268_984 ();
 FILLCELL_X32 FILLER_268_1016 ();
 FILLCELL_X32 FILLER_268_1048 ();
 FILLCELL_X32 FILLER_268_1080 ();
 FILLCELL_X32 FILLER_268_1112 ();
 FILLCELL_X32 FILLER_268_1144 ();
 FILLCELL_X32 FILLER_268_1176 ();
 FILLCELL_X32 FILLER_268_1208 ();
 FILLCELL_X32 FILLER_268_1240 ();
 FILLCELL_X32 FILLER_268_1272 ();
 FILLCELL_X32 FILLER_268_1304 ();
 FILLCELL_X32 FILLER_268_1336 ();
 FILLCELL_X32 FILLER_268_1368 ();
 FILLCELL_X32 FILLER_268_1400 ();
 FILLCELL_X32 FILLER_268_1432 ();
 FILLCELL_X32 FILLER_268_1464 ();
 FILLCELL_X32 FILLER_268_1496 ();
 FILLCELL_X32 FILLER_268_1528 ();
 FILLCELL_X32 FILLER_268_1560 ();
 FILLCELL_X32 FILLER_268_1592 ();
 FILLCELL_X32 FILLER_268_1624 ();
 FILLCELL_X32 FILLER_268_1656 ();
 FILLCELL_X32 FILLER_268_1688 ();
 FILLCELL_X32 FILLER_268_1720 ();
 FILLCELL_X32 FILLER_268_1752 ();
 FILLCELL_X32 FILLER_268_1784 ();
 FILLCELL_X32 FILLER_268_1816 ();
 FILLCELL_X32 FILLER_268_1848 ();
 FILLCELL_X8 FILLER_268_1880 ();
 FILLCELL_X4 FILLER_268_1888 ();
 FILLCELL_X2 FILLER_268_1892 ();
 FILLCELL_X32 FILLER_268_1895 ();
 FILLCELL_X32 FILLER_268_1927 ();
 FILLCELL_X32 FILLER_268_1959 ();
 FILLCELL_X32 FILLER_268_1991 ();
 FILLCELL_X32 FILLER_268_2023 ();
 FILLCELL_X32 FILLER_268_2055 ();
 FILLCELL_X16 FILLER_268_2087 ();
 FILLCELL_X8 FILLER_268_2103 ();
 FILLCELL_X4 FILLER_268_2111 ();
 FILLCELL_X32 FILLER_269_1 ();
 FILLCELL_X32 FILLER_269_33 ();
 FILLCELL_X32 FILLER_269_65 ();
 FILLCELL_X32 FILLER_269_97 ();
 FILLCELL_X32 FILLER_269_129 ();
 FILLCELL_X32 FILLER_269_161 ();
 FILLCELL_X32 FILLER_269_193 ();
 FILLCELL_X32 FILLER_269_225 ();
 FILLCELL_X32 FILLER_269_257 ();
 FILLCELL_X32 FILLER_269_289 ();
 FILLCELL_X32 FILLER_269_321 ();
 FILLCELL_X32 FILLER_269_353 ();
 FILLCELL_X32 FILLER_269_385 ();
 FILLCELL_X32 FILLER_269_417 ();
 FILLCELL_X32 FILLER_269_449 ();
 FILLCELL_X32 FILLER_269_481 ();
 FILLCELL_X32 FILLER_269_513 ();
 FILLCELL_X32 FILLER_269_545 ();
 FILLCELL_X32 FILLER_269_577 ();
 FILLCELL_X32 FILLER_269_609 ();
 FILLCELL_X32 FILLER_269_641 ();
 FILLCELL_X32 FILLER_269_673 ();
 FILLCELL_X32 FILLER_269_705 ();
 FILLCELL_X32 FILLER_269_737 ();
 FILLCELL_X32 FILLER_269_769 ();
 FILLCELL_X32 FILLER_269_801 ();
 FILLCELL_X32 FILLER_269_833 ();
 FILLCELL_X32 FILLER_269_865 ();
 FILLCELL_X32 FILLER_269_897 ();
 FILLCELL_X32 FILLER_269_929 ();
 FILLCELL_X32 FILLER_269_961 ();
 FILLCELL_X32 FILLER_269_993 ();
 FILLCELL_X32 FILLER_269_1025 ();
 FILLCELL_X32 FILLER_269_1057 ();
 FILLCELL_X32 FILLER_269_1089 ();
 FILLCELL_X32 FILLER_269_1121 ();
 FILLCELL_X32 FILLER_269_1153 ();
 FILLCELL_X32 FILLER_269_1185 ();
 FILLCELL_X32 FILLER_269_1217 ();
 FILLCELL_X8 FILLER_269_1249 ();
 FILLCELL_X4 FILLER_269_1257 ();
 FILLCELL_X2 FILLER_269_1261 ();
 FILLCELL_X32 FILLER_269_1264 ();
 FILLCELL_X32 FILLER_269_1296 ();
 FILLCELL_X32 FILLER_269_1328 ();
 FILLCELL_X32 FILLER_269_1360 ();
 FILLCELL_X32 FILLER_269_1392 ();
 FILLCELL_X32 FILLER_269_1424 ();
 FILLCELL_X32 FILLER_269_1456 ();
 FILLCELL_X32 FILLER_269_1488 ();
 FILLCELL_X32 FILLER_269_1520 ();
 FILLCELL_X32 FILLER_269_1552 ();
 FILLCELL_X32 FILLER_269_1584 ();
 FILLCELL_X32 FILLER_269_1616 ();
 FILLCELL_X32 FILLER_269_1648 ();
 FILLCELL_X32 FILLER_269_1680 ();
 FILLCELL_X32 FILLER_269_1712 ();
 FILLCELL_X32 FILLER_269_1744 ();
 FILLCELL_X32 FILLER_269_1776 ();
 FILLCELL_X32 FILLER_269_1808 ();
 FILLCELL_X32 FILLER_269_1840 ();
 FILLCELL_X32 FILLER_269_1872 ();
 FILLCELL_X32 FILLER_269_1904 ();
 FILLCELL_X32 FILLER_269_1936 ();
 FILLCELL_X32 FILLER_269_1968 ();
 FILLCELL_X32 FILLER_269_2000 ();
 FILLCELL_X32 FILLER_269_2032 ();
 FILLCELL_X32 FILLER_269_2064 ();
 FILLCELL_X16 FILLER_269_2096 ();
 FILLCELL_X2 FILLER_269_2112 ();
 FILLCELL_X1 FILLER_269_2114 ();
 FILLCELL_X32 FILLER_270_1 ();
 FILLCELL_X32 FILLER_270_33 ();
 FILLCELL_X32 FILLER_270_65 ();
 FILLCELL_X32 FILLER_270_97 ();
 FILLCELL_X32 FILLER_270_129 ();
 FILLCELL_X32 FILLER_270_161 ();
 FILLCELL_X32 FILLER_270_193 ();
 FILLCELL_X32 FILLER_270_225 ();
 FILLCELL_X32 FILLER_270_257 ();
 FILLCELL_X32 FILLER_270_289 ();
 FILLCELL_X32 FILLER_270_321 ();
 FILLCELL_X32 FILLER_270_353 ();
 FILLCELL_X32 FILLER_270_385 ();
 FILLCELL_X32 FILLER_270_417 ();
 FILLCELL_X32 FILLER_270_449 ();
 FILLCELL_X32 FILLER_270_481 ();
 FILLCELL_X32 FILLER_270_513 ();
 FILLCELL_X32 FILLER_270_545 ();
 FILLCELL_X32 FILLER_270_577 ();
 FILLCELL_X16 FILLER_270_609 ();
 FILLCELL_X4 FILLER_270_625 ();
 FILLCELL_X2 FILLER_270_629 ();
 FILLCELL_X32 FILLER_270_632 ();
 FILLCELL_X32 FILLER_270_664 ();
 FILLCELL_X32 FILLER_270_696 ();
 FILLCELL_X32 FILLER_270_728 ();
 FILLCELL_X32 FILLER_270_760 ();
 FILLCELL_X32 FILLER_270_792 ();
 FILLCELL_X32 FILLER_270_824 ();
 FILLCELL_X32 FILLER_270_856 ();
 FILLCELL_X32 FILLER_270_888 ();
 FILLCELL_X32 FILLER_270_920 ();
 FILLCELL_X32 FILLER_270_952 ();
 FILLCELL_X32 FILLER_270_984 ();
 FILLCELL_X32 FILLER_270_1016 ();
 FILLCELL_X32 FILLER_270_1048 ();
 FILLCELL_X32 FILLER_270_1080 ();
 FILLCELL_X32 FILLER_270_1112 ();
 FILLCELL_X32 FILLER_270_1144 ();
 FILLCELL_X32 FILLER_270_1176 ();
 FILLCELL_X32 FILLER_270_1208 ();
 FILLCELL_X32 FILLER_270_1240 ();
 FILLCELL_X32 FILLER_270_1272 ();
 FILLCELL_X32 FILLER_270_1304 ();
 FILLCELL_X32 FILLER_270_1336 ();
 FILLCELL_X32 FILLER_270_1368 ();
 FILLCELL_X32 FILLER_270_1400 ();
 FILLCELL_X32 FILLER_270_1432 ();
 FILLCELL_X32 FILLER_270_1464 ();
 FILLCELL_X32 FILLER_270_1496 ();
 FILLCELL_X32 FILLER_270_1528 ();
 FILLCELL_X32 FILLER_270_1560 ();
 FILLCELL_X32 FILLER_270_1592 ();
 FILLCELL_X32 FILLER_270_1624 ();
 FILLCELL_X32 FILLER_270_1656 ();
 FILLCELL_X32 FILLER_270_1688 ();
 FILLCELL_X32 FILLER_270_1720 ();
 FILLCELL_X32 FILLER_270_1752 ();
 FILLCELL_X32 FILLER_270_1784 ();
 FILLCELL_X32 FILLER_270_1816 ();
 FILLCELL_X32 FILLER_270_1848 ();
 FILLCELL_X8 FILLER_270_1880 ();
 FILLCELL_X4 FILLER_270_1888 ();
 FILLCELL_X2 FILLER_270_1892 ();
 FILLCELL_X32 FILLER_270_1895 ();
 FILLCELL_X32 FILLER_270_1927 ();
 FILLCELL_X32 FILLER_270_1959 ();
 FILLCELL_X32 FILLER_270_1991 ();
 FILLCELL_X32 FILLER_270_2023 ();
 FILLCELL_X32 FILLER_270_2055 ();
 FILLCELL_X16 FILLER_270_2087 ();
 FILLCELL_X8 FILLER_270_2103 ();
 FILLCELL_X4 FILLER_270_2111 ();
 FILLCELL_X32 FILLER_271_1 ();
 FILLCELL_X32 FILLER_271_33 ();
 FILLCELL_X32 FILLER_271_65 ();
 FILLCELL_X32 FILLER_271_97 ();
 FILLCELL_X32 FILLER_271_129 ();
 FILLCELL_X32 FILLER_271_161 ();
 FILLCELL_X32 FILLER_271_193 ();
 FILLCELL_X32 FILLER_271_225 ();
 FILLCELL_X32 FILLER_271_257 ();
 FILLCELL_X32 FILLER_271_289 ();
 FILLCELL_X32 FILLER_271_321 ();
 FILLCELL_X32 FILLER_271_353 ();
 FILLCELL_X32 FILLER_271_385 ();
 FILLCELL_X32 FILLER_271_417 ();
 FILLCELL_X32 FILLER_271_449 ();
 FILLCELL_X32 FILLER_271_481 ();
 FILLCELL_X32 FILLER_271_513 ();
 FILLCELL_X32 FILLER_271_545 ();
 FILLCELL_X32 FILLER_271_577 ();
 FILLCELL_X32 FILLER_271_609 ();
 FILLCELL_X32 FILLER_271_641 ();
 FILLCELL_X32 FILLER_271_673 ();
 FILLCELL_X32 FILLER_271_705 ();
 FILLCELL_X32 FILLER_271_737 ();
 FILLCELL_X32 FILLER_271_769 ();
 FILLCELL_X32 FILLER_271_801 ();
 FILLCELL_X32 FILLER_271_833 ();
 FILLCELL_X32 FILLER_271_865 ();
 FILLCELL_X32 FILLER_271_897 ();
 FILLCELL_X32 FILLER_271_929 ();
 FILLCELL_X32 FILLER_271_961 ();
 FILLCELL_X32 FILLER_271_993 ();
 FILLCELL_X32 FILLER_271_1025 ();
 FILLCELL_X32 FILLER_271_1057 ();
 FILLCELL_X32 FILLER_271_1089 ();
 FILLCELL_X32 FILLER_271_1121 ();
 FILLCELL_X32 FILLER_271_1153 ();
 FILLCELL_X32 FILLER_271_1185 ();
 FILLCELL_X32 FILLER_271_1217 ();
 FILLCELL_X8 FILLER_271_1249 ();
 FILLCELL_X4 FILLER_271_1257 ();
 FILLCELL_X2 FILLER_271_1261 ();
 FILLCELL_X32 FILLER_271_1264 ();
 FILLCELL_X32 FILLER_271_1296 ();
 FILLCELL_X32 FILLER_271_1328 ();
 FILLCELL_X32 FILLER_271_1360 ();
 FILLCELL_X32 FILLER_271_1392 ();
 FILLCELL_X32 FILLER_271_1424 ();
 FILLCELL_X32 FILLER_271_1456 ();
 FILLCELL_X32 FILLER_271_1488 ();
 FILLCELL_X32 FILLER_271_1520 ();
 FILLCELL_X32 FILLER_271_1552 ();
 FILLCELL_X32 FILLER_271_1584 ();
 FILLCELL_X32 FILLER_271_1616 ();
 FILLCELL_X32 FILLER_271_1648 ();
 FILLCELL_X32 FILLER_271_1680 ();
 FILLCELL_X32 FILLER_271_1712 ();
 FILLCELL_X32 FILLER_271_1744 ();
 FILLCELL_X32 FILLER_271_1776 ();
 FILLCELL_X32 FILLER_271_1808 ();
 FILLCELL_X32 FILLER_271_1840 ();
 FILLCELL_X32 FILLER_271_1872 ();
 FILLCELL_X32 FILLER_271_1904 ();
 FILLCELL_X32 FILLER_271_1936 ();
 FILLCELL_X32 FILLER_271_1968 ();
 FILLCELL_X32 FILLER_271_2000 ();
 FILLCELL_X32 FILLER_271_2032 ();
 FILLCELL_X32 FILLER_271_2064 ();
 FILLCELL_X16 FILLER_271_2096 ();
 FILLCELL_X2 FILLER_271_2112 ();
 FILLCELL_X1 FILLER_271_2114 ();
 FILLCELL_X32 FILLER_272_1 ();
 FILLCELL_X32 FILLER_272_33 ();
 FILLCELL_X32 FILLER_272_65 ();
 FILLCELL_X32 FILLER_272_97 ();
 FILLCELL_X32 FILLER_272_129 ();
 FILLCELL_X32 FILLER_272_161 ();
 FILLCELL_X32 FILLER_272_193 ();
 FILLCELL_X32 FILLER_272_225 ();
 FILLCELL_X32 FILLER_272_257 ();
 FILLCELL_X32 FILLER_272_289 ();
 FILLCELL_X32 FILLER_272_321 ();
 FILLCELL_X32 FILLER_272_353 ();
 FILLCELL_X32 FILLER_272_385 ();
 FILLCELL_X32 FILLER_272_417 ();
 FILLCELL_X32 FILLER_272_449 ();
 FILLCELL_X32 FILLER_272_481 ();
 FILLCELL_X32 FILLER_272_513 ();
 FILLCELL_X32 FILLER_272_545 ();
 FILLCELL_X32 FILLER_272_577 ();
 FILLCELL_X16 FILLER_272_609 ();
 FILLCELL_X4 FILLER_272_625 ();
 FILLCELL_X2 FILLER_272_629 ();
 FILLCELL_X32 FILLER_272_632 ();
 FILLCELL_X32 FILLER_272_664 ();
 FILLCELL_X32 FILLER_272_696 ();
 FILLCELL_X32 FILLER_272_728 ();
 FILLCELL_X32 FILLER_272_760 ();
 FILLCELL_X32 FILLER_272_792 ();
 FILLCELL_X32 FILLER_272_824 ();
 FILLCELL_X32 FILLER_272_856 ();
 FILLCELL_X32 FILLER_272_888 ();
 FILLCELL_X32 FILLER_272_920 ();
 FILLCELL_X32 FILLER_272_952 ();
 FILLCELL_X32 FILLER_272_984 ();
 FILLCELL_X32 FILLER_272_1016 ();
 FILLCELL_X32 FILLER_272_1048 ();
 FILLCELL_X32 FILLER_272_1080 ();
 FILLCELL_X32 FILLER_272_1112 ();
 FILLCELL_X32 FILLER_272_1144 ();
 FILLCELL_X32 FILLER_272_1176 ();
 FILLCELL_X32 FILLER_272_1208 ();
 FILLCELL_X32 FILLER_272_1240 ();
 FILLCELL_X32 FILLER_272_1272 ();
 FILLCELL_X32 FILLER_272_1304 ();
 FILLCELL_X32 FILLER_272_1336 ();
 FILLCELL_X32 FILLER_272_1368 ();
 FILLCELL_X32 FILLER_272_1400 ();
 FILLCELL_X32 FILLER_272_1432 ();
 FILLCELL_X32 FILLER_272_1464 ();
 FILLCELL_X32 FILLER_272_1496 ();
 FILLCELL_X32 FILLER_272_1528 ();
 FILLCELL_X32 FILLER_272_1560 ();
 FILLCELL_X32 FILLER_272_1592 ();
 FILLCELL_X32 FILLER_272_1624 ();
 FILLCELL_X32 FILLER_272_1656 ();
 FILLCELL_X32 FILLER_272_1688 ();
 FILLCELL_X32 FILLER_272_1720 ();
 FILLCELL_X32 FILLER_272_1752 ();
 FILLCELL_X32 FILLER_272_1784 ();
 FILLCELL_X32 FILLER_272_1816 ();
 FILLCELL_X32 FILLER_272_1848 ();
 FILLCELL_X8 FILLER_272_1880 ();
 FILLCELL_X4 FILLER_272_1888 ();
 FILLCELL_X2 FILLER_272_1892 ();
 FILLCELL_X32 FILLER_272_1895 ();
 FILLCELL_X32 FILLER_272_1927 ();
 FILLCELL_X32 FILLER_272_1959 ();
 FILLCELL_X32 FILLER_272_1991 ();
 FILLCELL_X32 FILLER_272_2023 ();
 FILLCELL_X32 FILLER_272_2055 ();
 FILLCELL_X16 FILLER_272_2087 ();
 FILLCELL_X8 FILLER_272_2103 ();
 FILLCELL_X4 FILLER_272_2111 ();
 FILLCELL_X32 FILLER_273_1 ();
 FILLCELL_X32 FILLER_273_33 ();
 FILLCELL_X32 FILLER_273_65 ();
 FILLCELL_X32 FILLER_273_97 ();
 FILLCELL_X32 FILLER_273_129 ();
 FILLCELL_X32 FILLER_273_161 ();
 FILLCELL_X32 FILLER_273_193 ();
 FILLCELL_X32 FILLER_273_225 ();
 FILLCELL_X32 FILLER_273_257 ();
 FILLCELL_X32 FILLER_273_289 ();
 FILLCELL_X32 FILLER_273_321 ();
 FILLCELL_X32 FILLER_273_353 ();
 FILLCELL_X32 FILLER_273_385 ();
 FILLCELL_X32 FILLER_273_417 ();
 FILLCELL_X32 FILLER_273_449 ();
 FILLCELL_X32 FILLER_273_481 ();
 FILLCELL_X32 FILLER_273_513 ();
 FILLCELL_X32 FILLER_273_545 ();
 FILLCELL_X32 FILLER_273_577 ();
 FILLCELL_X32 FILLER_273_609 ();
 FILLCELL_X32 FILLER_273_641 ();
 FILLCELL_X32 FILLER_273_673 ();
 FILLCELL_X32 FILLER_273_705 ();
 FILLCELL_X32 FILLER_273_737 ();
 FILLCELL_X32 FILLER_273_769 ();
 FILLCELL_X32 FILLER_273_801 ();
 FILLCELL_X32 FILLER_273_833 ();
 FILLCELL_X32 FILLER_273_865 ();
 FILLCELL_X32 FILLER_273_897 ();
 FILLCELL_X32 FILLER_273_929 ();
 FILLCELL_X32 FILLER_273_961 ();
 FILLCELL_X32 FILLER_273_993 ();
 FILLCELL_X32 FILLER_273_1025 ();
 FILLCELL_X32 FILLER_273_1057 ();
 FILLCELL_X32 FILLER_273_1089 ();
 FILLCELL_X32 FILLER_273_1121 ();
 FILLCELL_X32 FILLER_273_1153 ();
 FILLCELL_X32 FILLER_273_1185 ();
 FILLCELL_X32 FILLER_273_1217 ();
 FILLCELL_X8 FILLER_273_1249 ();
 FILLCELL_X4 FILLER_273_1257 ();
 FILLCELL_X2 FILLER_273_1261 ();
 FILLCELL_X32 FILLER_273_1264 ();
 FILLCELL_X32 FILLER_273_1296 ();
 FILLCELL_X32 FILLER_273_1328 ();
 FILLCELL_X32 FILLER_273_1360 ();
 FILLCELL_X32 FILLER_273_1392 ();
 FILLCELL_X32 FILLER_273_1424 ();
 FILLCELL_X32 FILLER_273_1456 ();
 FILLCELL_X32 FILLER_273_1488 ();
 FILLCELL_X32 FILLER_273_1520 ();
 FILLCELL_X32 FILLER_273_1552 ();
 FILLCELL_X32 FILLER_273_1584 ();
 FILLCELL_X32 FILLER_273_1616 ();
 FILLCELL_X32 FILLER_273_1648 ();
 FILLCELL_X32 FILLER_273_1680 ();
 FILLCELL_X32 FILLER_273_1712 ();
 FILLCELL_X32 FILLER_273_1744 ();
 FILLCELL_X32 FILLER_273_1776 ();
 FILLCELL_X32 FILLER_273_1808 ();
 FILLCELL_X32 FILLER_273_1840 ();
 FILLCELL_X32 FILLER_273_1872 ();
 FILLCELL_X32 FILLER_273_1904 ();
 FILLCELL_X32 FILLER_273_1936 ();
 FILLCELL_X32 FILLER_273_1968 ();
 FILLCELL_X32 FILLER_273_2000 ();
 FILLCELL_X32 FILLER_273_2032 ();
 FILLCELL_X32 FILLER_273_2064 ();
 FILLCELL_X16 FILLER_273_2096 ();
 FILLCELL_X2 FILLER_273_2112 ();
 FILLCELL_X1 FILLER_273_2114 ();
 FILLCELL_X32 FILLER_274_1 ();
 FILLCELL_X32 FILLER_274_33 ();
 FILLCELL_X32 FILLER_274_65 ();
 FILLCELL_X32 FILLER_274_97 ();
 FILLCELL_X32 FILLER_274_129 ();
 FILLCELL_X32 FILLER_274_161 ();
 FILLCELL_X32 FILLER_274_193 ();
 FILLCELL_X32 FILLER_274_225 ();
 FILLCELL_X32 FILLER_274_257 ();
 FILLCELL_X32 FILLER_274_289 ();
 FILLCELL_X32 FILLER_274_321 ();
 FILLCELL_X32 FILLER_274_353 ();
 FILLCELL_X32 FILLER_274_385 ();
 FILLCELL_X32 FILLER_274_417 ();
 FILLCELL_X32 FILLER_274_449 ();
 FILLCELL_X32 FILLER_274_481 ();
 FILLCELL_X32 FILLER_274_513 ();
 FILLCELL_X32 FILLER_274_545 ();
 FILLCELL_X32 FILLER_274_577 ();
 FILLCELL_X16 FILLER_274_609 ();
 FILLCELL_X4 FILLER_274_625 ();
 FILLCELL_X2 FILLER_274_629 ();
 FILLCELL_X32 FILLER_274_632 ();
 FILLCELL_X32 FILLER_274_664 ();
 FILLCELL_X32 FILLER_274_696 ();
 FILLCELL_X32 FILLER_274_728 ();
 FILLCELL_X32 FILLER_274_760 ();
 FILLCELL_X32 FILLER_274_792 ();
 FILLCELL_X32 FILLER_274_824 ();
 FILLCELL_X32 FILLER_274_856 ();
 FILLCELL_X32 FILLER_274_888 ();
 FILLCELL_X32 FILLER_274_920 ();
 FILLCELL_X32 FILLER_274_952 ();
 FILLCELL_X32 FILLER_274_984 ();
 FILLCELL_X32 FILLER_274_1016 ();
 FILLCELL_X32 FILLER_274_1048 ();
 FILLCELL_X32 FILLER_274_1080 ();
 FILLCELL_X32 FILLER_274_1112 ();
 FILLCELL_X32 FILLER_274_1144 ();
 FILLCELL_X32 FILLER_274_1176 ();
 FILLCELL_X32 FILLER_274_1208 ();
 FILLCELL_X32 FILLER_274_1240 ();
 FILLCELL_X32 FILLER_274_1272 ();
 FILLCELL_X32 FILLER_274_1304 ();
 FILLCELL_X32 FILLER_274_1336 ();
 FILLCELL_X32 FILLER_274_1368 ();
 FILLCELL_X32 FILLER_274_1400 ();
 FILLCELL_X32 FILLER_274_1432 ();
 FILLCELL_X32 FILLER_274_1464 ();
 FILLCELL_X32 FILLER_274_1496 ();
 FILLCELL_X32 FILLER_274_1528 ();
 FILLCELL_X32 FILLER_274_1560 ();
 FILLCELL_X32 FILLER_274_1592 ();
 FILLCELL_X32 FILLER_274_1624 ();
 FILLCELL_X32 FILLER_274_1656 ();
 FILLCELL_X32 FILLER_274_1688 ();
 FILLCELL_X32 FILLER_274_1720 ();
 FILLCELL_X32 FILLER_274_1752 ();
 FILLCELL_X32 FILLER_274_1784 ();
 FILLCELL_X32 FILLER_274_1816 ();
 FILLCELL_X32 FILLER_274_1848 ();
 FILLCELL_X8 FILLER_274_1880 ();
 FILLCELL_X4 FILLER_274_1888 ();
 FILLCELL_X2 FILLER_274_1892 ();
 FILLCELL_X32 FILLER_274_1895 ();
 FILLCELL_X32 FILLER_274_1927 ();
 FILLCELL_X32 FILLER_274_1959 ();
 FILLCELL_X32 FILLER_274_1991 ();
 FILLCELL_X32 FILLER_274_2023 ();
 FILLCELL_X32 FILLER_274_2055 ();
 FILLCELL_X16 FILLER_274_2087 ();
 FILLCELL_X8 FILLER_274_2103 ();
 FILLCELL_X4 FILLER_274_2111 ();
 FILLCELL_X32 FILLER_275_1 ();
 FILLCELL_X32 FILLER_275_33 ();
 FILLCELL_X32 FILLER_275_65 ();
 FILLCELL_X32 FILLER_275_97 ();
 FILLCELL_X32 FILLER_275_129 ();
 FILLCELL_X32 FILLER_275_161 ();
 FILLCELL_X32 FILLER_275_193 ();
 FILLCELL_X32 FILLER_275_225 ();
 FILLCELL_X32 FILLER_275_257 ();
 FILLCELL_X32 FILLER_275_289 ();
 FILLCELL_X32 FILLER_275_321 ();
 FILLCELL_X32 FILLER_275_353 ();
 FILLCELL_X32 FILLER_275_385 ();
 FILLCELL_X32 FILLER_275_417 ();
 FILLCELL_X32 FILLER_275_449 ();
 FILLCELL_X32 FILLER_275_481 ();
 FILLCELL_X32 FILLER_275_513 ();
 FILLCELL_X32 FILLER_275_545 ();
 FILLCELL_X32 FILLER_275_577 ();
 FILLCELL_X32 FILLER_275_609 ();
 FILLCELL_X32 FILLER_275_641 ();
 FILLCELL_X32 FILLER_275_673 ();
 FILLCELL_X32 FILLER_275_705 ();
 FILLCELL_X32 FILLER_275_737 ();
 FILLCELL_X32 FILLER_275_769 ();
 FILLCELL_X32 FILLER_275_801 ();
 FILLCELL_X32 FILLER_275_833 ();
 FILLCELL_X32 FILLER_275_865 ();
 FILLCELL_X32 FILLER_275_897 ();
 FILLCELL_X32 FILLER_275_929 ();
 FILLCELL_X32 FILLER_275_961 ();
 FILLCELL_X32 FILLER_275_993 ();
 FILLCELL_X32 FILLER_275_1025 ();
 FILLCELL_X32 FILLER_275_1057 ();
 FILLCELL_X32 FILLER_275_1089 ();
 FILLCELL_X32 FILLER_275_1121 ();
 FILLCELL_X32 FILLER_275_1153 ();
 FILLCELL_X32 FILLER_275_1185 ();
 FILLCELL_X32 FILLER_275_1217 ();
 FILLCELL_X8 FILLER_275_1249 ();
 FILLCELL_X4 FILLER_275_1257 ();
 FILLCELL_X2 FILLER_275_1261 ();
 FILLCELL_X32 FILLER_275_1264 ();
 FILLCELL_X32 FILLER_275_1296 ();
 FILLCELL_X32 FILLER_275_1328 ();
 FILLCELL_X32 FILLER_275_1360 ();
 FILLCELL_X32 FILLER_275_1392 ();
 FILLCELL_X32 FILLER_275_1424 ();
 FILLCELL_X32 FILLER_275_1456 ();
 FILLCELL_X32 FILLER_275_1488 ();
 FILLCELL_X32 FILLER_275_1520 ();
 FILLCELL_X32 FILLER_275_1552 ();
 FILLCELL_X32 FILLER_275_1584 ();
 FILLCELL_X32 FILLER_275_1616 ();
 FILLCELL_X32 FILLER_275_1648 ();
 FILLCELL_X32 FILLER_275_1680 ();
 FILLCELL_X32 FILLER_275_1712 ();
 FILLCELL_X32 FILLER_275_1744 ();
 FILLCELL_X32 FILLER_275_1776 ();
 FILLCELL_X32 FILLER_275_1808 ();
 FILLCELL_X32 FILLER_275_1840 ();
 FILLCELL_X32 FILLER_275_1872 ();
 FILLCELL_X32 FILLER_275_1904 ();
 FILLCELL_X32 FILLER_275_1936 ();
 FILLCELL_X32 FILLER_275_1968 ();
 FILLCELL_X32 FILLER_275_2000 ();
 FILLCELL_X32 FILLER_275_2032 ();
 FILLCELL_X32 FILLER_275_2064 ();
 FILLCELL_X16 FILLER_275_2096 ();
 FILLCELL_X2 FILLER_275_2112 ();
 FILLCELL_X1 FILLER_275_2114 ();
 FILLCELL_X32 FILLER_276_1 ();
 FILLCELL_X32 FILLER_276_33 ();
 FILLCELL_X32 FILLER_276_65 ();
 FILLCELL_X32 FILLER_276_97 ();
 FILLCELL_X32 FILLER_276_129 ();
 FILLCELL_X32 FILLER_276_161 ();
 FILLCELL_X32 FILLER_276_193 ();
 FILLCELL_X32 FILLER_276_225 ();
 FILLCELL_X32 FILLER_276_257 ();
 FILLCELL_X32 FILLER_276_289 ();
 FILLCELL_X32 FILLER_276_321 ();
 FILLCELL_X32 FILLER_276_353 ();
 FILLCELL_X32 FILLER_276_385 ();
 FILLCELL_X32 FILLER_276_417 ();
 FILLCELL_X32 FILLER_276_449 ();
 FILLCELL_X32 FILLER_276_481 ();
 FILLCELL_X32 FILLER_276_513 ();
 FILLCELL_X32 FILLER_276_545 ();
 FILLCELL_X32 FILLER_276_577 ();
 FILLCELL_X16 FILLER_276_609 ();
 FILLCELL_X4 FILLER_276_625 ();
 FILLCELL_X2 FILLER_276_629 ();
 FILLCELL_X32 FILLER_276_632 ();
 FILLCELL_X32 FILLER_276_664 ();
 FILLCELL_X32 FILLER_276_696 ();
 FILLCELL_X32 FILLER_276_728 ();
 FILLCELL_X32 FILLER_276_760 ();
 FILLCELL_X32 FILLER_276_792 ();
 FILLCELL_X32 FILLER_276_824 ();
 FILLCELL_X32 FILLER_276_856 ();
 FILLCELL_X32 FILLER_276_888 ();
 FILLCELL_X32 FILLER_276_920 ();
 FILLCELL_X32 FILLER_276_952 ();
 FILLCELL_X32 FILLER_276_984 ();
 FILLCELL_X32 FILLER_276_1016 ();
 FILLCELL_X32 FILLER_276_1048 ();
 FILLCELL_X32 FILLER_276_1080 ();
 FILLCELL_X32 FILLER_276_1112 ();
 FILLCELL_X32 FILLER_276_1144 ();
 FILLCELL_X32 FILLER_276_1176 ();
 FILLCELL_X32 FILLER_276_1208 ();
 FILLCELL_X32 FILLER_276_1240 ();
 FILLCELL_X32 FILLER_276_1272 ();
 FILLCELL_X32 FILLER_276_1304 ();
 FILLCELL_X32 FILLER_276_1336 ();
 FILLCELL_X32 FILLER_276_1368 ();
 FILLCELL_X32 FILLER_276_1400 ();
 FILLCELL_X32 FILLER_276_1432 ();
 FILLCELL_X32 FILLER_276_1464 ();
 FILLCELL_X32 FILLER_276_1496 ();
 FILLCELL_X32 FILLER_276_1528 ();
 FILLCELL_X32 FILLER_276_1560 ();
 FILLCELL_X32 FILLER_276_1592 ();
 FILLCELL_X32 FILLER_276_1624 ();
 FILLCELL_X32 FILLER_276_1656 ();
 FILLCELL_X32 FILLER_276_1688 ();
 FILLCELL_X32 FILLER_276_1720 ();
 FILLCELL_X32 FILLER_276_1752 ();
 FILLCELL_X32 FILLER_276_1784 ();
 FILLCELL_X32 FILLER_276_1816 ();
 FILLCELL_X32 FILLER_276_1848 ();
 FILLCELL_X8 FILLER_276_1880 ();
 FILLCELL_X4 FILLER_276_1888 ();
 FILLCELL_X2 FILLER_276_1892 ();
 FILLCELL_X32 FILLER_276_1895 ();
 FILLCELL_X32 FILLER_276_1927 ();
 FILLCELL_X32 FILLER_276_1959 ();
 FILLCELL_X32 FILLER_276_1991 ();
 FILLCELL_X32 FILLER_276_2023 ();
 FILLCELL_X32 FILLER_276_2055 ();
 FILLCELL_X16 FILLER_276_2087 ();
 FILLCELL_X8 FILLER_276_2103 ();
 FILLCELL_X4 FILLER_276_2111 ();
 FILLCELL_X32 FILLER_277_1 ();
 FILLCELL_X32 FILLER_277_33 ();
 FILLCELL_X32 FILLER_277_65 ();
 FILLCELL_X32 FILLER_277_97 ();
 FILLCELL_X32 FILLER_277_129 ();
 FILLCELL_X32 FILLER_277_161 ();
 FILLCELL_X32 FILLER_277_193 ();
 FILLCELL_X32 FILLER_277_225 ();
 FILLCELL_X32 FILLER_277_257 ();
 FILLCELL_X32 FILLER_277_289 ();
 FILLCELL_X32 FILLER_277_321 ();
 FILLCELL_X32 FILLER_277_353 ();
 FILLCELL_X32 FILLER_277_385 ();
 FILLCELL_X32 FILLER_277_417 ();
 FILLCELL_X32 FILLER_277_449 ();
 FILLCELL_X32 FILLER_277_481 ();
 FILLCELL_X32 FILLER_277_513 ();
 FILLCELL_X32 FILLER_277_545 ();
 FILLCELL_X32 FILLER_277_577 ();
 FILLCELL_X32 FILLER_277_609 ();
 FILLCELL_X32 FILLER_277_641 ();
 FILLCELL_X32 FILLER_277_673 ();
 FILLCELL_X32 FILLER_277_705 ();
 FILLCELL_X32 FILLER_277_737 ();
 FILLCELL_X32 FILLER_277_769 ();
 FILLCELL_X32 FILLER_277_801 ();
 FILLCELL_X32 FILLER_277_833 ();
 FILLCELL_X32 FILLER_277_865 ();
 FILLCELL_X32 FILLER_277_897 ();
 FILLCELL_X32 FILLER_277_929 ();
 FILLCELL_X32 FILLER_277_961 ();
 FILLCELL_X32 FILLER_277_993 ();
 FILLCELL_X32 FILLER_277_1025 ();
 FILLCELL_X32 FILLER_277_1057 ();
 FILLCELL_X32 FILLER_277_1089 ();
 FILLCELL_X32 FILLER_277_1121 ();
 FILLCELL_X32 FILLER_277_1153 ();
 FILLCELL_X32 FILLER_277_1185 ();
 FILLCELL_X32 FILLER_277_1217 ();
 FILLCELL_X8 FILLER_277_1249 ();
 FILLCELL_X4 FILLER_277_1257 ();
 FILLCELL_X2 FILLER_277_1261 ();
 FILLCELL_X32 FILLER_277_1264 ();
 FILLCELL_X32 FILLER_277_1296 ();
 FILLCELL_X32 FILLER_277_1328 ();
 FILLCELL_X32 FILLER_277_1360 ();
 FILLCELL_X32 FILLER_277_1392 ();
 FILLCELL_X32 FILLER_277_1424 ();
 FILLCELL_X32 FILLER_277_1456 ();
 FILLCELL_X32 FILLER_277_1488 ();
 FILLCELL_X32 FILLER_277_1520 ();
 FILLCELL_X32 FILLER_277_1552 ();
 FILLCELL_X32 FILLER_277_1584 ();
 FILLCELL_X32 FILLER_277_1616 ();
 FILLCELL_X32 FILLER_277_1648 ();
 FILLCELL_X32 FILLER_277_1680 ();
 FILLCELL_X32 FILLER_277_1712 ();
 FILLCELL_X32 FILLER_277_1744 ();
 FILLCELL_X32 FILLER_277_1776 ();
 FILLCELL_X32 FILLER_277_1808 ();
 FILLCELL_X32 FILLER_277_1840 ();
 FILLCELL_X32 FILLER_277_1872 ();
 FILLCELL_X32 FILLER_277_1904 ();
 FILLCELL_X32 FILLER_277_1936 ();
 FILLCELL_X32 FILLER_277_1968 ();
 FILLCELL_X32 FILLER_277_2000 ();
 FILLCELL_X32 FILLER_277_2032 ();
 FILLCELL_X32 FILLER_277_2064 ();
 FILLCELL_X16 FILLER_277_2096 ();
 FILLCELL_X2 FILLER_277_2112 ();
 FILLCELL_X1 FILLER_277_2114 ();
 FILLCELL_X32 FILLER_278_1 ();
 FILLCELL_X32 FILLER_278_33 ();
 FILLCELL_X32 FILLER_278_65 ();
 FILLCELL_X32 FILLER_278_97 ();
 FILLCELL_X32 FILLER_278_129 ();
 FILLCELL_X32 FILLER_278_161 ();
 FILLCELL_X32 FILLER_278_193 ();
 FILLCELL_X32 FILLER_278_225 ();
 FILLCELL_X32 FILLER_278_257 ();
 FILLCELL_X32 FILLER_278_289 ();
 FILLCELL_X32 FILLER_278_321 ();
 FILLCELL_X32 FILLER_278_353 ();
 FILLCELL_X32 FILLER_278_385 ();
 FILLCELL_X32 FILLER_278_417 ();
 FILLCELL_X32 FILLER_278_449 ();
 FILLCELL_X32 FILLER_278_481 ();
 FILLCELL_X32 FILLER_278_513 ();
 FILLCELL_X32 FILLER_278_545 ();
 FILLCELL_X32 FILLER_278_577 ();
 FILLCELL_X16 FILLER_278_609 ();
 FILLCELL_X4 FILLER_278_625 ();
 FILLCELL_X2 FILLER_278_629 ();
 FILLCELL_X32 FILLER_278_632 ();
 FILLCELL_X32 FILLER_278_664 ();
 FILLCELL_X32 FILLER_278_696 ();
 FILLCELL_X32 FILLER_278_728 ();
 FILLCELL_X32 FILLER_278_760 ();
 FILLCELL_X32 FILLER_278_792 ();
 FILLCELL_X32 FILLER_278_824 ();
 FILLCELL_X32 FILLER_278_856 ();
 FILLCELL_X32 FILLER_278_888 ();
 FILLCELL_X32 FILLER_278_920 ();
 FILLCELL_X32 FILLER_278_952 ();
 FILLCELL_X32 FILLER_278_984 ();
 FILLCELL_X32 FILLER_278_1016 ();
 FILLCELL_X32 FILLER_278_1048 ();
 FILLCELL_X32 FILLER_278_1080 ();
 FILLCELL_X32 FILLER_278_1112 ();
 FILLCELL_X32 FILLER_278_1144 ();
 FILLCELL_X32 FILLER_278_1176 ();
 FILLCELL_X32 FILLER_278_1208 ();
 FILLCELL_X32 FILLER_278_1240 ();
 FILLCELL_X32 FILLER_278_1272 ();
 FILLCELL_X32 FILLER_278_1304 ();
 FILLCELL_X32 FILLER_278_1336 ();
 FILLCELL_X32 FILLER_278_1368 ();
 FILLCELL_X32 FILLER_278_1400 ();
 FILLCELL_X32 FILLER_278_1432 ();
 FILLCELL_X32 FILLER_278_1464 ();
 FILLCELL_X32 FILLER_278_1496 ();
 FILLCELL_X32 FILLER_278_1528 ();
 FILLCELL_X32 FILLER_278_1560 ();
 FILLCELL_X32 FILLER_278_1592 ();
 FILLCELL_X32 FILLER_278_1624 ();
 FILLCELL_X32 FILLER_278_1656 ();
 FILLCELL_X32 FILLER_278_1688 ();
 FILLCELL_X32 FILLER_278_1720 ();
 FILLCELL_X32 FILLER_278_1752 ();
 FILLCELL_X32 FILLER_278_1784 ();
 FILLCELL_X32 FILLER_278_1816 ();
 FILLCELL_X32 FILLER_278_1848 ();
 FILLCELL_X8 FILLER_278_1880 ();
 FILLCELL_X4 FILLER_278_1888 ();
 FILLCELL_X2 FILLER_278_1892 ();
 FILLCELL_X32 FILLER_278_1895 ();
 FILLCELL_X32 FILLER_278_1927 ();
 FILLCELL_X32 FILLER_278_1959 ();
 FILLCELL_X32 FILLER_278_1991 ();
 FILLCELL_X32 FILLER_278_2023 ();
 FILLCELL_X32 FILLER_278_2055 ();
 FILLCELL_X16 FILLER_278_2087 ();
 FILLCELL_X8 FILLER_278_2103 ();
 FILLCELL_X4 FILLER_278_2111 ();
 FILLCELL_X32 FILLER_279_1 ();
 FILLCELL_X32 FILLER_279_33 ();
 FILLCELL_X32 FILLER_279_65 ();
 FILLCELL_X32 FILLER_279_97 ();
 FILLCELL_X32 FILLER_279_129 ();
 FILLCELL_X32 FILLER_279_161 ();
 FILLCELL_X32 FILLER_279_193 ();
 FILLCELL_X32 FILLER_279_225 ();
 FILLCELL_X32 FILLER_279_257 ();
 FILLCELL_X32 FILLER_279_289 ();
 FILLCELL_X32 FILLER_279_321 ();
 FILLCELL_X32 FILLER_279_353 ();
 FILLCELL_X32 FILLER_279_385 ();
 FILLCELL_X32 FILLER_279_417 ();
 FILLCELL_X32 FILLER_279_449 ();
 FILLCELL_X32 FILLER_279_481 ();
 FILLCELL_X32 FILLER_279_513 ();
 FILLCELL_X32 FILLER_279_545 ();
 FILLCELL_X32 FILLER_279_577 ();
 FILLCELL_X32 FILLER_279_609 ();
 FILLCELL_X32 FILLER_279_641 ();
 FILLCELL_X32 FILLER_279_673 ();
 FILLCELL_X32 FILLER_279_705 ();
 FILLCELL_X32 FILLER_279_737 ();
 FILLCELL_X32 FILLER_279_769 ();
 FILLCELL_X32 FILLER_279_801 ();
 FILLCELL_X32 FILLER_279_833 ();
 FILLCELL_X32 FILLER_279_865 ();
 FILLCELL_X32 FILLER_279_897 ();
 FILLCELL_X32 FILLER_279_929 ();
 FILLCELL_X32 FILLER_279_961 ();
 FILLCELL_X32 FILLER_279_993 ();
 FILLCELL_X32 FILLER_279_1025 ();
 FILLCELL_X32 FILLER_279_1057 ();
 FILLCELL_X32 FILLER_279_1089 ();
 FILLCELL_X32 FILLER_279_1121 ();
 FILLCELL_X32 FILLER_279_1153 ();
 FILLCELL_X32 FILLER_279_1185 ();
 FILLCELL_X32 FILLER_279_1217 ();
 FILLCELL_X8 FILLER_279_1249 ();
 FILLCELL_X4 FILLER_279_1257 ();
 FILLCELL_X2 FILLER_279_1261 ();
 FILLCELL_X32 FILLER_279_1264 ();
 FILLCELL_X32 FILLER_279_1296 ();
 FILLCELL_X32 FILLER_279_1328 ();
 FILLCELL_X32 FILLER_279_1360 ();
 FILLCELL_X32 FILLER_279_1392 ();
 FILLCELL_X32 FILLER_279_1424 ();
 FILLCELL_X32 FILLER_279_1456 ();
 FILLCELL_X32 FILLER_279_1488 ();
 FILLCELL_X32 FILLER_279_1520 ();
 FILLCELL_X32 FILLER_279_1552 ();
 FILLCELL_X32 FILLER_279_1584 ();
 FILLCELL_X32 FILLER_279_1616 ();
 FILLCELL_X32 FILLER_279_1648 ();
 FILLCELL_X32 FILLER_279_1680 ();
 FILLCELL_X32 FILLER_279_1712 ();
 FILLCELL_X32 FILLER_279_1744 ();
 FILLCELL_X32 FILLER_279_1776 ();
 FILLCELL_X32 FILLER_279_1808 ();
 FILLCELL_X32 FILLER_279_1840 ();
 FILLCELL_X32 FILLER_279_1872 ();
 FILLCELL_X32 FILLER_279_1904 ();
 FILLCELL_X32 FILLER_279_1936 ();
 FILLCELL_X32 FILLER_279_1968 ();
 FILLCELL_X32 FILLER_279_2000 ();
 FILLCELL_X32 FILLER_279_2032 ();
 FILLCELL_X32 FILLER_279_2064 ();
 FILLCELL_X16 FILLER_279_2096 ();
 FILLCELL_X2 FILLER_279_2112 ();
 FILLCELL_X1 FILLER_279_2114 ();
 FILLCELL_X32 FILLER_280_1 ();
 FILLCELL_X32 FILLER_280_33 ();
 FILLCELL_X32 FILLER_280_65 ();
 FILLCELL_X32 FILLER_280_97 ();
 FILLCELL_X32 FILLER_280_129 ();
 FILLCELL_X32 FILLER_280_161 ();
 FILLCELL_X32 FILLER_280_193 ();
 FILLCELL_X32 FILLER_280_225 ();
 FILLCELL_X32 FILLER_280_257 ();
 FILLCELL_X32 FILLER_280_289 ();
 FILLCELL_X32 FILLER_280_321 ();
 FILLCELL_X32 FILLER_280_353 ();
 FILLCELL_X32 FILLER_280_385 ();
 FILLCELL_X32 FILLER_280_417 ();
 FILLCELL_X32 FILLER_280_449 ();
 FILLCELL_X32 FILLER_280_481 ();
 FILLCELL_X32 FILLER_280_513 ();
 FILLCELL_X32 FILLER_280_545 ();
 FILLCELL_X32 FILLER_280_577 ();
 FILLCELL_X16 FILLER_280_609 ();
 FILLCELL_X4 FILLER_280_625 ();
 FILLCELL_X2 FILLER_280_629 ();
 FILLCELL_X32 FILLER_280_632 ();
 FILLCELL_X32 FILLER_280_664 ();
 FILLCELL_X32 FILLER_280_696 ();
 FILLCELL_X32 FILLER_280_728 ();
 FILLCELL_X32 FILLER_280_760 ();
 FILLCELL_X32 FILLER_280_792 ();
 FILLCELL_X32 FILLER_280_824 ();
 FILLCELL_X32 FILLER_280_856 ();
 FILLCELL_X32 FILLER_280_888 ();
 FILLCELL_X32 FILLER_280_920 ();
 FILLCELL_X32 FILLER_280_952 ();
 FILLCELL_X32 FILLER_280_984 ();
 FILLCELL_X32 FILLER_280_1016 ();
 FILLCELL_X32 FILLER_280_1048 ();
 FILLCELL_X32 FILLER_280_1080 ();
 FILLCELL_X32 FILLER_280_1112 ();
 FILLCELL_X32 FILLER_280_1144 ();
 FILLCELL_X32 FILLER_280_1176 ();
 FILLCELL_X32 FILLER_280_1208 ();
 FILLCELL_X32 FILLER_280_1240 ();
 FILLCELL_X32 FILLER_280_1272 ();
 FILLCELL_X32 FILLER_280_1304 ();
 FILLCELL_X32 FILLER_280_1336 ();
 FILLCELL_X32 FILLER_280_1368 ();
 FILLCELL_X32 FILLER_280_1400 ();
 FILLCELL_X32 FILLER_280_1432 ();
 FILLCELL_X32 FILLER_280_1464 ();
 FILLCELL_X32 FILLER_280_1496 ();
 FILLCELL_X32 FILLER_280_1528 ();
 FILLCELL_X32 FILLER_280_1560 ();
 FILLCELL_X32 FILLER_280_1592 ();
 FILLCELL_X32 FILLER_280_1624 ();
 FILLCELL_X32 FILLER_280_1656 ();
 FILLCELL_X32 FILLER_280_1688 ();
 FILLCELL_X32 FILLER_280_1720 ();
 FILLCELL_X32 FILLER_280_1752 ();
 FILLCELL_X32 FILLER_280_1784 ();
 FILLCELL_X32 FILLER_280_1816 ();
 FILLCELL_X32 FILLER_280_1848 ();
 FILLCELL_X8 FILLER_280_1880 ();
 FILLCELL_X4 FILLER_280_1888 ();
 FILLCELL_X2 FILLER_280_1892 ();
 FILLCELL_X32 FILLER_280_1895 ();
 FILLCELL_X32 FILLER_280_1927 ();
 FILLCELL_X32 FILLER_280_1959 ();
 FILLCELL_X32 FILLER_280_1991 ();
 FILLCELL_X32 FILLER_280_2023 ();
 FILLCELL_X32 FILLER_280_2055 ();
 FILLCELL_X16 FILLER_280_2087 ();
 FILLCELL_X8 FILLER_280_2103 ();
 FILLCELL_X4 FILLER_280_2111 ();
 FILLCELL_X32 FILLER_281_1 ();
 FILLCELL_X32 FILLER_281_33 ();
 FILLCELL_X32 FILLER_281_65 ();
 FILLCELL_X32 FILLER_281_97 ();
 FILLCELL_X32 FILLER_281_129 ();
 FILLCELL_X32 FILLER_281_161 ();
 FILLCELL_X32 FILLER_281_193 ();
 FILLCELL_X32 FILLER_281_225 ();
 FILLCELL_X32 FILLER_281_257 ();
 FILLCELL_X32 FILLER_281_289 ();
 FILLCELL_X32 FILLER_281_321 ();
 FILLCELL_X32 FILLER_281_353 ();
 FILLCELL_X32 FILLER_281_385 ();
 FILLCELL_X32 FILLER_281_417 ();
 FILLCELL_X32 FILLER_281_449 ();
 FILLCELL_X32 FILLER_281_481 ();
 FILLCELL_X32 FILLER_281_513 ();
 FILLCELL_X32 FILLER_281_545 ();
 FILLCELL_X32 FILLER_281_577 ();
 FILLCELL_X32 FILLER_281_609 ();
 FILLCELL_X32 FILLER_281_641 ();
 FILLCELL_X32 FILLER_281_673 ();
 FILLCELL_X32 FILLER_281_705 ();
 FILLCELL_X32 FILLER_281_737 ();
 FILLCELL_X32 FILLER_281_769 ();
 FILLCELL_X32 FILLER_281_801 ();
 FILLCELL_X32 FILLER_281_833 ();
 FILLCELL_X32 FILLER_281_865 ();
 FILLCELL_X32 FILLER_281_897 ();
 FILLCELL_X32 FILLER_281_929 ();
 FILLCELL_X32 FILLER_281_961 ();
 FILLCELL_X32 FILLER_281_993 ();
 FILLCELL_X32 FILLER_281_1025 ();
 FILLCELL_X32 FILLER_281_1057 ();
 FILLCELL_X32 FILLER_281_1089 ();
 FILLCELL_X32 FILLER_281_1121 ();
 FILLCELL_X32 FILLER_281_1153 ();
 FILLCELL_X32 FILLER_281_1185 ();
 FILLCELL_X32 FILLER_281_1217 ();
 FILLCELL_X8 FILLER_281_1249 ();
 FILLCELL_X4 FILLER_281_1257 ();
 FILLCELL_X2 FILLER_281_1261 ();
 FILLCELL_X32 FILLER_281_1264 ();
 FILLCELL_X32 FILLER_281_1296 ();
 FILLCELL_X32 FILLER_281_1328 ();
 FILLCELL_X32 FILLER_281_1360 ();
 FILLCELL_X32 FILLER_281_1392 ();
 FILLCELL_X32 FILLER_281_1424 ();
 FILLCELL_X32 FILLER_281_1456 ();
 FILLCELL_X32 FILLER_281_1488 ();
 FILLCELL_X32 FILLER_281_1520 ();
 FILLCELL_X32 FILLER_281_1552 ();
 FILLCELL_X32 FILLER_281_1584 ();
 FILLCELL_X32 FILLER_281_1616 ();
 FILLCELL_X32 FILLER_281_1648 ();
 FILLCELL_X32 FILLER_281_1680 ();
 FILLCELL_X32 FILLER_281_1712 ();
 FILLCELL_X32 FILLER_281_1744 ();
 FILLCELL_X32 FILLER_281_1776 ();
 FILLCELL_X32 FILLER_281_1808 ();
 FILLCELL_X32 FILLER_281_1840 ();
 FILLCELL_X32 FILLER_281_1872 ();
 FILLCELL_X32 FILLER_281_1904 ();
 FILLCELL_X32 FILLER_281_1936 ();
 FILLCELL_X32 FILLER_281_1968 ();
 FILLCELL_X32 FILLER_281_2000 ();
 FILLCELL_X32 FILLER_281_2032 ();
 FILLCELL_X32 FILLER_281_2064 ();
 FILLCELL_X16 FILLER_281_2096 ();
 FILLCELL_X2 FILLER_281_2112 ();
 FILLCELL_X1 FILLER_281_2114 ();
 FILLCELL_X32 FILLER_282_1 ();
 FILLCELL_X32 FILLER_282_33 ();
 FILLCELL_X32 FILLER_282_65 ();
 FILLCELL_X32 FILLER_282_97 ();
 FILLCELL_X32 FILLER_282_129 ();
 FILLCELL_X32 FILLER_282_161 ();
 FILLCELL_X32 FILLER_282_193 ();
 FILLCELL_X32 FILLER_282_225 ();
 FILLCELL_X32 FILLER_282_257 ();
 FILLCELL_X32 FILLER_282_289 ();
 FILLCELL_X32 FILLER_282_321 ();
 FILLCELL_X32 FILLER_282_353 ();
 FILLCELL_X32 FILLER_282_385 ();
 FILLCELL_X32 FILLER_282_417 ();
 FILLCELL_X32 FILLER_282_449 ();
 FILLCELL_X32 FILLER_282_481 ();
 FILLCELL_X32 FILLER_282_513 ();
 FILLCELL_X32 FILLER_282_545 ();
 FILLCELL_X32 FILLER_282_577 ();
 FILLCELL_X16 FILLER_282_609 ();
 FILLCELL_X4 FILLER_282_625 ();
 FILLCELL_X2 FILLER_282_629 ();
 FILLCELL_X32 FILLER_282_632 ();
 FILLCELL_X32 FILLER_282_664 ();
 FILLCELL_X32 FILLER_282_696 ();
 FILLCELL_X32 FILLER_282_728 ();
 FILLCELL_X32 FILLER_282_760 ();
 FILLCELL_X32 FILLER_282_792 ();
 FILLCELL_X32 FILLER_282_824 ();
 FILLCELL_X32 FILLER_282_856 ();
 FILLCELL_X32 FILLER_282_888 ();
 FILLCELL_X32 FILLER_282_920 ();
 FILLCELL_X32 FILLER_282_952 ();
 FILLCELL_X32 FILLER_282_984 ();
 FILLCELL_X32 FILLER_282_1016 ();
 FILLCELL_X32 FILLER_282_1048 ();
 FILLCELL_X32 FILLER_282_1080 ();
 FILLCELL_X32 FILLER_282_1112 ();
 FILLCELL_X32 FILLER_282_1144 ();
 FILLCELL_X32 FILLER_282_1176 ();
 FILLCELL_X32 FILLER_282_1208 ();
 FILLCELL_X32 FILLER_282_1240 ();
 FILLCELL_X32 FILLER_282_1272 ();
 FILLCELL_X32 FILLER_282_1304 ();
 FILLCELL_X32 FILLER_282_1336 ();
 FILLCELL_X32 FILLER_282_1368 ();
 FILLCELL_X32 FILLER_282_1400 ();
 FILLCELL_X32 FILLER_282_1432 ();
 FILLCELL_X32 FILLER_282_1464 ();
 FILLCELL_X32 FILLER_282_1496 ();
 FILLCELL_X32 FILLER_282_1528 ();
 FILLCELL_X32 FILLER_282_1560 ();
 FILLCELL_X32 FILLER_282_1592 ();
 FILLCELL_X32 FILLER_282_1624 ();
 FILLCELL_X32 FILLER_282_1656 ();
 FILLCELL_X32 FILLER_282_1688 ();
 FILLCELL_X32 FILLER_282_1720 ();
 FILLCELL_X32 FILLER_282_1752 ();
 FILLCELL_X32 FILLER_282_1784 ();
 FILLCELL_X32 FILLER_282_1816 ();
 FILLCELL_X32 FILLER_282_1848 ();
 FILLCELL_X8 FILLER_282_1880 ();
 FILLCELL_X4 FILLER_282_1888 ();
 FILLCELL_X2 FILLER_282_1892 ();
 FILLCELL_X32 FILLER_282_1895 ();
 FILLCELL_X32 FILLER_282_1927 ();
 FILLCELL_X32 FILLER_282_1959 ();
 FILLCELL_X32 FILLER_282_1991 ();
 FILLCELL_X32 FILLER_282_2023 ();
 FILLCELL_X32 FILLER_282_2055 ();
 FILLCELL_X16 FILLER_282_2087 ();
 FILLCELL_X8 FILLER_282_2103 ();
 FILLCELL_X4 FILLER_282_2111 ();
 FILLCELL_X32 FILLER_283_1 ();
 FILLCELL_X32 FILLER_283_33 ();
 FILLCELL_X32 FILLER_283_65 ();
 FILLCELL_X32 FILLER_283_97 ();
 FILLCELL_X32 FILLER_283_129 ();
 FILLCELL_X32 FILLER_283_161 ();
 FILLCELL_X32 FILLER_283_193 ();
 FILLCELL_X32 FILLER_283_225 ();
 FILLCELL_X32 FILLER_283_257 ();
 FILLCELL_X32 FILLER_283_289 ();
 FILLCELL_X32 FILLER_283_321 ();
 FILLCELL_X32 FILLER_283_353 ();
 FILLCELL_X32 FILLER_283_385 ();
 FILLCELL_X32 FILLER_283_417 ();
 FILLCELL_X32 FILLER_283_449 ();
 FILLCELL_X32 FILLER_283_481 ();
 FILLCELL_X32 FILLER_283_513 ();
 FILLCELL_X32 FILLER_283_545 ();
 FILLCELL_X32 FILLER_283_577 ();
 FILLCELL_X32 FILLER_283_609 ();
 FILLCELL_X32 FILLER_283_641 ();
 FILLCELL_X32 FILLER_283_673 ();
 FILLCELL_X32 FILLER_283_705 ();
 FILLCELL_X32 FILLER_283_737 ();
 FILLCELL_X32 FILLER_283_769 ();
 FILLCELL_X32 FILLER_283_801 ();
 FILLCELL_X32 FILLER_283_833 ();
 FILLCELL_X32 FILLER_283_865 ();
 FILLCELL_X32 FILLER_283_897 ();
 FILLCELL_X32 FILLER_283_929 ();
 FILLCELL_X32 FILLER_283_961 ();
 FILLCELL_X32 FILLER_283_993 ();
 FILLCELL_X32 FILLER_283_1025 ();
 FILLCELL_X32 FILLER_283_1057 ();
 FILLCELL_X32 FILLER_283_1089 ();
 FILLCELL_X32 FILLER_283_1121 ();
 FILLCELL_X32 FILLER_283_1153 ();
 FILLCELL_X16 FILLER_283_1185 ();
 FILLCELL_X4 FILLER_283_1201 ();
 FILLCELL_X2 FILLER_283_1205 ();
 FILLCELL_X32 FILLER_283_1209 ();
 FILLCELL_X16 FILLER_283_1241 ();
 FILLCELL_X4 FILLER_283_1257 ();
 FILLCELL_X2 FILLER_283_1261 ();
 FILLCELL_X32 FILLER_283_1264 ();
 FILLCELL_X32 FILLER_283_1296 ();
 FILLCELL_X32 FILLER_283_1328 ();
 FILLCELL_X32 FILLER_283_1360 ();
 FILLCELL_X32 FILLER_283_1392 ();
 FILLCELL_X32 FILLER_283_1424 ();
 FILLCELL_X32 FILLER_283_1456 ();
 FILLCELL_X32 FILLER_283_1488 ();
 FILLCELL_X32 FILLER_283_1520 ();
 FILLCELL_X32 FILLER_283_1552 ();
 FILLCELL_X32 FILLER_283_1584 ();
 FILLCELL_X32 FILLER_283_1616 ();
 FILLCELL_X32 FILLER_283_1648 ();
 FILLCELL_X32 FILLER_283_1680 ();
 FILLCELL_X32 FILLER_283_1712 ();
 FILLCELL_X32 FILLER_283_1744 ();
 FILLCELL_X32 FILLER_283_1776 ();
 FILLCELL_X32 FILLER_283_1808 ();
 FILLCELL_X32 FILLER_283_1840 ();
 FILLCELL_X32 FILLER_283_1872 ();
 FILLCELL_X32 FILLER_283_1904 ();
 FILLCELL_X32 FILLER_283_1936 ();
 FILLCELL_X32 FILLER_283_1968 ();
 FILLCELL_X32 FILLER_283_2000 ();
 FILLCELL_X32 FILLER_283_2032 ();
 FILLCELL_X32 FILLER_283_2064 ();
 FILLCELL_X16 FILLER_283_2096 ();
 FILLCELL_X2 FILLER_283_2112 ();
 FILLCELL_X1 FILLER_283_2114 ();
 FILLCELL_X32 FILLER_284_1 ();
 FILLCELL_X32 FILLER_284_33 ();
 FILLCELL_X32 FILLER_284_65 ();
 FILLCELL_X32 FILLER_284_97 ();
 FILLCELL_X32 FILLER_284_129 ();
 FILLCELL_X32 FILLER_284_161 ();
 FILLCELL_X32 FILLER_284_193 ();
 FILLCELL_X32 FILLER_284_225 ();
 FILLCELL_X32 FILLER_284_257 ();
 FILLCELL_X32 FILLER_284_289 ();
 FILLCELL_X32 FILLER_284_321 ();
 FILLCELL_X32 FILLER_284_353 ();
 FILLCELL_X32 FILLER_284_385 ();
 FILLCELL_X32 FILLER_284_417 ();
 FILLCELL_X32 FILLER_284_449 ();
 FILLCELL_X32 FILLER_284_481 ();
 FILLCELL_X32 FILLER_284_513 ();
 FILLCELL_X32 FILLER_284_545 ();
 FILLCELL_X32 FILLER_284_577 ();
 FILLCELL_X16 FILLER_284_609 ();
 FILLCELL_X4 FILLER_284_625 ();
 FILLCELL_X2 FILLER_284_629 ();
 FILLCELL_X32 FILLER_284_632 ();
 FILLCELL_X32 FILLER_284_664 ();
 FILLCELL_X32 FILLER_284_696 ();
 FILLCELL_X32 FILLER_284_728 ();
 FILLCELL_X32 FILLER_284_760 ();
 FILLCELL_X32 FILLER_284_792 ();
 FILLCELL_X32 FILLER_284_824 ();
 FILLCELL_X32 FILLER_284_856 ();
 FILLCELL_X32 FILLER_284_888 ();
 FILLCELL_X32 FILLER_284_920 ();
 FILLCELL_X32 FILLER_284_952 ();
 FILLCELL_X32 FILLER_284_984 ();
 FILLCELL_X32 FILLER_284_1016 ();
 FILLCELL_X32 FILLER_284_1048 ();
 FILLCELL_X32 FILLER_284_1080 ();
 FILLCELL_X32 FILLER_284_1112 ();
 FILLCELL_X32 FILLER_284_1144 ();
 FILLCELL_X16 FILLER_284_1176 ();
 FILLCELL_X2 FILLER_284_1192 ();
 FILLCELL_X1 FILLER_284_1194 ();
 FILLCELL_X4 FILLER_284_1197 ();
 FILLCELL_X1 FILLER_284_1201 ();
 FILLCELL_X8 FILLER_284_1207 ();
 FILLCELL_X32 FILLER_284_1220 ();
 FILLCELL_X32 FILLER_284_1252 ();
 FILLCELL_X32 FILLER_284_1284 ();
 FILLCELL_X32 FILLER_284_1316 ();
 FILLCELL_X32 FILLER_284_1348 ();
 FILLCELL_X32 FILLER_284_1380 ();
 FILLCELL_X32 FILLER_284_1412 ();
 FILLCELL_X32 FILLER_284_1444 ();
 FILLCELL_X32 FILLER_284_1476 ();
 FILLCELL_X32 FILLER_284_1508 ();
 FILLCELL_X32 FILLER_284_1540 ();
 FILLCELL_X32 FILLER_284_1572 ();
 FILLCELL_X32 FILLER_284_1604 ();
 FILLCELL_X32 FILLER_284_1636 ();
 FILLCELL_X32 FILLER_284_1668 ();
 FILLCELL_X32 FILLER_284_1700 ();
 FILLCELL_X32 FILLER_284_1732 ();
 FILLCELL_X32 FILLER_284_1764 ();
 FILLCELL_X32 FILLER_284_1796 ();
 FILLCELL_X32 FILLER_284_1828 ();
 FILLCELL_X32 FILLER_284_1860 ();
 FILLCELL_X2 FILLER_284_1892 ();
 FILLCELL_X32 FILLER_284_1895 ();
 FILLCELL_X32 FILLER_284_1927 ();
 FILLCELL_X32 FILLER_284_1959 ();
 FILLCELL_X32 FILLER_284_1991 ();
 FILLCELL_X32 FILLER_284_2023 ();
 FILLCELL_X32 FILLER_284_2055 ();
 FILLCELL_X16 FILLER_284_2087 ();
 FILLCELL_X8 FILLER_284_2103 ();
 FILLCELL_X4 FILLER_284_2111 ();
 FILLCELL_X32 FILLER_285_1 ();
 FILLCELL_X32 FILLER_285_33 ();
 FILLCELL_X32 FILLER_285_65 ();
 FILLCELL_X32 FILLER_285_97 ();
 FILLCELL_X32 FILLER_285_129 ();
 FILLCELL_X32 FILLER_285_161 ();
 FILLCELL_X32 FILLER_285_193 ();
 FILLCELL_X32 FILLER_285_225 ();
 FILLCELL_X32 FILLER_285_257 ();
 FILLCELL_X32 FILLER_285_289 ();
 FILLCELL_X32 FILLER_285_321 ();
 FILLCELL_X32 FILLER_285_353 ();
 FILLCELL_X32 FILLER_285_385 ();
 FILLCELL_X32 FILLER_285_417 ();
 FILLCELL_X32 FILLER_285_449 ();
 FILLCELL_X32 FILLER_285_481 ();
 FILLCELL_X32 FILLER_285_513 ();
 FILLCELL_X32 FILLER_285_545 ();
 FILLCELL_X32 FILLER_285_577 ();
 FILLCELL_X32 FILLER_285_609 ();
 FILLCELL_X32 FILLER_285_641 ();
 FILLCELL_X32 FILLER_285_673 ();
 FILLCELL_X32 FILLER_285_705 ();
 FILLCELL_X32 FILLER_285_737 ();
 FILLCELL_X32 FILLER_285_769 ();
 FILLCELL_X32 FILLER_285_801 ();
 FILLCELL_X32 FILLER_285_833 ();
 FILLCELL_X32 FILLER_285_865 ();
 FILLCELL_X32 FILLER_285_897 ();
 FILLCELL_X32 FILLER_285_929 ();
 FILLCELL_X32 FILLER_285_961 ();
 FILLCELL_X32 FILLER_285_993 ();
 FILLCELL_X32 FILLER_285_1025 ();
 FILLCELL_X32 FILLER_285_1057 ();
 FILLCELL_X32 FILLER_285_1089 ();
 FILLCELL_X2 FILLER_285_1121 ();
 FILLCELL_X8 FILLER_285_1126 ();
 FILLCELL_X4 FILLER_285_1134 ();
 FILLCELL_X2 FILLER_285_1138 ();
 FILLCELL_X1 FILLER_285_1140 ();
 FILLCELL_X32 FILLER_285_1144 ();
 FILLCELL_X32 FILLER_285_1176 ();
 FILLCELL_X32 FILLER_285_1221 ();
 FILLCELL_X8 FILLER_285_1253 ();
 FILLCELL_X2 FILLER_285_1261 ();
 FILLCELL_X32 FILLER_285_1264 ();
 FILLCELL_X32 FILLER_285_1296 ();
 FILLCELL_X32 FILLER_285_1328 ();
 FILLCELL_X32 FILLER_285_1360 ();
 FILLCELL_X32 FILLER_285_1392 ();
 FILLCELL_X32 FILLER_285_1424 ();
 FILLCELL_X32 FILLER_285_1456 ();
 FILLCELL_X32 FILLER_285_1488 ();
 FILLCELL_X32 FILLER_285_1520 ();
 FILLCELL_X32 FILLER_285_1552 ();
 FILLCELL_X32 FILLER_285_1584 ();
 FILLCELL_X32 FILLER_285_1616 ();
 FILLCELL_X32 FILLER_285_1648 ();
 FILLCELL_X32 FILLER_285_1680 ();
 FILLCELL_X32 FILLER_285_1712 ();
 FILLCELL_X32 FILLER_285_1744 ();
 FILLCELL_X32 FILLER_285_1776 ();
 FILLCELL_X32 FILLER_285_1808 ();
 FILLCELL_X32 FILLER_285_1840 ();
 FILLCELL_X32 FILLER_285_1872 ();
 FILLCELL_X32 FILLER_285_1904 ();
 FILLCELL_X32 FILLER_285_1936 ();
 FILLCELL_X32 FILLER_285_1968 ();
 FILLCELL_X32 FILLER_285_2000 ();
 FILLCELL_X32 FILLER_285_2032 ();
 FILLCELL_X32 FILLER_285_2064 ();
 FILLCELL_X16 FILLER_285_2096 ();
 FILLCELL_X2 FILLER_285_2112 ();
 FILLCELL_X1 FILLER_285_2114 ();
 FILLCELL_X32 FILLER_286_1 ();
 FILLCELL_X32 FILLER_286_33 ();
 FILLCELL_X32 FILLER_286_65 ();
 FILLCELL_X32 FILLER_286_97 ();
 FILLCELL_X32 FILLER_286_129 ();
 FILLCELL_X32 FILLER_286_161 ();
 FILLCELL_X32 FILLER_286_193 ();
 FILLCELL_X32 FILLER_286_225 ();
 FILLCELL_X32 FILLER_286_257 ();
 FILLCELL_X32 FILLER_286_289 ();
 FILLCELL_X32 FILLER_286_321 ();
 FILLCELL_X32 FILLER_286_353 ();
 FILLCELL_X32 FILLER_286_385 ();
 FILLCELL_X32 FILLER_286_417 ();
 FILLCELL_X32 FILLER_286_449 ();
 FILLCELL_X32 FILLER_286_481 ();
 FILLCELL_X32 FILLER_286_513 ();
 FILLCELL_X32 FILLER_286_545 ();
 FILLCELL_X32 FILLER_286_577 ();
 FILLCELL_X16 FILLER_286_609 ();
 FILLCELL_X4 FILLER_286_625 ();
 FILLCELL_X2 FILLER_286_629 ();
 FILLCELL_X32 FILLER_286_632 ();
 FILLCELL_X32 FILLER_286_664 ();
 FILLCELL_X32 FILLER_286_696 ();
 FILLCELL_X32 FILLER_286_728 ();
 FILLCELL_X32 FILLER_286_760 ();
 FILLCELL_X32 FILLER_286_792 ();
 FILLCELL_X32 FILLER_286_824 ();
 FILLCELL_X32 FILLER_286_856 ();
 FILLCELL_X32 FILLER_286_888 ();
 FILLCELL_X32 FILLER_286_920 ();
 FILLCELL_X32 FILLER_286_952 ();
 FILLCELL_X32 FILLER_286_984 ();
 FILLCELL_X32 FILLER_286_1016 ();
 FILLCELL_X32 FILLER_286_1048 ();
 FILLCELL_X16 FILLER_286_1080 ();
 FILLCELL_X8 FILLER_286_1096 ();
 FILLCELL_X4 FILLER_286_1104 ();
 FILLCELL_X1 FILLER_286_1108 ();
 FILLCELL_X32 FILLER_286_1121 ();
 FILLCELL_X32 FILLER_286_1153 ();
 FILLCELL_X8 FILLER_286_1185 ();
 FILLCELL_X1 FILLER_286_1193 ();
 FILLCELL_X2 FILLER_286_1197 ();
 FILLCELL_X1 FILLER_286_1199 ();
 FILLCELL_X1 FILLER_286_1216 ();
 FILLCELL_X8 FILLER_286_1220 ();
 FILLCELL_X1 FILLER_286_1228 ();
 FILLCELL_X16 FILLER_286_1242 ();
 FILLCELL_X4 FILLER_286_1258 ();
 FILLCELL_X32 FILLER_286_1263 ();
 FILLCELL_X32 FILLER_286_1295 ();
 FILLCELL_X32 FILLER_286_1327 ();
 FILLCELL_X32 FILLER_286_1359 ();
 FILLCELL_X32 FILLER_286_1391 ();
 FILLCELL_X32 FILLER_286_1423 ();
 FILLCELL_X32 FILLER_286_1455 ();
 FILLCELL_X32 FILLER_286_1487 ();
 FILLCELL_X32 FILLER_286_1519 ();
 FILLCELL_X32 FILLER_286_1551 ();
 FILLCELL_X32 FILLER_286_1583 ();
 FILLCELL_X32 FILLER_286_1615 ();
 FILLCELL_X32 FILLER_286_1647 ();
 FILLCELL_X32 FILLER_286_1679 ();
 FILLCELL_X32 FILLER_286_1711 ();
 FILLCELL_X32 FILLER_286_1743 ();
 FILLCELL_X32 FILLER_286_1775 ();
 FILLCELL_X32 FILLER_286_1807 ();
 FILLCELL_X32 FILLER_286_1839 ();
 FILLCELL_X16 FILLER_286_1871 ();
 FILLCELL_X4 FILLER_286_1887 ();
 FILLCELL_X2 FILLER_286_1891 ();
 FILLCELL_X32 FILLER_286_1894 ();
 FILLCELL_X32 FILLER_286_1926 ();
 FILLCELL_X32 FILLER_286_1958 ();
 FILLCELL_X32 FILLER_286_1990 ();
 FILLCELL_X32 FILLER_286_2022 ();
 FILLCELL_X32 FILLER_286_2054 ();
 FILLCELL_X16 FILLER_286_2086 ();
 FILLCELL_X8 FILLER_286_2102 ();
 FILLCELL_X4 FILLER_286_2110 ();
 FILLCELL_X1 FILLER_286_2114 ();
endmodule
