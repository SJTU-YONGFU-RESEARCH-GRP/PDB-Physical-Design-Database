module circular_buffer_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    peek_en,
    rd_en,
    rst_n,
    wr_en,
    fifo_count,
    peek_addr,
    peek_data,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input peek_en;
 input rd_en;
 input rst_n;
 input wr_en;
 output [4:0] fifo_count;
 input [3:0] peek_addr;
 output [7:0] peek_data;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 CLKBUF_X2 _0826_ (.A(net9),
    .Z(_0392_));
 INV_X1 _0827_ (.A(_0392_),
    .ZN(_0812_));
 BUF_X4 _0828_ (.A(_0800_),
    .Z(_0393_));
 INV_X1 _0829_ (.A(_0393_),
    .ZN(_0394_));
 AND2_X1 _0830_ (.A1(_0805_),
    .A2(_0802_),
    .ZN(_0395_));
 INV_X1 _0831_ (.A(_0824_),
    .ZN(_0792_));
 AOI221_X2 _0832_ (.A(_0804_),
    .B1(_0395_),
    .B2(_0792_),
    .C1(_0801_),
    .C2(_0805_),
    .ZN(_0396_));
 XNOR2_X1 _0833_ (.A(_0394_),
    .B(_0396_),
    .ZN(_0397_));
 INV_X1 _0834_ (.A(_0397_),
    .ZN(net11));
 XNOR2_X2 _0835_ (.A(_0805_),
    .B(_0793_),
    .ZN(_0398_));
 INV_X1 _0836_ (.A(_0398_),
    .ZN(net10));
 CLKBUF_X2 _0837_ (.A(_0825_),
    .Z(_0399_));
 INV_X1 _0838_ (.A(_0399_),
    .ZN(net8));
 AND2_X1 _0839_ (.A1(_0393_),
    .A2(_0805_),
    .ZN(_0400_));
 AOI221_X2 _0840_ (.A(_0799_),
    .B1(_0804_),
    .B2(_0393_),
    .C1(_0400_),
    .C2(_0793_),
    .ZN(_0401_));
 XNOR2_X1 _0841_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .ZN(_0402_));
 XOR2_X2 _0842_ (.A(_0401_),
    .B(_0402_),
    .Z(_0403_));
 INV_X2 _0843_ (.A(_0403_),
    .ZN(_0404_));
 BUF_X4 _0844_ (.A(_0404_),
    .Z(_0405_));
 CLKBUF_X3 _0845_ (.A(_0405_),
    .Z(net12));
 BUF_X4 _0846_ (.A(net30),
    .Z(_0406_));
 CLKBUF_X3 _0847_ (.A(_0406_),
    .Z(_0407_));
 NAND4_X1 _0848_ (.A1(_0393_),
    .A2(_0399_),
    .A3(_0812_),
    .A4(_0398_),
    .ZN(_0408_));
 NAND4_X1 _0849_ (.A1(_0394_),
    .A2(_0399_),
    .A3(_0812_),
    .A4(_0398_),
    .ZN(_0409_));
 MUX2_X1 _0850_ (.A(_0408_),
    .B(_0409_),
    .S(_0396_),
    .Z(_0410_));
 BUF_X4 _0851_ (.A(_0410_),
    .Z(_0411_));
 BUF_X8 _0852_ (.A(_0411_),
    .Z(_0412_));
 BUF_X4 _0853_ (.A(_0412_),
    .Z(_0413_));
 NOR2_X1 _0854_ (.A1(_0407_),
    .A2(_0413_),
    .ZN(net13));
 NOR2_X1 _0855_ (.A1(net12),
    .A2(_0413_),
    .ZN(net7));
 INV_X1 _0856_ (.A(net2),
    .ZN(_0794_));
 INV_X1 _0857_ (.A(_0806_),
    .ZN(_0795_));
 BUF_X1 _0858_ (.A(wr_data[0]),
    .Z(_0414_));
 BUF_X2 _0859_ (.A(_0414_),
    .Z(_0415_));
 INV_X1 _0860_ (.A(\wr_ptr[3] ),
    .ZN(_0416_));
 INV_X1 _0861_ (.A(\wr_ptr[2] ),
    .ZN(_0417_));
 NAND2_X1 _0862_ (.A1(_0416_),
    .A2(_0417_),
    .ZN(_0418_));
 CLKBUF_X3 _0863_ (.A(wr_en),
    .Z(_0419_));
 NAND2_X1 _0864_ (.A1(_0419_),
    .A2(_0817_),
    .ZN(_0420_));
 NOR2_X1 _0865_ (.A1(_0418_),
    .A2(_0420_),
    .ZN(_0421_));
 OAI21_X4 _0866_ (.A(_0421_),
    .B1(_0412_),
    .B2(_0406_),
    .ZN(_0422_));
 MUX2_X1 _0867_ (.A(_0415_),
    .B(\mem[0][0] ),
    .S(_0422_),
    .Z(_0116_));
 CLKBUF_X2 _0868_ (.A(wr_data[1]),
    .Z(_0423_));
 BUF_X2 _0869_ (.A(_0423_),
    .Z(_0424_));
 MUX2_X1 _0870_ (.A(_0424_),
    .B(\mem[0][1] ),
    .S(_0422_),
    .Z(_0117_));
 CLKBUF_X2 _0871_ (.A(wr_data[2]),
    .Z(_0425_));
 BUF_X2 _0872_ (.A(_0425_),
    .Z(_0426_));
 MUX2_X1 _0873_ (.A(_0426_),
    .B(\mem[0][2] ),
    .S(_0422_),
    .Z(_0118_));
 CLKBUF_X2 _0874_ (.A(wr_data[3]),
    .Z(_0427_));
 BUF_X2 _0875_ (.A(_0427_),
    .Z(_0428_));
 MUX2_X1 _0876_ (.A(_0428_),
    .B(\mem[0][3] ),
    .S(_0422_),
    .Z(_0119_));
 CLKBUF_X2 _0877_ (.A(wr_data[4]),
    .Z(_0429_));
 BUF_X2 _0878_ (.A(_0429_),
    .Z(_0430_));
 MUX2_X1 _0879_ (.A(_0430_),
    .B(\mem[0][4] ),
    .S(_0422_),
    .Z(_0120_));
 BUF_X2 _0880_ (.A(wr_data[5]),
    .Z(_0431_));
 BUF_X2 _0881_ (.A(_0431_),
    .Z(_0432_));
 MUX2_X1 _0882_ (.A(_0432_),
    .B(\mem[0][5] ),
    .S(_0422_),
    .Z(_0121_));
 CLKBUF_X2 _0883_ (.A(wr_data[6]),
    .Z(_0433_));
 BUF_X2 _0884_ (.A(_0433_),
    .Z(_0434_));
 MUX2_X1 _0885_ (.A(_0434_),
    .B(\mem[0][6] ),
    .S(_0422_),
    .Z(_0122_));
 CLKBUF_X2 _0886_ (.A(wr_data[7]),
    .Z(_0435_));
 BUF_X2 _0887_ (.A(_0435_),
    .Z(_0436_));
 MUX2_X1 _0888_ (.A(_0436_),
    .B(\mem[0][7] ),
    .S(_0422_),
    .Z(_0123_));
 NAND2_X1 _0889_ (.A1(\wr_ptr[3] ),
    .A2(_0417_),
    .ZN(_0437_));
 NAND2_X1 _0890_ (.A1(_0419_),
    .A2(_0818_),
    .ZN(_0438_));
 NOR2_X1 _0891_ (.A1(_0437_),
    .A2(_0438_),
    .ZN(_0439_));
 OAI21_X4 _0892_ (.A(_0439_),
    .B1(_0412_),
    .B2(_0406_),
    .ZN(_0440_));
 MUX2_X1 _0893_ (.A(_0415_),
    .B(\mem[10][0] ),
    .S(_0440_),
    .Z(_0124_));
 MUX2_X1 _0894_ (.A(_0424_),
    .B(\mem[10][1] ),
    .S(_0440_),
    .Z(_0125_));
 MUX2_X1 _0895_ (.A(_0426_),
    .B(\mem[10][2] ),
    .S(_0440_),
    .Z(_0126_));
 MUX2_X1 _0896_ (.A(_0428_),
    .B(\mem[10][3] ),
    .S(_0440_),
    .Z(_0127_));
 MUX2_X1 _0897_ (.A(_0430_),
    .B(\mem[10][4] ),
    .S(_0440_),
    .Z(_0128_));
 MUX2_X1 _0898_ (.A(_0432_),
    .B(\mem[10][5] ),
    .S(_0440_),
    .Z(_0129_));
 MUX2_X1 _0899_ (.A(_0434_),
    .B(\mem[10][6] ),
    .S(_0440_),
    .Z(_0130_));
 MUX2_X1 _0900_ (.A(_0436_),
    .B(\mem[10][7] ),
    .S(_0440_),
    .Z(_0131_));
 NAND2_X1 _0901_ (.A1(_0419_),
    .A2(_0822_),
    .ZN(_0441_));
 NOR2_X1 _0902_ (.A1(_0437_),
    .A2(_0441_),
    .ZN(_0442_));
 OAI21_X4 _0903_ (.A(_0442_),
    .B1(_0412_),
    .B2(_0406_),
    .ZN(_0443_));
 MUX2_X1 _0904_ (.A(_0415_),
    .B(\mem[11][0] ),
    .S(_0443_),
    .Z(_0132_));
 MUX2_X1 _0905_ (.A(_0424_),
    .B(\mem[11][1] ),
    .S(_0443_),
    .Z(_0133_));
 MUX2_X1 _0906_ (.A(_0426_),
    .B(\mem[11][2] ),
    .S(_0443_),
    .Z(_0134_));
 MUX2_X1 _0907_ (.A(_0428_),
    .B(\mem[11][3] ),
    .S(_0443_),
    .Z(_0135_));
 MUX2_X1 _0908_ (.A(_0430_),
    .B(\mem[11][4] ),
    .S(_0443_),
    .Z(_0136_));
 MUX2_X1 _0909_ (.A(_0432_),
    .B(\mem[11][5] ),
    .S(_0443_),
    .Z(_0137_));
 MUX2_X1 _0910_ (.A(_0434_),
    .B(\mem[11][6] ),
    .S(_0443_),
    .Z(_0138_));
 MUX2_X1 _0911_ (.A(_0436_),
    .B(\mem[11][7] ),
    .S(_0443_),
    .Z(_0139_));
 NOR2_X2 _0912_ (.A1(_0416_),
    .A2(_0417_),
    .ZN(_0444_));
 NAND3_X2 _0913_ (.A1(_0419_),
    .A2(_0817_),
    .A3(_0444_),
    .ZN(_0445_));
 NOR4_X1 _0914_ (.A1(_0394_),
    .A2(net8),
    .A3(_0392_),
    .A4(net10),
    .ZN(_0446_));
 NOR4_X1 _0915_ (.A1(_0393_),
    .A2(net8),
    .A3(_0392_),
    .A4(net10),
    .ZN(_0447_));
 MUX2_X1 _0916_ (.A(_0446_),
    .B(_0447_),
    .S(_0396_),
    .Z(_0448_));
 BUF_X4 _0917_ (.A(_0448_),
    .Z(_0449_));
 AOI21_X4 _0918_ (.A(_0445_),
    .B1(_0449_),
    .B2(_0405_),
    .ZN(_0450_));
 MUX2_X1 _0919_ (.A(\mem[12][0] ),
    .B(_0415_),
    .S(_0450_),
    .Z(_0140_));
 MUX2_X1 _0920_ (.A(\mem[12][1] ),
    .B(_0424_),
    .S(_0450_),
    .Z(_0141_));
 MUX2_X1 _0921_ (.A(\mem[12][2] ),
    .B(_0426_),
    .S(_0450_),
    .Z(_0142_));
 MUX2_X1 _0922_ (.A(\mem[12][3] ),
    .B(_0428_),
    .S(_0450_),
    .Z(_0143_));
 MUX2_X1 _0923_ (.A(\mem[12][4] ),
    .B(_0430_),
    .S(_0450_),
    .Z(_0144_));
 MUX2_X1 _0924_ (.A(\mem[12][5] ),
    .B(_0432_),
    .S(_0450_),
    .Z(_0145_));
 MUX2_X1 _0925_ (.A(\mem[12][6] ),
    .B(_0434_),
    .S(_0450_),
    .Z(_0146_));
 MUX2_X1 _0926_ (.A(\mem[12][7] ),
    .B(_0436_),
    .S(_0450_),
    .Z(_0147_));
 NAND3_X2 _0927_ (.A1(_0419_),
    .A2(_0820_),
    .A3(_0444_),
    .ZN(_0451_));
 AOI21_X4 _0928_ (.A(_0451_),
    .B1(_0449_),
    .B2(_0405_),
    .ZN(_0452_));
 MUX2_X1 _0929_ (.A(\mem[13][0] ),
    .B(_0415_),
    .S(_0452_),
    .Z(_0148_));
 MUX2_X1 _0930_ (.A(\mem[13][1] ),
    .B(_0424_),
    .S(_0452_),
    .Z(_0149_));
 MUX2_X1 _0931_ (.A(\mem[13][2] ),
    .B(_0426_),
    .S(_0452_),
    .Z(_0150_));
 MUX2_X1 _0932_ (.A(\mem[13][3] ),
    .B(_0428_),
    .S(_0452_),
    .Z(_0151_));
 MUX2_X1 _0933_ (.A(\mem[13][4] ),
    .B(_0430_),
    .S(_0452_),
    .Z(_0152_));
 MUX2_X1 _0934_ (.A(\mem[13][5] ),
    .B(_0432_),
    .S(_0452_),
    .Z(_0153_));
 MUX2_X1 _0935_ (.A(\mem[13][6] ),
    .B(_0434_),
    .S(_0452_),
    .Z(_0154_));
 MUX2_X1 _0936_ (.A(\mem[13][7] ),
    .B(_0436_),
    .S(_0452_),
    .Z(_0155_));
 NAND3_X2 _0937_ (.A1(_0419_),
    .A2(_0818_),
    .A3(_0444_),
    .ZN(_0453_));
 AOI21_X4 _0938_ (.A(_0453_),
    .B1(_0449_),
    .B2(_0405_),
    .ZN(_0454_));
 MUX2_X1 _0939_ (.A(\mem[14][0] ),
    .B(_0415_),
    .S(_0454_),
    .Z(_0156_));
 MUX2_X1 _0940_ (.A(\mem[14][1] ),
    .B(_0424_),
    .S(_0454_),
    .Z(_0157_));
 MUX2_X1 _0941_ (.A(\mem[14][2] ),
    .B(_0426_),
    .S(_0454_),
    .Z(_0158_));
 MUX2_X1 _0942_ (.A(\mem[14][3] ),
    .B(_0428_),
    .S(_0454_),
    .Z(_0159_));
 MUX2_X1 _0943_ (.A(\mem[14][4] ),
    .B(_0430_),
    .S(_0454_),
    .Z(_0160_));
 MUX2_X1 _0944_ (.A(\mem[14][5] ),
    .B(_0432_),
    .S(_0454_),
    .Z(_0161_));
 MUX2_X1 _0945_ (.A(\mem[14][6] ),
    .B(_0434_),
    .S(_0454_),
    .Z(_0162_));
 MUX2_X1 _0946_ (.A(\mem[14][7] ),
    .B(_0436_),
    .S(_0454_),
    .Z(_0163_));
 NAND3_X1 _0947_ (.A1(_0419_),
    .A2(_0822_),
    .A3(_0444_),
    .ZN(_0455_));
 AOI21_X4 _0948_ (.A(_0455_),
    .B1(_0449_),
    .B2(_0405_),
    .ZN(_0456_));
 MUX2_X1 _0949_ (.A(\mem[15][0] ),
    .B(_0415_),
    .S(_0456_),
    .Z(_0164_));
 MUX2_X1 _0950_ (.A(\mem[15][1] ),
    .B(_0424_),
    .S(_0456_),
    .Z(_0165_));
 MUX2_X1 _0951_ (.A(\mem[15][2] ),
    .B(_0426_),
    .S(_0456_),
    .Z(_0166_));
 MUX2_X1 _0952_ (.A(\mem[15][3] ),
    .B(_0428_),
    .S(_0456_),
    .Z(_0167_));
 MUX2_X1 _0953_ (.A(\mem[15][4] ),
    .B(_0430_),
    .S(_0456_),
    .Z(_0168_));
 MUX2_X1 _0954_ (.A(\mem[15][5] ),
    .B(_0432_),
    .S(_0456_),
    .Z(_0169_));
 MUX2_X1 _0955_ (.A(\mem[15][6] ),
    .B(_0434_),
    .S(_0456_),
    .Z(_0170_));
 MUX2_X1 _0956_ (.A(\mem[15][7] ),
    .B(_0436_),
    .S(_0456_),
    .Z(_0171_));
 NAND2_X1 _0957_ (.A1(_0419_),
    .A2(_0820_),
    .ZN(_0457_));
 NOR2_X1 _0958_ (.A1(_0418_),
    .A2(_0457_),
    .ZN(_0458_));
 OAI21_X4 _0959_ (.A(_0458_),
    .B1(_0412_),
    .B2(_0406_),
    .ZN(_0459_));
 MUX2_X1 _0960_ (.A(_0415_),
    .B(\mem[1][0] ),
    .S(_0459_),
    .Z(_0172_));
 MUX2_X1 _0961_ (.A(_0424_),
    .B(\mem[1][1] ),
    .S(_0459_),
    .Z(_0173_));
 MUX2_X1 _0962_ (.A(_0426_),
    .B(\mem[1][2] ),
    .S(_0459_),
    .Z(_0174_));
 MUX2_X1 _0963_ (.A(_0428_),
    .B(\mem[1][3] ),
    .S(_0459_),
    .Z(_0175_));
 MUX2_X1 _0964_ (.A(_0430_),
    .B(\mem[1][4] ),
    .S(_0459_),
    .Z(_0176_));
 MUX2_X1 _0965_ (.A(_0432_),
    .B(\mem[1][5] ),
    .S(_0459_),
    .Z(_0177_));
 MUX2_X1 _0966_ (.A(_0434_),
    .B(\mem[1][6] ),
    .S(_0459_),
    .Z(_0178_));
 MUX2_X1 _0967_ (.A(_0436_),
    .B(\mem[1][7] ),
    .S(_0459_),
    .Z(_0179_));
 NOR2_X1 _0968_ (.A1(_0418_),
    .A2(_0438_),
    .ZN(_0460_));
 OAI21_X4 _0969_ (.A(_0460_),
    .B1(_0412_),
    .B2(_0406_),
    .ZN(_0461_));
 MUX2_X1 _0970_ (.A(_0415_),
    .B(\mem[2][0] ),
    .S(_0461_),
    .Z(_0180_));
 MUX2_X1 _0971_ (.A(_0424_),
    .B(\mem[2][1] ),
    .S(_0461_),
    .Z(_0181_));
 MUX2_X1 _0972_ (.A(_0426_),
    .B(\mem[2][2] ),
    .S(_0461_),
    .Z(_0182_));
 MUX2_X1 _0973_ (.A(_0428_),
    .B(\mem[2][3] ),
    .S(_0461_),
    .Z(_0183_));
 MUX2_X1 _0974_ (.A(_0430_),
    .B(\mem[2][4] ),
    .S(_0461_),
    .Z(_0184_));
 MUX2_X1 _0975_ (.A(_0432_),
    .B(\mem[2][5] ),
    .S(_0461_),
    .Z(_0185_));
 MUX2_X1 _0976_ (.A(_0434_),
    .B(\mem[2][6] ),
    .S(_0461_),
    .Z(_0186_));
 MUX2_X1 _0977_ (.A(_0436_),
    .B(\mem[2][7] ),
    .S(_0461_),
    .Z(_0187_));
 NOR2_X1 _0978_ (.A1(_0418_),
    .A2(_0441_),
    .ZN(_0462_));
 OAI21_X4 _0979_ (.A(_0462_),
    .B1(_0412_),
    .B2(net30),
    .ZN(_0463_));
 MUX2_X1 _0980_ (.A(_0415_),
    .B(\mem[3][0] ),
    .S(_0463_),
    .Z(_0188_));
 MUX2_X1 _0981_ (.A(_0424_),
    .B(\mem[3][1] ),
    .S(_0463_),
    .Z(_0189_));
 MUX2_X1 _0982_ (.A(_0426_),
    .B(\mem[3][2] ),
    .S(_0463_),
    .Z(_0190_));
 MUX2_X1 _0983_ (.A(_0428_),
    .B(\mem[3][3] ),
    .S(_0463_),
    .Z(_0191_));
 MUX2_X1 _0984_ (.A(_0430_),
    .B(\mem[3][4] ),
    .S(_0463_),
    .Z(_0192_));
 MUX2_X1 _0985_ (.A(_0432_),
    .B(\mem[3][5] ),
    .S(_0463_),
    .Z(_0193_));
 MUX2_X1 _0986_ (.A(_0434_),
    .B(\mem[3][6] ),
    .S(_0463_),
    .Z(_0194_));
 MUX2_X1 _0987_ (.A(_0436_),
    .B(\mem[3][7] ),
    .S(_0463_),
    .Z(_0195_));
 NAND2_X1 _0988_ (.A1(_0416_),
    .A2(\wr_ptr[2] ),
    .ZN(_0464_));
 NOR2_X1 _0989_ (.A1(_0420_),
    .A2(_0464_),
    .ZN(_0465_));
 OAI21_X4 _0990_ (.A(_0465_),
    .B1(_0412_),
    .B2(net30),
    .ZN(_0466_));
 MUX2_X1 _0991_ (.A(_0414_),
    .B(\mem[4][0] ),
    .S(_0466_),
    .Z(_0196_));
 MUX2_X1 _0992_ (.A(_0423_),
    .B(\mem[4][1] ),
    .S(_0466_),
    .Z(_0197_));
 MUX2_X1 _0993_ (.A(_0425_),
    .B(\mem[4][2] ),
    .S(_0466_),
    .Z(_0198_));
 MUX2_X1 _0994_ (.A(_0427_),
    .B(\mem[4][3] ),
    .S(_0466_),
    .Z(_0199_));
 MUX2_X1 _0995_ (.A(_0429_),
    .B(\mem[4][4] ),
    .S(_0466_),
    .Z(_0200_));
 MUX2_X1 _0996_ (.A(_0431_),
    .B(\mem[4][5] ),
    .S(_0466_),
    .Z(_0201_));
 MUX2_X1 _0997_ (.A(_0433_),
    .B(\mem[4][6] ),
    .S(_0466_),
    .Z(_0202_));
 MUX2_X1 _0998_ (.A(_0435_),
    .B(\mem[4][7] ),
    .S(_0466_),
    .Z(_0203_));
 NOR2_X1 _0999_ (.A1(_0457_),
    .A2(_0464_),
    .ZN(_0467_));
 OAI21_X4 _1000_ (.A(_0467_),
    .B1(_0411_),
    .B2(net30),
    .ZN(_0468_));
 MUX2_X1 _1001_ (.A(_0414_),
    .B(\mem[5][0] ),
    .S(_0468_),
    .Z(_0204_));
 MUX2_X1 _1002_ (.A(_0423_),
    .B(\mem[5][1] ),
    .S(_0468_),
    .Z(_0205_));
 MUX2_X1 _1003_ (.A(_0425_),
    .B(\mem[5][2] ),
    .S(_0468_),
    .Z(_0206_));
 MUX2_X1 _1004_ (.A(_0427_),
    .B(\mem[5][3] ),
    .S(_0468_),
    .Z(_0207_));
 MUX2_X1 _1005_ (.A(_0429_),
    .B(\mem[5][4] ),
    .S(_0468_),
    .Z(_0208_));
 MUX2_X1 _1006_ (.A(_0431_),
    .B(\mem[5][5] ),
    .S(_0468_),
    .Z(_0209_));
 MUX2_X1 _1007_ (.A(_0433_),
    .B(\mem[5][6] ),
    .S(_0468_),
    .Z(_0210_));
 MUX2_X1 _1008_ (.A(_0435_),
    .B(\mem[5][7] ),
    .S(_0468_),
    .Z(_0211_));
 NOR2_X1 _1009_ (.A1(_0438_),
    .A2(_0464_),
    .ZN(_0469_));
 OAI21_X4 _1010_ (.A(_0469_),
    .B1(_0411_),
    .B2(net30),
    .ZN(_0470_));
 MUX2_X1 _1011_ (.A(_0414_),
    .B(\mem[6][0] ),
    .S(_0470_),
    .Z(_0212_));
 MUX2_X1 _1012_ (.A(_0423_),
    .B(\mem[6][1] ),
    .S(_0470_),
    .Z(_0213_));
 MUX2_X1 _1013_ (.A(_0425_),
    .B(\mem[6][2] ),
    .S(_0470_),
    .Z(_0214_));
 MUX2_X1 _1014_ (.A(_0427_),
    .B(\mem[6][3] ),
    .S(_0470_),
    .Z(_0215_));
 MUX2_X1 _1015_ (.A(_0429_),
    .B(\mem[6][4] ),
    .S(_0470_),
    .Z(_0216_));
 MUX2_X1 _1016_ (.A(_0431_),
    .B(\mem[6][5] ),
    .S(_0470_),
    .Z(_0217_));
 MUX2_X1 _1017_ (.A(_0433_),
    .B(\mem[6][6] ),
    .S(_0470_),
    .Z(_0218_));
 MUX2_X1 _1018_ (.A(_0435_),
    .B(\mem[6][7] ),
    .S(_0470_),
    .Z(_0219_));
 NOR2_X1 _1019_ (.A1(_0441_),
    .A2(_0464_),
    .ZN(_0471_));
 OAI21_X4 _1020_ (.A(_0471_),
    .B1(_0411_),
    .B2(net30),
    .ZN(_0472_));
 MUX2_X1 _1021_ (.A(_0414_),
    .B(\mem[7][0] ),
    .S(_0472_),
    .Z(_0220_));
 MUX2_X1 _1022_ (.A(_0423_),
    .B(\mem[7][1] ),
    .S(_0472_),
    .Z(_0221_));
 MUX2_X1 _1023_ (.A(_0425_),
    .B(\mem[7][2] ),
    .S(_0472_),
    .Z(_0222_));
 MUX2_X1 _1024_ (.A(_0427_),
    .B(\mem[7][3] ),
    .S(_0472_),
    .Z(_0223_));
 MUX2_X1 _1025_ (.A(_0429_),
    .B(\mem[7][4] ),
    .S(_0472_),
    .Z(_0224_));
 MUX2_X1 _1026_ (.A(_0431_),
    .B(\mem[7][5] ),
    .S(_0472_),
    .Z(_0225_));
 MUX2_X1 _1027_ (.A(_0433_),
    .B(\mem[7][6] ),
    .S(_0472_),
    .Z(_0226_));
 MUX2_X1 _1028_ (.A(_0435_),
    .B(\mem[7][7] ),
    .S(_0472_),
    .Z(_0227_));
 NOR2_X1 _1029_ (.A1(_0420_),
    .A2(_0437_),
    .ZN(_0473_));
 OAI21_X4 _1030_ (.A(_0473_),
    .B1(_0411_),
    .B2(net30),
    .ZN(_0474_));
 MUX2_X1 _1031_ (.A(_0414_),
    .B(\mem[8][0] ),
    .S(_0474_),
    .Z(_0228_));
 MUX2_X1 _1032_ (.A(_0423_),
    .B(\mem[8][1] ),
    .S(_0474_),
    .Z(_0229_));
 MUX2_X1 _1033_ (.A(_0425_),
    .B(\mem[8][2] ),
    .S(_0474_),
    .Z(_0230_));
 MUX2_X1 _1034_ (.A(_0427_),
    .B(\mem[8][3] ),
    .S(_0474_),
    .Z(_0231_));
 MUX2_X1 _1035_ (.A(_0429_),
    .B(\mem[8][4] ),
    .S(_0474_),
    .Z(_0232_));
 MUX2_X1 _1036_ (.A(_0431_),
    .B(\mem[8][5] ),
    .S(_0474_),
    .Z(_0233_));
 MUX2_X1 _1037_ (.A(_0433_),
    .B(\mem[8][6] ),
    .S(_0474_),
    .Z(_0234_));
 MUX2_X1 _1038_ (.A(_0435_),
    .B(\mem[8][7] ),
    .S(_0474_),
    .Z(_0235_));
 NOR2_X1 _1039_ (.A1(_0437_),
    .A2(_0457_),
    .ZN(_0475_));
 OAI21_X4 _1040_ (.A(_0475_),
    .B1(_0411_),
    .B2(net30),
    .ZN(_0476_));
 MUX2_X1 _1041_ (.A(_0414_),
    .B(\mem[9][0] ),
    .S(_0476_),
    .Z(_0236_));
 MUX2_X1 _1042_ (.A(_0423_),
    .B(\mem[9][1] ),
    .S(_0476_),
    .Z(_0237_));
 MUX2_X1 _1043_ (.A(_0425_),
    .B(\mem[9][2] ),
    .S(_0476_),
    .Z(_0238_));
 MUX2_X1 _1044_ (.A(_0427_),
    .B(\mem[9][3] ),
    .S(_0476_),
    .Z(_0239_));
 MUX2_X1 _1045_ (.A(_0429_),
    .B(\mem[9][4] ),
    .S(_0476_),
    .Z(_0240_));
 MUX2_X1 _1046_ (.A(_0431_),
    .B(\mem[9][5] ),
    .S(_0476_),
    .Z(_0241_));
 MUX2_X1 _1047_ (.A(_0433_),
    .B(\mem[9][6] ),
    .S(_0476_),
    .Z(_0242_));
 MUX2_X1 _1048_ (.A(_0435_),
    .B(\mem[9][7] ),
    .S(_0476_),
    .Z(_0243_));
 CLKBUF_X2 _1049_ (.A(rd_en),
    .Z(_0477_));
 INV_X2 _1050_ (.A(_0477_),
    .ZN(_0478_));
 BUF_X2 _1051_ (.A(rst_n),
    .Z(_0479_));
 INV_X2 _1052_ (.A(_0479_),
    .ZN(_0480_));
 NOR2_X4 _1053_ (.A1(_0478_),
    .A2(_0480_),
    .ZN(_0481_));
 BUF_X2 _1054_ (.A(\rd_ptr[0] ),
    .Z(_0482_));
 CLKBUF_X3 _1055_ (.A(_0482_),
    .Z(_0483_));
 CLKBUF_X2 _1056_ (.A(\rd_ptr[1] ),
    .Z(_0484_));
 BUF_X4 _1057_ (.A(_0484_),
    .Z(_0485_));
 CLKBUF_X3 _1058_ (.A(_0485_),
    .Z(_0486_));
 MUX2_X1 _1059_ (.A(\mem[8][0] ),
    .B(\mem[10][0] ),
    .S(_0486_),
    .Z(_0487_));
 NOR2_X1 _1060_ (.A1(_0483_),
    .A2(_0487_),
    .ZN(_0488_));
 INV_X2 _1061_ (.A(_0482_),
    .ZN(_0489_));
 CLKBUF_X3 _1062_ (.A(_0489_),
    .Z(_0490_));
 MUX2_X1 _1063_ (.A(\mem[9][0] ),
    .B(\mem[11][0] ),
    .S(_0486_),
    .Z(_0491_));
 NOR2_X1 _1064_ (.A1(_0490_),
    .A2(_0491_),
    .ZN(_0492_));
 BUF_X2 _1065_ (.A(\rd_ptr[3] ),
    .Z(_0493_));
 BUF_X2 _1066_ (.A(\rd_ptr[2] ),
    .Z(_0494_));
 INV_X1 _1067_ (.A(_0494_),
    .ZN(_0495_));
 NAND2_X2 _1068_ (.A1(_0493_),
    .A2(_0495_),
    .ZN(_0496_));
 NAND2_X2 _1069_ (.A1(_0493_),
    .A2(_0494_),
    .ZN(_0497_));
 BUF_X4 _1070_ (.A(_0484_),
    .Z(_0498_));
 MUX2_X1 _1071_ (.A(\mem[12][0] ),
    .B(\mem[14][0] ),
    .S(_0498_),
    .Z(_0499_));
 NOR2_X1 _1072_ (.A1(_0482_),
    .A2(_0499_),
    .ZN(_0500_));
 CLKBUF_X3 _1073_ (.A(_0489_),
    .Z(_0501_));
 BUF_X4 _1074_ (.A(_0484_),
    .Z(_0502_));
 MUX2_X1 _1075_ (.A(\mem[13][0] ),
    .B(\mem[15][0] ),
    .S(_0502_),
    .Z(_0503_));
 NOR2_X1 _1076_ (.A1(_0501_),
    .A2(_0503_),
    .ZN(_0504_));
 OAI33_X1 _1077_ (.A1(_0488_),
    .A2(_0492_),
    .A3(_0496_),
    .B1(_0497_),
    .B2(_0500_),
    .B3(_0504_),
    .ZN(_0505_));
 MUX2_X1 _1078_ (.A(\mem[0][0] ),
    .B(\mem[2][0] ),
    .S(_0486_),
    .Z(_0506_));
 NOR2_X1 _1079_ (.A1(_0483_),
    .A2(_0506_),
    .ZN(_0507_));
 CLKBUF_X3 _1080_ (.A(_0485_),
    .Z(_0508_));
 MUX2_X1 _1081_ (.A(\mem[1][0] ),
    .B(\mem[3][0] ),
    .S(_0508_),
    .Z(_0509_));
 NOR2_X1 _1082_ (.A1(_0490_),
    .A2(_0509_),
    .ZN(_0510_));
 INV_X1 _1083_ (.A(_0493_),
    .ZN(_0511_));
 NAND2_X2 _1084_ (.A1(_0511_),
    .A2(_0495_),
    .ZN(_0512_));
 NAND2_X2 _1085_ (.A1(_0511_),
    .A2(_0494_),
    .ZN(_0513_));
 MUX2_X1 _1086_ (.A(\mem[4][0] ),
    .B(\mem[6][0] ),
    .S(_0502_),
    .Z(_0514_));
 NOR2_X1 _1087_ (.A1(_0482_),
    .A2(_0514_),
    .ZN(_0515_));
 MUX2_X1 _1088_ (.A(\mem[5][0] ),
    .B(\mem[7][0] ),
    .S(_0485_),
    .Z(_0516_));
 NOR2_X1 _1089_ (.A1(_0489_),
    .A2(_0516_),
    .ZN(_0517_));
 OAI33_X1 _1090_ (.A1(_0507_),
    .A2(_0510_),
    .A3(_0512_),
    .B1(_0513_),
    .B2(_0515_),
    .B3(_0517_),
    .ZN(_0518_));
 OAI221_X1 _1091_ (.A(_0481_),
    .B1(_0505_),
    .B2(_0518_),
    .C1(net12),
    .C2(_0413_),
    .ZN(_0519_));
 BUF_X2 _1092_ (.A(_0479_),
    .Z(_0520_));
 BUF_X4 _1093_ (.A(_0449_),
    .Z(_0521_));
 NAND4_X1 _1094_ (.A1(net22),
    .A2(_0520_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0522_));
 NAND3_X1 _1095_ (.A1(_0478_),
    .A2(net22),
    .A3(_0520_),
    .ZN(_0523_));
 NAND3_X1 _1096_ (.A1(_0519_),
    .A2(_0522_),
    .A3(_0523_),
    .ZN(_0244_));
 MUX2_X1 _1097_ (.A(\mem[4][1] ),
    .B(\mem[6][1] ),
    .S(_0486_),
    .Z(_0524_));
 NOR2_X1 _1098_ (.A1(_0483_),
    .A2(_0524_),
    .ZN(_0525_));
 MUX2_X1 _1099_ (.A(\mem[5][1] ),
    .B(\mem[7][1] ),
    .S(_0508_),
    .Z(_0526_));
 NOR2_X1 _1100_ (.A1(_0490_),
    .A2(_0526_),
    .ZN(_0527_));
 CLKBUF_X3 _1101_ (.A(_0482_),
    .Z(_0528_));
 CLKBUF_X3 _1102_ (.A(_0485_),
    .Z(_0529_));
 MUX2_X1 _1103_ (.A(\mem[0][1] ),
    .B(\mem[2][1] ),
    .S(_0529_),
    .Z(_0530_));
 NOR2_X1 _1104_ (.A1(_0528_),
    .A2(_0530_),
    .ZN(_0531_));
 CLKBUF_X3 _1105_ (.A(_0489_),
    .Z(_0532_));
 MUX2_X1 _1106_ (.A(\mem[1][1] ),
    .B(\mem[3][1] ),
    .S(_0498_),
    .Z(_0533_));
 NOR2_X1 _1107_ (.A1(_0532_),
    .A2(_0533_),
    .ZN(_0534_));
 OAI33_X1 _1108_ (.A1(_0513_),
    .A2(_0525_),
    .A3(_0527_),
    .B1(_0531_),
    .B2(_0534_),
    .B3(_0512_),
    .ZN(_0535_));
 MUX2_X1 _1109_ (.A(\mem[12][1] ),
    .B(\mem[14][1] ),
    .S(_0529_),
    .Z(_0536_));
 NOR2_X1 _1110_ (.A1(_0528_),
    .A2(_0536_),
    .ZN(_0537_));
 CLKBUF_X3 _1111_ (.A(_0485_),
    .Z(_0538_));
 MUX2_X1 _1112_ (.A(\mem[13][1] ),
    .B(\mem[15][1] ),
    .S(_0538_),
    .Z(_0539_));
 NOR2_X1 _1113_ (.A1(_0532_),
    .A2(_0539_),
    .ZN(_0540_));
 CLKBUF_X3 _1114_ (.A(_0482_),
    .Z(_0541_));
 MUX2_X1 _1115_ (.A(\mem[8][1] ),
    .B(\mem[10][1] ),
    .S(_0498_),
    .Z(_0542_));
 NOR2_X1 _1116_ (.A1(_0541_),
    .A2(_0542_),
    .ZN(_0543_));
 MUX2_X1 _1117_ (.A(\mem[9][1] ),
    .B(\mem[11][1] ),
    .S(_0502_),
    .Z(_0544_));
 NOR2_X1 _1118_ (.A1(_0501_),
    .A2(_0544_),
    .ZN(_0545_));
 OAI33_X1 _1119_ (.A1(_0497_),
    .A2(_0537_),
    .A3(_0540_),
    .B1(_0543_),
    .B2(_0545_),
    .B3(_0496_),
    .ZN(_0546_));
 OAI221_X2 _1120_ (.A(_0481_),
    .B1(_0535_),
    .B2(_0546_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0547_));
 NAND4_X1 _1121_ (.A1(net23),
    .A2(_0520_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0548_));
 NAND3_X1 _1122_ (.A1(_0478_),
    .A2(net23),
    .A3(_0520_),
    .ZN(_0549_));
 NAND3_X1 _1123_ (.A1(_0547_),
    .A2(_0548_),
    .A3(_0549_),
    .ZN(_0245_));
 MUX2_X1 _1124_ (.A(\mem[4][2] ),
    .B(\mem[6][2] ),
    .S(_0486_),
    .Z(_0550_));
 NOR2_X1 _1125_ (.A1(_0483_),
    .A2(_0550_),
    .ZN(_0551_));
 MUX2_X1 _1126_ (.A(\mem[5][2] ),
    .B(\mem[7][2] ),
    .S(_0508_),
    .Z(_0552_));
 NOR2_X1 _1127_ (.A1(_0490_),
    .A2(_0552_),
    .ZN(_0553_));
 MUX2_X1 _1128_ (.A(\mem[0][2] ),
    .B(\mem[2][2] ),
    .S(_0529_),
    .Z(_0554_));
 NOR2_X1 _1129_ (.A1(_0528_),
    .A2(_0554_),
    .ZN(_0555_));
 MUX2_X1 _1130_ (.A(\mem[1][2] ),
    .B(\mem[3][2] ),
    .S(_0502_),
    .Z(_0556_));
 NOR2_X1 _1131_ (.A1(_0532_),
    .A2(_0556_),
    .ZN(_0557_));
 OAI33_X1 _1132_ (.A1(_0513_),
    .A2(_0551_),
    .A3(_0553_),
    .B1(_0555_),
    .B2(_0557_),
    .B3(_0512_),
    .ZN(_0558_));
 MUX2_X1 _1133_ (.A(\mem[12][2] ),
    .B(\mem[14][2] ),
    .S(_0529_),
    .Z(_0559_));
 NOR2_X1 _1134_ (.A1(_0528_),
    .A2(_0559_),
    .ZN(_0560_));
 MUX2_X1 _1135_ (.A(\mem[13][2] ),
    .B(\mem[15][2] ),
    .S(_0538_),
    .Z(_0561_));
 NOR2_X1 _1136_ (.A1(_0532_),
    .A2(_0561_),
    .ZN(_0562_));
 MUX2_X1 _1137_ (.A(\mem[8][2] ),
    .B(\mem[10][2] ),
    .S(_0498_),
    .Z(_0563_));
 NOR2_X1 _1138_ (.A1(_0541_),
    .A2(_0563_),
    .ZN(_0564_));
 MUX2_X1 _1139_ (.A(\mem[9][2] ),
    .B(\mem[11][2] ),
    .S(_0502_),
    .Z(_0565_));
 NOR2_X1 _1140_ (.A1(_0501_),
    .A2(_0565_),
    .ZN(_0566_));
 OAI33_X1 _1141_ (.A1(_0497_),
    .A2(_0560_),
    .A3(_0562_),
    .B1(_0564_),
    .B2(_0566_),
    .B3(_0496_),
    .ZN(_0567_));
 OAI221_X2 _1142_ (.A(_0481_),
    .B1(_0558_),
    .B2(_0567_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0568_));
 BUF_X2 _1143_ (.A(_0479_),
    .Z(_0569_));
 NAND4_X1 _1144_ (.A1(net24),
    .A2(_0569_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0570_));
 NAND3_X1 _1145_ (.A1(_0478_),
    .A2(net24),
    .A3(_0520_),
    .ZN(_0571_));
 NAND3_X1 _1146_ (.A1(_0568_),
    .A2(_0570_),
    .A3(_0571_),
    .ZN(_0246_));
 MUX2_X1 _1147_ (.A(\mem[4][3] ),
    .B(\mem[6][3] ),
    .S(_0486_),
    .Z(_0572_));
 NOR2_X1 _1148_ (.A1(_0483_),
    .A2(_0572_),
    .ZN(_0573_));
 MUX2_X1 _1149_ (.A(\mem[5][3] ),
    .B(\mem[7][3] ),
    .S(_0508_),
    .Z(_0574_));
 NOR2_X1 _1150_ (.A1(_0490_),
    .A2(_0574_),
    .ZN(_0575_));
 MUX2_X1 _1151_ (.A(\mem[0][3] ),
    .B(\mem[2][3] ),
    .S(_0529_),
    .Z(_0576_));
 NOR2_X1 _1152_ (.A1(_0528_),
    .A2(_0576_),
    .ZN(_0577_));
 MUX2_X1 _1153_ (.A(\mem[1][3] ),
    .B(\mem[3][3] ),
    .S(_0502_),
    .Z(_0578_));
 NOR2_X1 _1154_ (.A1(_0532_),
    .A2(_0578_),
    .ZN(_0579_));
 OAI33_X1 _1155_ (.A1(_0513_),
    .A2(_0573_),
    .A3(_0575_),
    .B1(_0577_),
    .B2(_0579_),
    .B3(_0512_),
    .ZN(_0580_));
 MUX2_X1 _1156_ (.A(\mem[12][3] ),
    .B(\mem[14][3] ),
    .S(_0529_),
    .Z(_0581_));
 NOR2_X1 _1157_ (.A1(_0528_),
    .A2(_0581_),
    .ZN(_0582_));
 MUX2_X1 _1158_ (.A(\mem[13][3] ),
    .B(\mem[15][3] ),
    .S(_0538_),
    .Z(_0583_));
 NOR2_X1 _1159_ (.A1(_0532_),
    .A2(_0583_),
    .ZN(_0584_));
 MUX2_X1 _1160_ (.A(\mem[8][3] ),
    .B(\mem[10][3] ),
    .S(_0498_),
    .Z(_0585_));
 NOR2_X1 _1161_ (.A1(_0541_),
    .A2(_0585_),
    .ZN(_0586_));
 MUX2_X1 _1162_ (.A(\mem[9][3] ),
    .B(\mem[11][3] ),
    .S(_0485_),
    .Z(_0587_));
 NOR2_X1 _1163_ (.A1(_0501_),
    .A2(_0587_),
    .ZN(_0588_));
 OAI33_X1 _1164_ (.A1(_0497_),
    .A2(_0582_),
    .A3(_0584_),
    .B1(_0586_),
    .B2(_0588_),
    .B3(_0496_),
    .ZN(_0589_));
 OAI221_X1 _1165_ (.A(_0481_),
    .B1(_0580_),
    .B2(_0589_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0590_));
 NAND4_X1 _1166_ (.A1(net25),
    .A2(_0569_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0591_));
 NAND3_X1 _1167_ (.A1(_0478_),
    .A2(net25),
    .A3(_0520_),
    .ZN(_0592_));
 NAND3_X1 _1168_ (.A1(_0590_),
    .A2(_0591_),
    .A3(_0592_),
    .ZN(_0247_));
 MUX2_X1 _1169_ (.A(\mem[4][4] ),
    .B(\mem[6][4] ),
    .S(_0486_),
    .Z(_0593_));
 NOR2_X1 _1170_ (.A1(_0483_),
    .A2(_0593_),
    .ZN(_0594_));
 MUX2_X1 _1171_ (.A(\mem[5][4] ),
    .B(\mem[7][4] ),
    .S(_0508_),
    .Z(_0595_));
 NOR2_X1 _1172_ (.A1(_0490_),
    .A2(_0595_),
    .ZN(_0596_));
 MUX2_X1 _1173_ (.A(\mem[0][4] ),
    .B(\mem[2][4] ),
    .S(_0538_),
    .Z(_0597_));
 NOR2_X1 _1174_ (.A1(_0541_),
    .A2(_0597_),
    .ZN(_0598_));
 MUX2_X1 _1175_ (.A(\mem[1][4] ),
    .B(\mem[3][4] ),
    .S(_0502_),
    .Z(_0599_));
 NOR2_X1 _1176_ (.A1(_0501_),
    .A2(_0599_),
    .ZN(_0600_));
 OAI33_X1 _1177_ (.A1(_0513_),
    .A2(_0594_),
    .A3(_0596_),
    .B1(_0598_),
    .B2(_0600_),
    .B3(_0512_),
    .ZN(_0601_));
 MUX2_X1 _1178_ (.A(\mem[12][4] ),
    .B(\mem[14][4] ),
    .S(_0529_),
    .Z(_0602_));
 NOR2_X1 _1179_ (.A1(_0528_),
    .A2(_0602_),
    .ZN(_0603_));
 MUX2_X1 _1180_ (.A(\mem[13][4] ),
    .B(\mem[15][4] ),
    .S(_0538_),
    .Z(_0604_));
 NOR2_X1 _1181_ (.A1(_0532_),
    .A2(_0604_),
    .ZN(_0605_));
 MUX2_X1 _1182_ (.A(\mem[8][4] ),
    .B(\mem[10][4] ),
    .S(_0498_),
    .Z(_0606_));
 NOR2_X1 _1183_ (.A1(_0541_),
    .A2(_0606_),
    .ZN(_0607_));
 MUX2_X1 _1184_ (.A(\mem[9][4] ),
    .B(\mem[11][4] ),
    .S(_0485_),
    .Z(_0608_));
 NOR2_X1 _1185_ (.A1(_0501_),
    .A2(_0608_),
    .ZN(_0609_));
 OAI33_X1 _1186_ (.A1(_0497_),
    .A2(_0603_),
    .A3(_0605_),
    .B1(_0607_),
    .B2(_0609_),
    .B3(_0496_),
    .ZN(_0610_));
 OAI221_X1 _1187_ (.A(_0481_),
    .B1(_0601_),
    .B2(_0610_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0611_));
 NAND4_X1 _1188_ (.A1(net26),
    .A2(_0569_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0612_));
 NAND3_X1 _1189_ (.A1(_0478_),
    .A2(net26),
    .A3(_0520_),
    .ZN(_0613_));
 NAND3_X1 _1190_ (.A1(_0611_),
    .A2(_0612_),
    .A3(_0613_),
    .ZN(_0248_));
 MUX2_X1 _1191_ (.A(\mem[4][5] ),
    .B(\mem[6][5] ),
    .S(_0486_),
    .Z(_0614_));
 NOR2_X1 _1192_ (.A1(_0483_),
    .A2(_0614_),
    .ZN(_0615_));
 MUX2_X1 _1193_ (.A(\mem[5][5] ),
    .B(\mem[7][5] ),
    .S(_0508_),
    .Z(_0616_));
 NOR2_X1 _1194_ (.A1(_0490_),
    .A2(_0616_),
    .ZN(_0617_));
 MUX2_X1 _1195_ (.A(\mem[0][5] ),
    .B(\mem[2][5] ),
    .S(_0538_),
    .Z(_0618_));
 NOR2_X1 _1196_ (.A1(_0541_),
    .A2(_0618_),
    .ZN(_0619_));
 MUX2_X1 _1197_ (.A(\mem[1][5] ),
    .B(\mem[3][5] ),
    .S(_0502_),
    .Z(_0620_));
 NOR2_X1 _1198_ (.A1(_0501_),
    .A2(_0620_),
    .ZN(_0621_));
 OAI33_X1 _1199_ (.A1(_0513_),
    .A2(_0615_),
    .A3(_0617_),
    .B1(_0619_),
    .B2(_0621_),
    .B3(_0512_),
    .ZN(_0622_));
 MUX2_X1 _1200_ (.A(\mem[12][5] ),
    .B(\mem[14][5] ),
    .S(_0529_),
    .Z(_0623_));
 NOR2_X1 _1201_ (.A1(_0528_),
    .A2(_0623_),
    .ZN(_0624_));
 MUX2_X1 _1202_ (.A(\mem[13][5] ),
    .B(\mem[15][5] ),
    .S(_0538_),
    .Z(_0625_));
 NOR2_X1 _1203_ (.A1(_0532_),
    .A2(_0625_),
    .ZN(_0626_));
 MUX2_X1 _1204_ (.A(\mem[8][5] ),
    .B(\mem[10][5] ),
    .S(_0498_),
    .Z(_0627_));
 NOR2_X1 _1205_ (.A1(_0541_),
    .A2(_0627_),
    .ZN(_0628_));
 MUX2_X1 _1206_ (.A(\mem[9][5] ),
    .B(\mem[11][5] ),
    .S(_0485_),
    .Z(_0629_));
 NOR2_X1 _1207_ (.A1(_0501_),
    .A2(_0629_),
    .ZN(_0630_));
 OAI33_X1 _1208_ (.A1(_0497_),
    .A2(_0624_),
    .A3(_0626_),
    .B1(_0628_),
    .B2(_0630_),
    .B3(_0496_),
    .ZN(_0631_));
 OAI221_X1 _1209_ (.A(_0481_),
    .B1(_0622_),
    .B2(_0631_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0632_));
 NAND4_X1 _1210_ (.A1(net27),
    .A2(_0569_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0633_));
 NAND3_X1 _1211_ (.A1(_0478_),
    .A2(net27),
    .A3(_0520_),
    .ZN(_0634_));
 NAND3_X1 _1212_ (.A1(_0632_),
    .A2(_0633_),
    .A3(_0634_),
    .ZN(_0249_));
 MUX2_X1 _1213_ (.A(\mem[4][6] ),
    .B(\mem[6][6] ),
    .S(_0508_),
    .Z(_0635_));
 NOR2_X1 _1214_ (.A1(_0483_),
    .A2(_0635_),
    .ZN(_0636_));
 MUX2_X1 _1215_ (.A(\mem[5][6] ),
    .B(\mem[7][6] ),
    .S(_0508_),
    .Z(_0637_));
 NOR2_X1 _1216_ (.A1(_0490_),
    .A2(_0637_),
    .ZN(_0638_));
 MUX2_X1 _1217_ (.A(\mem[0][6] ),
    .B(\mem[2][6] ),
    .S(_0538_),
    .Z(_0639_));
 NOR2_X1 _1218_ (.A1(_0541_),
    .A2(_0639_),
    .ZN(_0640_));
 MUX2_X1 _1219_ (.A(\mem[1][6] ),
    .B(\mem[3][6] ),
    .S(_0502_),
    .Z(_0641_));
 NOR2_X1 _1220_ (.A1(_0501_),
    .A2(_0641_),
    .ZN(_0642_));
 OAI33_X1 _1221_ (.A1(_0513_),
    .A2(_0636_),
    .A3(_0638_),
    .B1(_0640_),
    .B2(_0642_),
    .B3(_0512_),
    .ZN(_0643_));
 MUX2_X1 _1222_ (.A(\mem[12][6] ),
    .B(\mem[14][6] ),
    .S(_0529_),
    .Z(_0644_));
 NOR2_X1 _1223_ (.A1(_0528_),
    .A2(_0644_),
    .ZN(_0645_));
 MUX2_X1 _1224_ (.A(\mem[13][6] ),
    .B(\mem[15][6] ),
    .S(_0538_),
    .Z(_0646_));
 NOR2_X1 _1225_ (.A1(_0532_),
    .A2(_0646_),
    .ZN(_0647_));
 MUX2_X1 _1226_ (.A(\mem[8][6] ),
    .B(\mem[10][6] ),
    .S(_0498_),
    .Z(_0648_));
 NOR2_X1 _1227_ (.A1(_0541_),
    .A2(_0648_),
    .ZN(_0649_));
 MUX2_X1 _1228_ (.A(\mem[9][6] ),
    .B(\mem[11][6] ),
    .S(_0485_),
    .Z(_0650_));
 NOR2_X1 _1229_ (.A1(_0489_),
    .A2(_0650_),
    .ZN(_0651_));
 OAI33_X1 _1230_ (.A1(_0497_),
    .A2(_0645_),
    .A3(_0647_),
    .B1(_0649_),
    .B2(_0651_),
    .B3(_0496_),
    .ZN(_0652_));
 OAI221_X2 _1231_ (.A(_0481_),
    .B1(_0643_),
    .B2(_0652_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0653_));
 NAND4_X1 _1232_ (.A1(net28),
    .A2(_0569_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0654_));
 NAND3_X1 _1233_ (.A1(_0478_),
    .A2(net28),
    .A3(_0520_),
    .ZN(_0655_));
 NAND3_X1 _1234_ (.A1(_0653_),
    .A2(_0654_),
    .A3(_0655_),
    .ZN(_0250_));
 MUX2_X1 _1235_ (.A(\mem[4][7] ),
    .B(\mem[6][7] ),
    .S(_0508_),
    .Z(_0656_));
 NOR2_X1 _1236_ (.A1(_0483_),
    .A2(_0656_),
    .ZN(_0657_));
 MUX2_X1 _1237_ (.A(\mem[5][7] ),
    .B(\mem[7][7] ),
    .S(_0508_),
    .Z(_0658_));
 NOR2_X1 _1238_ (.A1(_0490_),
    .A2(_0658_),
    .ZN(_0659_));
 MUX2_X1 _1239_ (.A(\mem[0][7] ),
    .B(\mem[2][7] ),
    .S(_0538_),
    .Z(_0660_));
 NOR2_X1 _1240_ (.A1(_0541_),
    .A2(_0660_),
    .ZN(_0661_));
 MUX2_X1 _1241_ (.A(\mem[1][7] ),
    .B(\mem[3][7] ),
    .S(_0502_),
    .Z(_0662_));
 NOR2_X1 _1242_ (.A1(_0501_),
    .A2(_0662_),
    .ZN(_0663_));
 OAI33_X1 _1243_ (.A1(_0513_),
    .A2(_0657_),
    .A3(_0659_),
    .B1(_0661_),
    .B2(_0663_),
    .B3(_0512_),
    .ZN(_0664_));
 MUX2_X1 _1244_ (.A(\mem[12][7] ),
    .B(\mem[14][7] ),
    .S(_0529_),
    .Z(_0665_));
 NOR2_X1 _1245_ (.A1(_0528_),
    .A2(_0665_),
    .ZN(_0666_));
 MUX2_X1 _1246_ (.A(\mem[13][7] ),
    .B(\mem[15][7] ),
    .S(_0498_),
    .Z(_0667_));
 NOR2_X1 _1247_ (.A1(_0532_),
    .A2(_0667_),
    .ZN(_0668_));
 MUX2_X1 _1248_ (.A(\mem[8][7] ),
    .B(\mem[10][7] ),
    .S(_0498_),
    .Z(_0669_));
 NOR2_X1 _1249_ (.A1(_0482_),
    .A2(_0669_),
    .ZN(_0670_));
 MUX2_X1 _1250_ (.A(\mem[9][7] ),
    .B(\mem[11][7] ),
    .S(_0485_),
    .Z(_0671_));
 NOR2_X1 _1251_ (.A1(_0489_),
    .A2(_0671_),
    .ZN(_0672_));
 OAI33_X1 _1252_ (.A1(_0497_),
    .A2(_0666_),
    .A3(_0668_),
    .B1(_0670_),
    .B2(_0672_),
    .B3(_0496_),
    .ZN(_0673_));
 OAI221_X2 _1253_ (.A(_0481_),
    .B1(_0664_),
    .B2(_0673_),
    .C1(_0413_),
    .C2(net12),
    .ZN(_0674_));
 NAND4_X1 _1254_ (.A1(net29),
    .A2(_0569_),
    .A3(_0407_),
    .A4(_0521_),
    .ZN(_0675_));
 NAND3_X1 _1255_ (.A1(_0478_),
    .A2(net29),
    .A3(_0520_),
    .ZN(_0676_));
 NAND3_X1 _1256_ (.A1(_0674_),
    .A2(_0675_),
    .A3(_0676_),
    .ZN(_0251_));
 AND2_X1 _1257_ (.A1(_0114_),
    .A2(_0569_),
    .ZN(_0677_));
 CLKBUF_X3 _1258_ (.A(_0480_),
    .Z(_0678_));
 NOR2_X1 _1259_ (.A1(_0490_),
    .A2(_0678_),
    .ZN(_0679_));
 OAI21_X1 _1260_ (.A(_0477_),
    .B1(_0405_),
    .B2(_0412_),
    .ZN(_0680_));
 MUX2_X1 _1261_ (.A(_0677_),
    .B(_0679_),
    .S(_0680_),
    .Z(_0252_));
 AND2_X1 _1262_ (.A1(_0115_),
    .A2(_0479_),
    .ZN(_0681_));
 AND2_X1 _1263_ (.A1(_0486_),
    .A2(_0569_),
    .ZN(_0682_));
 MUX2_X1 _1264_ (.A(_0681_),
    .B(_0682_),
    .S(_0680_),
    .Z(_0253_));
 NOR2_X1 _1265_ (.A1(_0495_),
    .A2(_0678_),
    .ZN(_0683_));
 NOR2_X1 _1266_ (.A1(_0494_),
    .A2(_0678_),
    .ZN(_0684_));
 NAND2_X1 _1267_ (.A1(_0477_),
    .A2(_0815_),
    .ZN(_0685_));
 AOI21_X1 _1268_ (.A(_0685_),
    .B1(_0521_),
    .B2(_0406_),
    .ZN(_0686_));
 MUX2_X1 _1269_ (.A(_0683_),
    .B(_0684_),
    .S(_0686_),
    .Z(_0254_));
 NOR2_X1 _1270_ (.A1(_0511_),
    .A2(_0678_),
    .ZN(_0687_));
 NOR2_X1 _1271_ (.A1(_0493_),
    .A2(_0678_),
    .ZN(_0688_));
 NAND4_X1 _1272_ (.A1(_0477_),
    .A2(_0483_),
    .A3(_0486_),
    .A4(_0494_),
    .ZN(_0689_));
 AOI21_X1 _1273_ (.A(_0689_),
    .B1(_0449_),
    .B2(_0406_),
    .ZN(_0690_));
 MUX2_X1 _1274_ (.A(_0687_),
    .B(_0688_),
    .S(_0690_),
    .Z(_0255_));
 AND2_X1 _1275_ (.A1(\rd_ptr[4] ),
    .A2(_0479_),
    .ZN(_0691_));
 NOR2_X1 _1276_ (.A1(\rd_ptr[4] ),
    .A2(_0678_),
    .ZN(_0692_));
 NAND4_X1 _1277_ (.A1(_0477_),
    .A2(_0493_),
    .A3(_0494_),
    .A4(_0815_),
    .ZN(_0693_));
 AOI21_X1 _1278_ (.A(_0693_),
    .B1(_0449_),
    .B2(_0406_),
    .ZN(_0694_));
 MUX2_X1 _1279_ (.A(_0691_),
    .B(_0692_),
    .S(_0694_),
    .Z(_0256_));
 AND2_X1 _1280_ (.A1(_0112_),
    .A2(_0479_),
    .ZN(_0695_));
 AND2_X1 _1281_ (.A1(\wr_ptr[0] ),
    .A2(_0569_),
    .ZN(_0696_));
 OAI21_X1 _1282_ (.A(_0419_),
    .B1(_0406_),
    .B2(_0412_),
    .ZN(_0697_));
 MUX2_X1 _1283_ (.A(_0695_),
    .B(_0696_),
    .S(_0697_),
    .Z(_0257_));
 AND2_X1 _1284_ (.A1(_0113_),
    .A2(_0479_),
    .ZN(_0698_));
 AND2_X1 _1285_ (.A1(\wr_ptr[1] ),
    .A2(_0569_),
    .ZN(_0699_));
 MUX2_X1 _1286_ (.A(_0698_),
    .B(_0699_),
    .S(_0697_),
    .Z(_0258_));
 NOR2_X1 _1287_ (.A1(_0417_),
    .A2(_0678_),
    .ZN(_0700_));
 NOR2_X1 _1288_ (.A1(\wr_ptr[2] ),
    .A2(_0678_),
    .ZN(_0701_));
 AOI21_X1 _1289_ (.A(_0441_),
    .B1(_0521_),
    .B2(_0405_),
    .ZN(_0702_));
 MUX2_X1 _1290_ (.A(_0700_),
    .B(_0701_),
    .S(_0702_),
    .Z(_0259_));
 NOR2_X1 _1291_ (.A1(_0416_),
    .A2(_0480_),
    .ZN(_0703_));
 NOR2_X1 _1292_ (.A1(\wr_ptr[3] ),
    .A2(_0678_),
    .ZN(_0704_));
 NAND4_X1 _1293_ (.A1(_0419_),
    .A2(\wr_ptr[2] ),
    .A3(\wr_ptr[1] ),
    .A4(\wr_ptr[0] ),
    .ZN(_0705_));
 AOI21_X1 _1294_ (.A(_0705_),
    .B1(_0449_),
    .B2(_0405_),
    .ZN(_0706_));
 MUX2_X1 _1295_ (.A(_0703_),
    .B(_0704_),
    .S(_0706_),
    .Z(_0260_));
 AND2_X1 _1296_ (.A1(\wr_ptr[4] ),
    .A2(_0479_),
    .ZN(_0707_));
 NOR2_X1 _1297_ (.A1(\wr_ptr[4] ),
    .A2(_0678_),
    .ZN(_0708_));
 MUX2_X1 _1298_ (.A(_0707_),
    .B(_0708_),
    .S(_0456_),
    .Z(_0261_));
 XOR2_X1 _1299_ (.A(_0399_),
    .B(_0392_),
    .Z(_0709_));
 NOR4_X1 _1300_ (.A1(net11),
    .A2(net10),
    .A3(_0405_),
    .A4(_0709_),
    .ZN(net5));
 NOR3_X1 _1301_ (.A1(net8),
    .A2(_0392_),
    .A3(net10),
    .ZN(_0710_));
 AOI21_X1 _1302_ (.A(_0405_),
    .B1(net10),
    .B2(_0392_),
    .ZN(_0711_));
 OAI22_X1 _1303_ (.A1(_0407_),
    .A2(_0710_),
    .B1(_0711_),
    .B2(_0397_),
    .ZN(net6));
 INV_X2 _1304_ (.A(net4),
    .ZN(_0712_));
 CLKBUF_X2 _1305_ (.A(peek_addr[3]),
    .Z(_0713_));
 NOR2_X1 _1306_ (.A1(_0393_),
    .A2(_0713_),
    .ZN(_0714_));
 NOR2_X1 _1307_ (.A1(_0394_),
    .A2(_0713_),
    .ZN(_0715_));
 MUX2_X1 _1308_ (.A(_0714_),
    .B(_0715_),
    .S(_0396_),
    .Z(_0716_));
 INV_X1 _1309_ (.A(net3),
    .ZN(_0717_));
 INV_X1 _1310_ (.A(_0813_),
    .ZN(_0718_));
 OAI21_X1 _1311_ (.A(_0814_),
    .B1(net1),
    .B2(_0399_),
    .ZN(_0719_));
 NAND3_X1 _1312_ (.A1(_0717_),
    .A2(_0718_),
    .A3(_0719_),
    .ZN(_0720_));
 AOI21_X1 _1313_ (.A(_0717_),
    .B1(_0718_),
    .B2(_0719_),
    .ZN(_0721_));
 OAI21_X1 _1314_ (.A(_0720_),
    .B1(_0721_),
    .B2(_0398_),
    .ZN(_0722_));
 NAND2_X1 _1315_ (.A1(_0393_),
    .A2(_0713_),
    .ZN(_0723_));
 NAND2_X1 _1316_ (.A1(_0394_),
    .A2(_0713_),
    .ZN(_0724_));
 MUX2_X1 _1317_ (.A(_0723_),
    .B(_0724_),
    .S(_0396_),
    .Z(_0725_));
 AOI211_X4 _1318_ (.A(_0404_),
    .B(_0716_),
    .C1(_0722_),
    .C2(_0725_),
    .ZN(_0726_));
 BUF_X2 _1319_ (.A(_0811_),
    .Z(_0727_));
 XNOR2_X2 _1320_ (.A(_0796_),
    .B(_0727_),
    .ZN(_0728_));
 BUF_X2 _1321_ (.A(_0728_),
    .Z(_0729_));
 BUF_X8 _1322_ (.A(_0797_),
    .Z(_0730_));
 BUF_X4 _1323_ (.A(_0730_),
    .Z(_0731_));
 MUX2_X1 _1324_ (.A(\mem[12][0] ),
    .B(\mem[14][0] ),
    .S(_0731_),
    .Z(_0732_));
 MUX2_X1 _1325_ (.A(\mem[13][0] ),
    .B(\mem[15][0] ),
    .S(_0731_),
    .Z(_0733_));
 BUF_X2 _1326_ (.A(_0807_),
    .Z(_0734_));
 BUF_X4 _1327_ (.A(_0734_),
    .Z(_0735_));
 MUX2_X1 _1328_ (.A(_0732_),
    .B(_0733_),
    .S(_0735_),
    .Z(_0736_));
 NAND2_X1 _1329_ (.A1(_0729_),
    .A2(_0736_),
    .ZN(_0737_));
 MUX2_X1 _1330_ (.A(\mem[4][0] ),
    .B(\mem[6][0] ),
    .S(_0731_),
    .Z(_0738_));
 MUX2_X1 _1331_ (.A(\mem[5][0] ),
    .B(\mem[7][0] ),
    .S(_0731_),
    .Z(_0739_));
 MUX2_X1 _1332_ (.A(_0738_),
    .B(_0739_),
    .S(_0735_),
    .Z(_0740_));
 NAND2_X1 _1333_ (.A1(_0729_),
    .A2(_0740_),
    .ZN(_0741_));
 NAND3_X1 _1334_ (.A1(_0806_),
    .A2(_0809_),
    .A3(_0727_),
    .ZN(_0742_));
 AOI21_X1 _1335_ (.A(_0810_),
    .B1(_0808_),
    .B2(_0727_),
    .ZN(_0743_));
 NAND2_X1 _1336_ (.A1(_0742_),
    .A2(_0743_),
    .ZN(_0744_));
 XOR2_X2 _1337_ (.A(_0713_),
    .B(_0493_),
    .Z(_0745_));
 XNOR2_X2 _1338_ (.A(_0744_),
    .B(_0745_),
    .ZN(_0746_));
 MUX2_X1 _1339_ (.A(_0737_),
    .B(_0741_),
    .S(_0746_),
    .Z(_0747_));
 XOR2_X2 _1340_ (.A(_0796_),
    .B(_0727_),
    .Z(_0748_));
 BUF_X2 _1341_ (.A(_0748_),
    .Z(_0749_));
 MUX2_X1 _1342_ (.A(\mem[8][0] ),
    .B(\mem[10][0] ),
    .S(_0731_),
    .Z(_0750_));
 MUX2_X1 _1343_ (.A(\mem[9][0] ),
    .B(\mem[11][0] ),
    .S(_0731_),
    .Z(_0751_));
 MUX2_X1 _1344_ (.A(_0750_),
    .B(_0751_),
    .S(_0735_),
    .Z(_0752_));
 NAND2_X1 _1345_ (.A1(_0749_),
    .A2(_0752_),
    .ZN(_0753_));
 MUX2_X1 _1346_ (.A(\mem[0][0] ),
    .B(\mem[2][0] ),
    .S(_0731_),
    .Z(_0754_));
 MUX2_X1 _1347_ (.A(\mem[1][0] ),
    .B(\mem[3][0] ),
    .S(_0731_),
    .Z(_0755_));
 MUX2_X1 _1348_ (.A(_0754_),
    .B(_0755_),
    .S(_0735_),
    .Z(_0756_));
 NAND2_X1 _1349_ (.A1(_0749_),
    .A2(_0756_),
    .ZN(_0757_));
 MUX2_X1 _1350_ (.A(_0753_),
    .B(_0757_),
    .S(_0746_),
    .Z(_0758_));
 AOI211_X2 _1351_ (.A(_0712_),
    .B(_0726_),
    .C1(_0747_),
    .C2(_0758_),
    .ZN(net14));
 BUF_X4 _1352_ (.A(_0730_),
    .Z(_0759_));
 MUX2_X1 _1353_ (.A(_0012_),
    .B(_0014_),
    .S(_0759_),
    .Z(_0760_));
 MUX2_X1 _1354_ (.A(_0013_),
    .B(_0015_),
    .S(_0759_),
    .Z(_0761_));
 BUF_X4 _1355_ (.A(_0734_),
    .Z(_0762_));
 MUX2_X1 _1356_ (.A(_0760_),
    .B(_0761_),
    .S(_0762_),
    .Z(_0262_));
 AND2_X1 _1357_ (.A1(_0729_),
    .A2(_0262_),
    .ZN(_0263_));
 BUF_X4 _1358_ (.A(_0730_),
    .Z(_0264_));
 MUX2_X1 _1359_ (.A(_0004_),
    .B(_0006_),
    .S(_0264_),
    .Z(_0265_));
 MUX2_X1 _1360_ (.A(_0005_),
    .B(_0007_),
    .S(_0731_),
    .Z(_0266_));
 MUX2_X1 _1361_ (.A(_0265_),
    .B(_0266_),
    .S(_0735_),
    .Z(_0267_));
 AND2_X1 _1362_ (.A1(_0729_),
    .A2(_0267_),
    .ZN(_0268_));
 CLKBUF_X3 _1363_ (.A(_0746_),
    .Z(_0269_));
 MUX2_X1 _1364_ (.A(_0263_),
    .B(_0268_),
    .S(_0269_),
    .Z(_0270_));
 BUF_X4 _1365_ (.A(_0730_),
    .Z(_0271_));
 MUX2_X1 _1366_ (.A(_0008_),
    .B(_0010_),
    .S(_0271_),
    .Z(_0272_));
 MUX2_X1 _1367_ (.A(_0009_),
    .B(_0011_),
    .S(_0271_),
    .Z(_0273_));
 BUF_X4 _1368_ (.A(_0734_),
    .Z(_0274_));
 MUX2_X1 _1369_ (.A(_0272_),
    .B(_0273_),
    .S(_0274_),
    .Z(_0275_));
 AND2_X1 _1370_ (.A1(_0749_),
    .A2(_0275_),
    .ZN(_0276_));
 BUF_X4 _1371_ (.A(_0730_),
    .Z(_0277_));
 MUX2_X1 _1372_ (.A(_0000_),
    .B(_0002_),
    .S(_0277_),
    .Z(_0278_));
 BUF_X4 _1373_ (.A(_0730_),
    .Z(_0279_));
 MUX2_X1 _1374_ (.A(_0001_),
    .B(_0003_),
    .S(_0279_),
    .Z(_0280_));
 MUX2_X1 _1375_ (.A(_0278_),
    .B(_0280_),
    .S(_0762_),
    .Z(_0281_));
 AND2_X1 _1376_ (.A1(_0749_),
    .A2(_0281_),
    .ZN(_0282_));
 MUX2_X1 _1377_ (.A(_0276_),
    .B(_0282_),
    .S(_0269_),
    .Z(_0283_));
 NOR4_X1 _1378_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0270_),
    .A4(_0283_),
    .ZN(net15));
 MUX2_X1 _1379_ (.A(_0028_),
    .B(_0030_),
    .S(_0279_),
    .Z(_0284_));
 MUX2_X1 _1380_ (.A(_0029_),
    .B(_0031_),
    .S(_0759_),
    .Z(_0285_));
 MUX2_X1 _1381_ (.A(_0284_),
    .B(_0285_),
    .S(_0762_),
    .Z(_0286_));
 AND2_X1 _1382_ (.A1(_0728_),
    .A2(_0286_),
    .ZN(_0287_));
 MUX2_X1 _1383_ (.A(_0020_),
    .B(_0022_),
    .S(_0264_),
    .Z(_0288_));
 MUX2_X1 _1384_ (.A(_0021_),
    .B(_0023_),
    .S(_0731_),
    .Z(_0289_));
 MUX2_X1 _1385_ (.A(_0288_),
    .B(_0289_),
    .S(_0735_),
    .Z(_0290_));
 AND2_X1 _1386_ (.A1(_0729_),
    .A2(_0290_),
    .ZN(_0291_));
 MUX2_X1 _1387_ (.A(_0287_),
    .B(_0291_),
    .S(_0269_),
    .Z(_0292_));
 MUX2_X1 _1388_ (.A(_0024_),
    .B(_0026_),
    .S(_0271_),
    .Z(_0293_));
 MUX2_X1 _1389_ (.A(_0025_),
    .B(_0027_),
    .S(_0271_),
    .Z(_0294_));
 MUX2_X1 _1390_ (.A(_0293_),
    .B(_0294_),
    .S(_0274_),
    .Z(_0295_));
 AND2_X1 _1391_ (.A1(_0748_),
    .A2(_0295_),
    .ZN(_0296_));
 MUX2_X1 _1392_ (.A(_0016_),
    .B(_0018_),
    .S(_0277_),
    .Z(_0297_));
 MUX2_X1 _1393_ (.A(_0017_),
    .B(_0019_),
    .S(_0279_),
    .Z(_0298_));
 MUX2_X1 _1394_ (.A(_0297_),
    .B(_0298_),
    .S(_0762_),
    .Z(_0299_));
 AND2_X1 _1395_ (.A1(_0749_),
    .A2(_0299_),
    .ZN(_0300_));
 MUX2_X1 _1396_ (.A(_0296_),
    .B(_0300_),
    .S(_0269_),
    .Z(_0301_));
 NOR4_X1 _1397_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0292_),
    .A4(_0301_),
    .ZN(net16));
 MUX2_X1 _1398_ (.A(_0044_),
    .B(_0046_),
    .S(_0279_),
    .Z(_0302_));
 MUX2_X1 _1399_ (.A(_0045_),
    .B(_0047_),
    .S(_0759_),
    .Z(_0303_));
 MUX2_X1 _1400_ (.A(_0302_),
    .B(_0303_),
    .S(_0762_),
    .Z(_0304_));
 AND2_X1 _1401_ (.A1(_0728_),
    .A2(_0304_),
    .ZN(_0305_));
 MUX2_X1 _1402_ (.A(_0036_),
    .B(_0038_),
    .S(_0264_),
    .Z(_0306_));
 MUX2_X1 _1403_ (.A(_0037_),
    .B(_0039_),
    .S(_0264_),
    .Z(_0307_));
 MUX2_X1 _1404_ (.A(_0306_),
    .B(_0307_),
    .S(_0735_),
    .Z(_0308_));
 AND2_X1 _1405_ (.A1(_0729_),
    .A2(_0308_),
    .ZN(_0309_));
 MUX2_X1 _1406_ (.A(_0305_),
    .B(_0309_),
    .S(_0269_),
    .Z(_0310_));
 MUX2_X1 _1407_ (.A(_0040_),
    .B(_0042_),
    .S(_0271_),
    .Z(_0311_));
 MUX2_X1 _1408_ (.A(_0041_),
    .B(_0043_),
    .S(_0271_),
    .Z(_0312_));
 MUX2_X1 _1409_ (.A(_0311_),
    .B(_0312_),
    .S(_0274_),
    .Z(_0313_));
 AND2_X1 _1410_ (.A1(_0748_),
    .A2(_0313_),
    .ZN(_0314_));
 MUX2_X1 _1411_ (.A(_0032_),
    .B(_0034_),
    .S(_0277_),
    .Z(_0315_));
 MUX2_X1 _1412_ (.A(_0033_),
    .B(_0035_),
    .S(_0279_),
    .Z(_0316_));
 MUX2_X1 _1413_ (.A(_0315_),
    .B(_0316_),
    .S(_0274_),
    .Z(_0317_));
 AND2_X1 _1414_ (.A1(_0749_),
    .A2(_0317_),
    .ZN(_0318_));
 MUX2_X1 _1415_ (.A(_0314_),
    .B(_0318_),
    .S(_0269_),
    .Z(_0319_));
 NOR4_X1 _1416_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0310_),
    .A4(_0319_),
    .ZN(net17));
 MUX2_X1 _1417_ (.A(_0060_),
    .B(_0062_),
    .S(_0279_),
    .Z(_0320_));
 MUX2_X1 _1418_ (.A(_0061_),
    .B(_0063_),
    .S(_0759_),
    .Z(_0321_));
 MUX2_X1 _1419_ (.A(_0320_),
    .B(_0321_),
    .S(_0762_),
    .Z(_0322_));
 AND2_X1 _1420_ (.A1(_0728_),
    .A2(_0322_),
    .ZN(_0323_));
 MUX2_X1 _1421_ (.A(_0052_),
    .B(_0054_),
    .S(_0264_),
    .Z(_0324_));
 MUX2_X1 _1422_ (.A(_0053_),
    .B(_0055_),
    .S(_0264_),
    .Z(_0325_));
 MUX2_X1 _1423_ (.A(_0324_),
    .B(_0325_),
    .S(_0735_),
    .Z(_0326_));
 AND2_X1 _1424_ (.A1(_0729_),
    .A2(_0326_),
    .ZN(_0327_));
 MUX2_X1 _1425_ (.A(_0323_),
    .B(_0327_),
    .S(_0269_),
    .Z(_0328_));
 MUX2_X1 _1426_ (.A(_0056_),
    .B(_0058_),
    .S(_0730_),
    .Z(_0329_));
 MUX2_X1 _1427_ (.A(_0057_),
    .B(_0059_),
    .S(_0271_),
    .Z(_0330_));
 MUX2_X1 _1428_ (.A(_0329_),
    .B(_0330_),
    .S(_0274_),
    .Z(_0331_));
 AND2_X1 _1429_ (.A1(_0748_),
    .A2(_0331_),
    .ZN(_0332_));
 MUX2_X1 _1430_ (.A(_0048_),
    .B(_0050_),
    .S(_0277_),
    .Z(_0333_));
 MUX2_X1 _1431_ (.A(_0049_),
    .B(_0051_),
    .S(_0279_),
    .Z(_0334_));
 MUX2_X1 _1432_ (.A(_0333_),
    .B(_0334_),
    .S(_0274_),
    .Z(_0335_));
 AND2_X1 _1433_ (.A1(_0749_),
    .A2(_0335_),
    .ZN(_0336_));
 MUX2_X1 _1434_ (.A(_0332_),
    .B(_0336_),
    .S(_0746_),
    .Z(_0337_));
 NOR4_X2 _1435_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0328_),
    .A4(_0337_),
    .ZN(net18));
 MUX2_X1 _1436_ (.A(_0076_),
    .B(_0078_),
    .S(_0279_),
    .Z(_0338_));
 MUX2_X1 _1437_ (.A(_0077_),
    .B(_0079_),
    .S(_0759_),
    .Z(_0339_));
 MUX2_X1 _1438_ (.A(_0338_),
    .B(_0339_),
    .S(_0762_),
    .Z(_0340_));
 AND2_X1 _1439_ (.A1(_0728_),
    .A2(_0340_),
    .ZN(_0341_));
 MUX2_X1 _1440_ (.A(_0068_),
    .B(_0070_),
    .S(_0264_),
    .Z(_0342_));
 MUX2_X1 _1441_ (.A(_0069_),
    .B(_0071_),
    .S(_0264_),
    .Z(_0343_));
 MUX2_X1 _1442_ (.A(_0342_),
    .B(_0343_),
    .S(_0735_),
    .Z(_0344_));
 AND2_X1 _1443_ (.A1(_0729_),
    .A2(_0344_),
    .ZN(_0345_));
 MUX2_X1 _1444_ (.A(_0341_),
    .B(_0345_),
    .S(_0269_),
    .Z(_0346_));
 MUX2_X1 _1445_ (.A(_0072_),
    .B(_0074_),
    .S(_0730_),
    .Z(_0347_));
 MUX2_X1 _1446_ (.A(_0073_),
    .B(_0075_),
    .S(_0271_),
    .Z(_0348_));
 MUX2_X1 _1447_ (.A(_0347_),
    .B(_0348_),
    .S(_0274_),
    .Z(_0349_));
 AND2_X1 _1448_ (.A1(_0748_),
    .A2(_0349_),
    .ZN(_0350_));
 MUX2_X1 _1449_ (.A(_0064_),
    .B(_0066_),
    .S(_0277_),
    .Z(_0351_));
 MUX2_X1 _1450_ (.A(_0065_),
    .B(_0067_),
    .S(_0277_),
    .Z(_0352_));
 MUX2_X1 _1451_ (.A(_0351_),
    .B(_0352_),
    .S(_0274_),
    .Z(_0353_));
 AND2_X1 _1452_ (.A1(_0749_),
    .A2(_0353_),
    .ZN(_0354_));
 MUX2_X1 _1453_ (.A(_0350_),
    .B(_0354_),
    .S(_0746_),
    .Z(_0355_));
 NOR4_X2 _1454_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0346_),
    .A4(_0355_),
    .ZN(net19));
 MUX2_X1 _1455_ (.A(_0092_),
    .B(_0094_),
    .S(_0279_),
    .Z(_0356_));
 MUX2_X1 _1456_ (.A(_0093_),
    .B(_0095_),
    .S(_0759_),
    .Z(_0357_));
 MUX2_X1 _1457_ (.A(_0356_),
    .B(_0357_),
    .S(_0762_),
    .Z(_0358_));
 AND2_X1 _1458_ (.A1(_0728_),
    .A2(_0358_),
    .ZN(_0359_));
 MUX2_X1 _1459_ (.A(_0084_),
    .B(_0086_),
    .S(_0759_),
    .Z(_0360_));
 MUX2_X1 _1460_ (.A(_0085_),
    .B(_0087_),
    .S(_0264_),
    .Z(_0361_));
 MUX2_X1 _1461_ (.A(_0360_),
    .B(_0361_),
    .S(_0735_),
    .Z(_0362_));
 AND2_X1 _1462_ (.A1(_0729_),
    .A2(_0362_),
    .ZN(_0363_));
 MUX2_X1 _1463_ (.A(_0359_),
    .B(_0363_),
    .S(_0269_),
    .Z(_0364_));
 MUX2_X1 _1464_ (.A(_0088_),
    .B(_0090_),
    .S(_0730_),
    .Z(_0365_));
 MUX2_X1 _1465_ (.A(_0089_),
    .B(_0091_),
    .S(_0271_),
    .Z(_0366_));
 MUX2_X1 _1466_ (.A(_0365_),
    .B(_0366_),
    .S(_0734_),
    .Z(_0367_));
 AND2_X1 _1467_ (.A1(_0748_),
    .A2(_0367_),
    .ZN(_0368_));
 MUX2_X1 _1468_ (.A(_0080_),
    .B(_0082_),
    .S(_0277_),
    .Z(_0369_));
 MUX2_X1 _1469_ (.A(_0081_),
    .B(_0083_),
    .S(_0277_),
    .Z(_0370_));
 MUX2_X1 _1470_ (.A(_0369_),
    .B(_0370_),
    .S(_0274_),
    .Z(_0371_));
 AND2_X1 _1471_ (.A1(_0749_),
    .A2(_0371_),
    .ZN(_0372_));
 MUX2_X1 _1472_ (.A(_0368_),
    .B(_0372_),
    .S(_0746_),
    .Z(_0373_));
 NOR4_X2 _1473_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0364_),
    .A4(_0373_),
    .ZN(net20));
 MUX2_X1 _1474_ (.A(_0108_),
    .B(_0110_),
    .S(_0279_),
    .Z(_0374_));
 MUX2_X1 _1475_ (.A(_0109_),
    .B(_0111_),
    .S(_0759_),
    .Z(_0375_));
 MUX2_X1 _1476_ (.A(_0374_),
    .B(_0375_),
    .S(_0762_),
    .Z(_0376_));
 AND2_X1 _1477_ (.A1(_0728_),
    .A2(_0376_),
    .ZN(_0377_));
 MUX2_X1 _1478_ (.A(_0100_),
    .B(_0102_),
    .S(_0759_),
    .Z(_0378_));
 MUX2_X1 _1479_ (.A(_0101_),
    .B(_0103_),
    .S(_0264_),
    .Z(_0379_));
 MUX2_X1 _1480_ (.A(_0378_),
    .B(_0379_),
    .S(_0762_),
    .Z(_0380_));
 AND2_X1 _1481_ (.A1(_0729_),
    .A2(_0380_),
    .ZN(_0381_));
 MUX2_X1 _1482_ (.A(_0377_),
    .B(_0381_),
    .S(_0269_),
    .Z(_0382_));
 MUX2_X1 _1483_ (.A(_0104_),
    .B(_0106_),
    .S(_0730_),
    .Z(_0383_));
 MUX2_X1 _1484_ (.A(_0105_),
    .B(_0107_),
    .S(_0271_),
    .Z(_0384_));
 MUX2_X1 _1485_ (.A(_0383_),
    .B(_0384_),
    .S(_0734_),
    .Z(_0385_));
 AND2_X1 _1486_ (.A1(_0748_),
    .A2(_0385_),
    .ZN(_0386_));
 MUX2_X1 _1487_ (.A(_0096_),
    .B(_0098_),
    .S(_0277_),
    .Z(_0387_));
 MUX2_X1 _1488_ (.A(_0097_),
    .B(_0099_),
    .S(_0277_),
    .Z(_0388_));
 MUX2_X1 _1489_ (.A(_0387_),
    .B(_0388_),
    .S(_0274_),
    .Z(_0389_));
 AND2_X1 _1490_ (.A1(_0749_),
    .A2(_0389_),
    .ZN(_0390_));
 MUX2_X1 _1491_ (.A(_0386_),
    .B(_0390_),
    .S(_0746_),
    .Z(_0391_));
 NOR4_X2 _1492_ (.A1(_0712_),
    .A2(_0726_),
    .A3(_0382_),
    .A4(_0391_),
    .ZN(net21));
 FA_X1 _1493_ (.A(_0791_),
    .B(\wr_ptr[1] ),
    .CI(_0792_),
    .CO(_0793_),
    .S(net9));
 FA_X1 _1494_ (.A(_0794_),
    .B(_0791_),
    .CI(_0795_),
    .CO(_0796_),
    .S(_0797_));
 HA_X1 _1495_ (.A(_0798_),
    .B(\wr_ptr[3] ),
    .CO(_0799_),
    .S(_0800_));
 HA_X1 _1496_ (.A(_0791_),
    .B(\wr_ptr[1] ),
    .CO(_0801_),
    .S(_0802_));
 HA_X1 _1497_ (.A(_0803_),
    .B(\wr_ptr[2] ),
    .CO(_0804_),
    .S(_0805_));
 HA_X1 _1498_ (.A(net1),
    .B(\rd_ptr[0] ),
    .CO(_0806_),
    .S(_0807_));
 HA_X1 _1499_ (.A(net2),
    .B(\rd_ptr[1] ),
    .CO(_0808_),
    .S(_0809_));
 HA_X1 _1500_ (.A(net3),
    .B(\rd_ptr[2] ),
    .CO(_0810_),
    .S(_0811_));
 HA_X1 _1501_ (.A(net2),
    .B(_0812_),
    .CO(_0813_),
    .S(_0814_));
 HA_X1 _1502_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .CO(_0815_),
    .S(_0115_));
 HA_X1 _1503_ (.A(_0112_),
    .B(_0816_),
    .CO(_0817_),
    .S(_0113_));
 HA_X1 _1504_ (.A(_0112_),
    .B(\wr_ptr[1] ),
    .CO(_0818_),
    .S(_0819_));
 HA_X1 _1505_ (.A(\wr_ptr[0] ),
    .B(_0816_),
    .CO(_0820_),
    .S(_0821_));
 HA_X1 _1506_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_0822_),
    .S(_0823_));
 HA_X1 _1507_ (.A(\rd_ptr[0] ),
    .B(_0112_),
    .CO(_0824_),
    .S(_0825_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[0][0] ),
    .QN(_0790_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[0][1] ),
    .QN(_0000_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[0][2] ),
    .QN(_0016_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[0][3] ),
    .QN(_0032_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[0][4] ),
    .QN(_0048_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[0][5] ),
    .QN(_0064_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[0][6] ),
    .QN(_0080_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[0][7] ),
    .QN(_0096_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[10][0] ),
    .QN(_0789_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][1] ),
    .QN(_0010_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][2] ),
    .QN(_0026_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[10][3] ),
    .QN(_0042_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[10][4] ),
    .QN(_0058_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[10][5] ),
    .QN(_0074_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[10][6] ),
    .QN(_0090_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[10][7] ),
    .QN(_0106_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[11][0] ),
    .QN(_0788_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][1] ),
    .QN(_0011_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][2] ),
    .QN(_0027_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[11][3] ),
    .QN(_0043_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[11][4] ),
    .QN(_0059_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[11][5] ),
    .QN(_0075_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[11][6] ),
    .QN(_0091_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[11][7] ),
    .QN(_0107_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[12][0] ),
    .QN(_0787_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[12][1] ),
    .QN(_0012_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[12][2] ),
    .QN(_0028_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[12][3] ),
    .QN(_0044_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[12][4] ),
    .QN(_0060_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[12][5] ),
    .QN(_0076_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[12][6] ),
    .QN(_0092_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[12][7] ),
    .QN(_0108_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][0] ),
    .QN(_0786_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0149_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[13][1] ),
    .QN(_0013_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0150_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[13][2] ),
    .QN(_0029_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0151_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[13][3] ),
    .QN(_0045_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0152_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[13][4] ),
    .QN(_0061_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0153_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][5] ),
    .QN(_0077_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0154_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[13][6] ),
    .QN(_0093_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0155_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][7] ),
    .QN(_0109_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0156_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[14][0] ),
    .QN(_0785_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0157_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[14][1] ),
    .QN(_0014_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0158_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[14][2] ),
    .QN(_0030_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0159_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[14][3] ),
    .QN(_0046_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0160_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[14][4] ),
    .QN(_0062_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0161_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[14][5] ),
    .QN(_0078_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0162_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[14][6] ),
    .QN(_0094_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0163_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[14][7] ),
    .QN(_0110_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0164_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[15][0] ),
    .QN(_0784_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0165_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[15][1] ),
    .QN(_0015_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0166_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[15][2] ),
    .QN(_0031_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[15][3] ),
    .QN(_0047_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[15][4] ),
    .QN(_0063_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[15][5] ),
    .QN(_0079_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[15][6] ),
    .QN(_0095_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[15][7] ),
    .QN(_0111_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[1][0] ),
    .QN(_0783_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[1][1] ),
    .QN(_0001_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[1][2] ),
    .QN(_0017_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[1][3] ),
    .QN(_0033_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[1][4] ),
    .QN(_0049_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[1][5] ),
    .QN(_0065_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[1][6] ),
    .QN(_0081_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[1][7] ),
    .QN(_0097_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[2][0] ),
    .QN(_0782_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[2][1] ),
    .QN(_0002_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[2][2] ),
    .QN(_0018_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[2][3] ),
    .QN(_0034_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[2][4] ),
    .QN(_0050_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[2][5] ),
    .QN(_0066_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[2][6] ),
    .QN(_0082_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[2][7] ),
    .QN(_0098_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[3][0] ),
    .QN(_0781_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[3][1] ),
    .QN(_0003_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[3][2] ),
    .QN(_0019_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[3][3] ),
    .QN(_0035_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0192_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[3][4] ),
    .QN(_0051_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0193_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[3][5] ),
    .QN(_0067_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0194_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[3][6] ),
    .QN(_0083_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0195_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[3][7] ),
    .QN(_0099_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0196_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[4][0] ),
    .QN(_0780_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0197_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[4][1] ),
    .QN(_0004_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0198_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[4][2] ),
    .QN(_0020_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0199_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[4][3] ),
    .QN(_0036_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0200_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[4][4] ),
    .QN(_0052_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0201_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[4][5] ),
    .QN(_0068_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0202_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[4][6] ),
    .QN(_0084_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0203_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[4][7] ),
    .QN(_0100_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0204_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[5][0] ),
    .QN(_0779_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0205_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[5][1] ),
    .QN(_0005_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0206_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[5][2] ),
    .QN(_0021_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0207_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[5][3] ),
    .QN(_0037_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0208_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[5][4] ),
    .QN(_0053_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0209_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[5][5] ),
    .QN(_0069_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0210_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[5][6] ),
    .QN(_0085_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0211_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[5][7] ),
    .QN(_0101_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0212_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[6][0] ),
    .QN(_0778_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0213_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[6][1] ),
    .QN(_0006_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0214_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[6][2] ),
    .QN(_0022_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0215_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[6][3] ),
    .QN(_0038_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0216_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[6][4] ),
    .QN(_0054_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0217_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[6][5] ),
    .QN(_0070_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0218_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[6][6] ),
    .QN(_0086_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0219_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[6][7] ),
    .QN(_0102_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0220_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[7][0] ),
    .QN(_0777_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0221_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[7][1] ),
    .QN(_0007_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0222_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[7][2] ),
    .QN(_0023_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0223_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[7][3] ),
    .QN(_0039_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0224_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[7][4] ),
    .QN(_0055_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0225_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[7][5] ),
    .QN(_0071_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0226_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[7][6] ),
    .QN(_0087_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0227_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[7][7] ),
    .QN(_0103_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0228_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[8][0] ),
    .QN(_0776_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0229_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[8][1] ),
    .QN(_0008_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0230_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[8][2] ),
    .QN(_0024_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0231_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[8][3] ),
    .QN(_0040_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0232_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[8][4] ),
    .QN(_0056_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0233_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[8][5] ),
    .QN(_0072_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0234_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[8][6] ),
    .QN(_0088_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0235_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[8][7] ),
    .QN(_0104_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0236_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[9][0] ),
    .QN(_0775_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0237_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[9][1] ),
    .QN(_0009_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0238_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[9][2] ),
    .QN(_0025_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0239_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[9][3] ),
    .QN(_0041_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0240_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[9][4] ),
    .QN(_0057_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0241_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[9][5] ),
    .QN(_0073_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0242_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[9][6] ),
    .QN(_0089_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0243_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[9][7] ),
    .QN(_0105_));
 DFF_X1 \rd_data[0]$_SDFFE_PN0P_  (.D(_0244_),
    .CK(clknet_4_7_0_clk),
    .Q(net22),
    .QN(_0774_));
 DFF_X1 \rd_data[1]$_SDFFE_PN0P_  (.D(_0245_),
    .CK(clknet_4_7_0_clk),
    .Q(net23),
    .QN(_0773_));
 DFF_X1 \rd_data[2]$_SDFFE_PN0P_  (.D(_0246_),
    .CK(clknet_4_13_0_clk),
    .Q(net24),
    .QN(_0772_));
 DFF_X1 \rd_data[3]$_SDFFE_PN0P_  (.D(_0247_),
    .CK(clknet_4_13_0_clk),
    .Q(net25),
    .QN(_0771_));
 DFF_X1 \rd_data[4]$_SDFFE_PN0P_  (.D(_0248_),
    .CK(clknet_4_7_0_clk),
    .Q(net26),
    .QN(_0770_));
 DFF_X1 \rd_data[5]$_SDFFE_PN0P_  (.D(_0249_),
    .CK(clknet_4_7_0_clk),
    .Q(net27),
    .QN(_0769_));
 DFF_X1 \rd_data[6]$_SDFFE_PN0P_  (.D(_0250_),
    .CK(clknet_4_7_0_clk),
    .Q(net28),
    .QN(_0768_));
 DFF_X1 \rd_data[7]$_SDFFE_PN0P_  (.D(_0251_),
    .CK(clknet_4_7_0_clk),
    .Q(net29),
    .QN(_0767_));
 DFF_X2 \rd_ptr[0]$_SDFFE_PN0P_  (.D(_0252_),
    .CK(clknet_4_13_0_clk),
    .Q(\rd_ptr[0] ),
    .QN(_0114_));
 DFF_X2 \rd_ptr[1]$_SDFFE_PN0P_  (.D(_0253_),
    .CK(clknet_4_13_0_clk),
    .Q(\rd_ptr[1] ),
    .QN(_0791_));
 DFF_X1 \rd_ptr[2]$_SDFFE_PN0P_  (.D(_0254_),
    .CK(clknet_4_13_0_clk),
    .Q(\rd_ptr[2] ),
    .QN(_0803_));
 DFF_X1 \rd_ptr[3]$_SDFFE_PN0P_  (.D(_0255_),
    .CK(clknet_4_15_0_clk),
    .Q(\rd_ptr[3] ),
    .QN(_0798_));
 DFF_X1 \rd_ptr[4]$_SDFFE_PN0P_  (.D(_0256_),
    .CK(clknet_4_15_0_clk),
    .Q(\rd_ptr[4] ),
    .QN(_0766_));
 DFF_X2 \wr_ptr[0]$_SDFFE_PN0P_  (.D(_0257_),
    .CK(clknet_4_15_0_clk),
    .Q(\wr_ptr[0] ),
    .QN(_0112_));
 DFF_X2 \wr_ptr[1]$_SDFFE_PN0P_  (.D(_0258_),
    .CK(clknet_4_14_0_clk),
    .Q(\wr_ptr[1] ),
    .QN(_0816_));
 DFF_X2 \wr_ptr[2]$_SDFFE_PN0P_  (.D(_0259_),
    .CK(clknet_4_15_0_clk),
    .Q(\wr_ptr[2] ),
    .QN(_0765_));
 DFF_X2 \wr_ptr[3]$_SDFFE_PN0P_  (.D(_0260_),
    .CK(clknet_4_15_0_clk),
    .Q(\wr_ptr[3] ),
    .QN(_0764_));
 DFF_X1 \wr_ptr[4]$_SDFFE_PN0P_  (.D(_0261_),
    .CK(clknet_4_15_0_clk),
    .Q(\wr_ptr[4] ),
    .QN(_0763_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_77 ();
 BUF_X1 input1 (.A(peek_addr[0]),
    .Z(net1));
 BUF_X1 input2 (.A(peek_addr[1]),
    .Z(net2));
 BUF_X1 input3 (.A(peek_addr[2]),
    .Z(net3));
 BUF_X1 input4 (.A(peek_en),
    .Z(net4));
 BUF_X1 output5 (.A(net5),
    .Z(almost_empty));
 BUF_X1 output6 (.A(net6),
    .Z(almost_full));
 BUF_X1 output7 (.A(net7),
    .Z(empty));
 BUF_X1 output8 (.A(net8),
    .Z(fifo_count[0]));
 BUF_X1 output9 (.A(net9),
    .Z(fifo_count[1]));
 BUF_X1 output10 (.A(net10),
    .Z(fifo_count[2]));
 BUF_X1 output11 (.A(net11),
    .Z(fifo_count[3]));
 BUF_X1 output12 (.A(net12),
    .Z(fifo_count[4]));
 BUF_X1 output13 (.A(net13),
    .Z(full));
 BUF_X1 output14 (.A(net14),
    .Z(peek_data[0]));
 BUF_X1 output15 (.A(net15),
    .Z(peek_data[1]));
 BUF_X1 output16 (.A(net16),
    .Z(peek_data[2]));
 BUF_X1 output17 (.A(net17),
    .Z(peek_data[3]));
 BUF_X1 output18 (.A(net18),
    .Z(peek_data[4]));
 BUF_X1 output19 (.A(net19),
    .Z(peek_data[5]));
 BUF_X1 output20 (.A(net20),
    .Z(peek_data[6]));
 BUF_X1 output21 (.A(net21),
    .Z(peek_data[7]));
 BUF_X1 output22 (.A(net22),
    .Z(rd_data[0]));
 BUF_X1 output23 (.A(net23),
    .Z(rd_data[1]));
 BUF_X1 output24 (.A(net24),
    .Z(rd_data[2]));
 BUF_X1 output25 (.A(net25),
    .Z(rd_data[3]));
 BUF_X1 output26 (.A(net26),
    .Z(rd_data[4]));
 BUF_X1 output27 (.A(net27),
    .Z(rd_data[5]));
 BUF_X1 output28 (.A(net28),
    .Z(rd_data[6]));
 BUF_X1 output29 (.A(net29),
    .Z(rd_data[7]));
 BUF_X8 max_cap30 (.A(_0403_),
    .Z(net30));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X2 clkload0 (.A(clknet_4_0_0_clk));
 INV_X1 clkload1 (.A(clknet_4_1_0_clk));
 CLKBUF_X1 clkload2 (.A(clknet_4_2_0_clk));
 INV_X2 clkload3 (.A(clknet_4_3_0_clk));
 CLKBUF_X1 clkload4 (.A(clknet_4_5_0_clk));
 INV_X2 clkload5 (.A(clknet_4_6_0_clk));
 CLKBUF_X1 clkload6 (.A(clknet_4_8_0_clk));
 INV_X1 clkload7 (.A(clknet_4_9_0_clk));
 CLKBUF_X1 clkload8 (.A(clknet_4_10_0_clk));
 INV_X1 clkload9 (.A(clknet_4_12_0_clk));
 INV_X2 clkload10 (.A(clknet_4_13_0_clk));
 INV_X1 clkload11 (.A(clknet_4_14_0_clk));
 INV_X2 clkload12 (.A(clknet_4_15_0_clk));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_21 ();
 FILLCELL_X16 FILLER_0_53 ();
 FILLCELL_X4 FILLER_0_69 ();
 FILLCELL_X1 FILLER_0_84 ();
 FILLCELL_X8 FILLER_0_89 ();
 FILLCELL_X4 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_103 ();
 FILLCELL_X8 FILLER_0_128 ();
 FILLCELL_X4 FILLER_0_136 ();
 FILLCELL_X2 FILLER_0_140 ();
 FILLCELL_X1 FILLER_0_142 ();
 FILLCELL_X1 FILLER_0_147 ();
 FILLCELL_X8 FILLER_0_154 ();
 FILLCELL_X2 FILLER_0_162 ();
 FILLCELL_X1 FILLER_0_164 ();
 FILLCELL_X16 FILLER_0_185 ();
 FILLCELL_X16 FILLER_0_225 ();
 FILLCELL_X8 FILLER_0_241 ();
 FILLCELL_X4 FILLER_0_249 ();
 FILLCELL_X16 FILLER_0_260 ();
 FILLCELL_X8 FILLER_0_276 ();
 FILLCELL_X4 FILLER_0_284 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X8 FILLER_1_23 ();
 FILLCELL_X2 FILLER_1_31 ();
 FILLCELL_X2 FILLER_1_50 ();
 FILLCELL_X1 FILLER_1_52 ();
 FILLCELL_X2 FILLER_1_60 ();
 FILLCELL_X1 FILLER_1_62 ();
 FILLCELL_X16 FILLER_1_80 ();
 FILLCELL_X8 FILLER_1_96 ();
 FILLCELL_X4 FILLER_1_104 ();
 FILLCELL_X8 FILLER_1_125 ();
 FILLCELL_X4 FILLER_1_133 ();
 FILLCELL_X8 FILLER_1_157 ();
 FILLCELL_X4 FILLER_1_189 ();
 FILLCELL_X2 FILLER_1_193 ();
 FILLCELL_X1 FILLER_1_195 ();
 FILLCELL_X16 FILLER_1_220 ();
 FILLCELL_X4 FILLER_1_236 ();
 FILLCELL_X4 FILLER_1_264 ();
 FILLCELL_X2 FILLER_1_285 ();
 FILLCELL_X1 FILLER_1_287 ();
 FILLCELL_X8 FILLER_2_1 ();
 FILLCELL_X2 FILLER_2_9 ();
 FILLCELL_X1 FILLER_2_11 ();
 FILLCELL_X1 FILLER_2_29 ();
 FILLCELL_X2 FILLER_2_37 ();
 FILLCELL_X2 FILLER_2_56 ();
 FILLCELL_X2 FILLER_2_75 ();
 FILLCELL_X16 FILLER_2_91 ();
 FILLCELL_X2 FILLER_2_107 ();
 FILLCELL_X1 FILLER_2_109 ();
 FILLCELL_X8 FILLER_2_131 ();
 FILLCELL_X4 FILLER_2_139 ();
 FILLCELL_X2 FILLER_2_143 ();
 FILLCELL_X1 FILLER_2_145 ();
 FILLCELL_X8 FILLER_2_153 ();
 FILLCELL_X4 FILLER_2_161 ();
 FILLCELL_X2 FILLER_2_165 ();
 FILLCELL_X1 FILLER_2_167 ();
 FILLCELL_X8 FILLER_2_189 ();
 FILLCELL_X2 FILLER_2_197 ();
 FILLCELL_X8 FILLER_2_211 ();
 FILLCELL_X1 FILLER_2_219 ();
 FILLCELL_X8 FILLER_2_227 ();
 FILLCELL_X2 FILLER_2_235 ();
 FILLCELL_X4 FILLER_2_268 ();
 FILLCELL_X2 FILLER_2_272 ();
 FILLCELL_X1 FILLER_2_274 ();
 FILLCELL_X4 FILLER_2_282 ();
 FILLCELL_X2 FILLER_2_286 ();
 FILLCELL_X1 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_19 ();
 FILLCELL_X1 FILLER_3_27 ();
 FILLCELL_X8 FILLER_3_35 ();
 FILLCELL_X1 FILLER_3_43 ();
 FILLCELL_X2 FILLER_3_51 ();
 FILLCELL_X1 FILLER_3_60 ();
 FILLCELL_X1 FILLER_3_68 ();
 FILLCELL_X8 FILLER_3_102 ();
 FILLCELL_X1 FILLER_3_110 ();
 FILLCELL_X1 FILLER_3_118 ();
 FILLCELL_X8 FILLER_3_133 ();
 FILLCELL_X4 FILLER_3_141 ();
 FILLCELL_X2 FILLER_3_145 ();
 FILLCELL_X1 FILLER_3_164 ();
 FILLCELL_X8 FILLER_3_172 ();
 FILLCELL_X2 FILLER_3_180 ();
 FILLCELL_X4 FILLER_3_199 ();
 FILLCELL_X4 FILLER_3_232 ();
 FILLCELL_X2 FILLER_3_236 ();
 FILLCELL_X16 FILLER_3_269 ();
 FILLCELL_X2 FILLER_3_285 ();
 FILLCELL_X1 FILLER_3_287 ();
 FILLCELL_X8 FILLER_4_1 ();
 FILLCELL_X4 FILLER_4_9 ();
 FILLCELL_X2 FILLER_4_13 ();
 FILLCELL_X1 FILLER_4_15 ();
 FILLCELL_X2 FILLER_4_23 ();
 FILLCELL_X16 FILLER_4_32 ();
 FILLCELL_X2 FILLER_4_48 ();
 FILLCELL_X8 FILLER_4_57 ();
 FILLCELL_X4 FILLER_4_65 ();
 FILLCELL_X4 FILLER_4_103 ();
 FILLCELL_X2 FILLER_4_107 ();
 FILLCELL_X8 FILLER_4_133 ();
 FILLCELL_X4 FILLER_4_141 ();
 FILLCELL_X1 FILLER_4_145 ();
 FILLCELL_X1 FILLER_4_167 ();
 FILLCELL_X4 FILLER_4_175 ();
 FILLCELL_X2 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_195 ();
 FILLCELL_X2 FILLER_4_234 ();
 FILLCELL_X32 FILLER_4_253 ();
 FILLCELL_X2 FILLER_4_285 ();
 FILLCELL_X1 FILLER_4_287 ();
 FILLCELL_X8 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_9 ();
 FILLCELL_X1 FILLER_5_13 ();
 FILLCELL_X16 FILLER_5_21 ();
 FILLCELL_X8 FILLER_5_37 ();
 FILLCELL_X2 FILLER_5_45 ();
 FILLCELL_X16 FILLER_5_54 ();
 FILLCELL_X8 FILLER_5_70 ();
 FILLCELL_X2 FILLER_5_78 ();
 FILLCELL_X1 FILLER_5_80 ();
 FILLCELL_X2 FILLER_5_88 ();
 FILLCELL_X8 FILLER_5_97 ();
 FILLCELL_X4 FILLER_5_105 ();
 FILLCELL_X1 FILLER_5_109 ();
 FILLCELL_X4 FILLER_5_141 ();
 FILLCELL_X2 FILLER_5_145 ();
 FILLCELL_X1 FILLER_5_147 ();
 FILLCELL_X8 FILLER_5_172 ();
 FILLCELL_X2 FILLER_5_180 ();
 FILLCELL_X8 FILLER_5_206 ();
 FILLCELL_X2 FILLER_5_214 ();
 FILLCELL_X4 FILLER_5_221 ();
 FILLCELL_X8 FILLER_5_232 ();
 FILLCELL_X2 FILLER_5_245 ();
 FILLCELL_X8 FILLER_5_275 ();
 FILLCELL_X4 FILLER_5_283 ();
 FILLCELL_X1 FILLER_5_287 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_30 ();
 FILLCELL_X2 FILLER_6_38 ();
 FILLCELL_X2 FILLER_6_44 ();
 FILLCELL_X8 FILLER_6_63 ();
 FILLCELL_X1 FILLER_6_71 ();
 FILLCELL_X16 FILLER_6_89 ();
 FILLCELL_X8 FILLER_6_105 ();
 FILLCELL_X1 FILLER_6_113 ();
 FILLCELL_X2 FILLER_6_121 ();
 FILLCELL_X1 FILLER_6_123 ();
 FILLCELL_X16 FILLER_6_128 ();
 FILLCELL_X4 FILLER_6_144 ();
 FILLCELL_X8 FILLER_6_179 ();
 FILLCELL_X4 FILLER_6_187 ();
 FILLCELL_X2 FILLER_6_191 ();
 FILLCELL_X16 FILLER_6_207 ();
 FILLCELL_X8 FILLER_6_223 ();
 FILLCELL_X2 FILLER_6_231 ();
 FILLCELL_X4 FILLER_6_257 ();
 FILLCELL_X1 FILLER_6_261 ();
 FILLCELL_X8 FILLER_6_279 ();
 FILLCELL_X1 FILLER_6_287 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_5 ();
 FILLCELL_X2 FILLER_7_34 ();
 FILLCELL_X1 FILLER_7_36 ();
 FILLCELL_X2 FILLER_7_68 ();
 FILLCELL_X32 FILLER_7_101 ();
 FILLCELL_X8 FILLER_7_133 ();
 FILLCELL_X1 FILLER_7_141 ();
 FILLCELL_X16 FILLER_7_166 ();
 FILLCELL_X16 FILLER_7_206 ();
 FILLCELL_X2 FILLER_7_222 ();
 FILLCELL_X16 FILLER_7_231 ();
 FILLCELL_X4 FILLER_7_247 ();
 FILLCELL_X1 FILLER_7_251 ();
 FILLCELL_X8 FILLER_7_259 ();
 FILLCELL_X1 FILLER_7_267 ();
 FILLCELL_X2 FILLER_7_285 ();
 FILLCELL_X1 FILLER_7_287 ();
 FILLCELL_X8 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_9 ();
 FILLCELL_X1 FILLER_8_13 ();
 FILLCELL_X1 FILLER_8_21 ();
 FILLCELL_X16 FILLER_8_29 ();
 FILLCELL_X16 FILLER_8_59 ();
 FILLCELL_X1 FILLER_8_75 ();
 FILLCELL_X16 FILLER_8_94 ();
 FILLCELL_X1 FILLER_8_110 ();
 FILLCELL_X2 FILLER_8_135 ();
 FILLCELL_X8 FILLER_8_168 ();
 FILLCELL_X8 FILLER_8_200 ();
 FILLCELL_X2 FILLER_8_208 ();
 FILLCELL_X1 FILLER_8_210 ();
 FILLCELL_X16 FILLER_8_228 ();
 FILLCELL_X4 FILLER_8_244 ();
 FILLCELL_X1 FILLER_8_248 ();
 FILLCELL_X4 FILLER_8_280 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_9 ();
 FILLCELL_X1 FILLER_9_11 ();
 FILLCELL_X2 FILLER_9_19 ();
 FILLCELL_X1 FILLER_9_21 ();
 FILLCELL_X8 FILLER_9_26 ();
 FILLCELL_X2 FILLER_9_34 ();
 FILLCELL_X1 FILLER_9_36 ();
 FILLCELL_X4 FILLER_9_44 ();
 FILLCELL_X16 FILLER_9_55 ();
 FILLCELL_X8 FILLER_9_71 ();
 FILLCELL_X1 FILLER_9_79 ();
 FILLCELL_X2 FILLER_9_97 ();
 FILLCELL_X4 FILLER_9_106 ();
 FILLCELL_X2 FILLER_9_110 ();
 FILLCELL_X1 FILLER_9_112 ();
 FILLCELL_X16 FILLER_9_130 ();
 FILLCELL_X4 FILLER_9_146 ();
 FILLCELL_X2 FILLER_9_150 ();
 FILLCELL_X2 FILLER_9_155 ();
 FILLCELL_X1 FILLER_9_157 ();
 FILLCELL_X16 FILLER_9_165 ();
 FILLCELL_X4 FILLER_9_181 ();
 FILLCELL_X4 FILLER_9_199 ();
 FILLCELL_X1 FILLER_9_203 ();
 FILLCELL_X1 FILLER_9_211 ();
 FILLCELL_X16 FILLER_9_233 ();
 FILLCELL_X2 FILLER_9_249 ();
 FILLCELL_X1 FILLER_9_251 ();
 FILLCELL_X8 FILLER_9_259 ();
 FILLCELL_X4 FILLER_9_274 ();
 FILLCELL_X2 FILLER_9_285 ();
 FILLCELL_X1 FILLER_9_287 ();
 FILLCELL_X4 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_22 ();
 FILLCELL_X1 FILLER_10_54 ();
 FILLCELL_X8 FILLER_10_67 ();
 FILLCELL_X2 FILLER_10_75 ();
 FILLCELL_X1 FILLER_10_77 ();
 FILLCELL_X2 FILLER_10_110 ();
 FILLCELL_X1 FILLER_10_112 ();
 FILLCELL_X4 FILLER_10_127 ();
 FILLCELL_X8 FILLER_10_138 ();
 FILLCELL_X2 FILLER_10_146 ();
 FILLCELL_X2 FILLER_10_152 ();
 FILLCELL_X8 FILLER_10_178 ();
 FILLCELL_X4 FILLER_10_186 ();
 FILLCELL_X32 FILLER_10_248 ();
 FILLCELL_X8 FILLER_10_280 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_5 ();
 FILLCELL_X8 FILLER_11_24 ();
 FILLCELL_X8 FILLER_11_60 ();
 FILLCELL_X4 FILLER_11_68 ();
 FILLCELL_X1 FILLER_11_72 ();
 FILLCELL_X2 FILLER_11_77 ();
 FILLCELL_X2 FILLER_11_83 ();
 FILLCELL_X2 FILLER_11_92 ();
 FILLCELL_X16 FILLER_11_108 ();
 FILLCELL_X1 FILLER_11_124 ();
 FILLCELL_X8 FILLER_11_136 ();
 FILLCELL_X4 FILLER_11_144 ();
 FILLCELL_X2 FILLER_11_148 ();
 FILLCELL_X1 FILLER_11_150 ();
 FILLCELL_X16 FILLER_11_186 ();
 FILLCELL_X2 FILLER_11_202 ();
 FILLCELL_X4 FILLER_11_218 ();
 FILLCELL_X1 FILLER_11_222 ();
 FILLCELL_X8 FILLER_11_230 ();
 FILLCELL_X2 FILLER_11_238 ();
 FILLCELL_X4 FILLER_11_257 ();
 FILLCELL_X2 FILLER_11_261 ();
 FILLCELL_X1 FILLER_11_263 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_9 ();
 FILLCELL_X1 FILLER_12_11 ();
 FILLCELL_X1 FILLER_12_19 ();
 FILLCELL_X8 FILLER_12_27 ();
 FILLCELL_X4 FILLER_12_35 ();
 FILLCELL_X1 FILLER_12_39 ();
 FILLCELL_X2 FILLER_12_47 ();
 FILLCELL_X1 FILLER_12_49 ();
 FILLCELL_X4 FILLER_12_68 ();
 FILLCELL_X2 FILLER_12_72 ();
 FILLCELL_X1 FILLER_12_74 ();
 FILLCELL_X2 FILLER_12_82 ();
 FILLCELL_X1 FILLER_12_84 ();
 FILLCELL_X8 FILLER_12_93 ();
 FILLCELL_X2 FILLER_12_101 ();
 FILLCELL_X1 FILLER_12_103 ();
 FILLCELL_X4 FILLER_12_108 ();
 FILLCELL_X2 FILLER_12_112 ();
 FILLCELL_X1 FILLER_12_114 ();
 FILLCELL_X2 FILLER_12_119 ();
 FILLCELL_X4 FILLER_12_125 ();
 FILLCELL_X1 FILLER_12_129 ();
 FILLCELL_X1 FILLER_12_134 ();
 FILLCELL_X2 FILLER_12_142 ();
 FILLCELL_X1 FILLER_12_144 ();
 FILLCELL_X2 FILLER_12_165 ();
 FILLCELL_X1 FILLER_12_167 ();
 FILLCELL_X8 FILLER_12_182 ();
 FILLCELL_X8 FILLER_12_193 ();
 FILLCELL_X4 FILLER_12_201 ();
 FILLCELL_X2 FILLER_12_205 ();
 FILLCELL_X4 FILLER_12_247 ();
 FILLCELL_X8 FILLER_12_278 ();
 FILLCELL_X2 FILLER_12_286 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X16 FILLER_13_6 ();
 FILLCELL_X8 FILLER_13_22 ();
 FILLCELL_X2 FILLER_13_30 ();
 FILLCELL_X1 FILLER_13_32 ();
 FILLCELL_X8 FILLER_13_36 ();
 FILLCELL_X4 FILLER_13_44 ();
 FILLCELL_X1 FILLER_13_48 ();
 FILLCELL_X1 FILLER_13_53 ();
 FILLCELL_X2 FILLER_13_71 ();
 FILLCELL_X8 FILLER_13_77 ();
 FILLCELL_X2 FILLER_13_85 ();
 FILLCELL_X2 FILLER_13_94 ();
 FILLCELL_X1 FILLER_13_96 ();
 FILLCELL_X2 FILLER_13_111 ();
 FILLCELL_X1 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_137 ();
 FILLCELL_X1 FILLER_13_145 ();
 FILLCELL_X2 FILLER_13_155 ();
 FILLCELL_X1 FILLER_13_157 ();
 FILLCELL_X2 FILLER_13_165 ();
 FILLCELL_X1 FILLER_13_176 ();
 FILLCELL_X1 FILLER_13_184 ();
 FILLCELL_X1 FILLER_13_188 ();
 FILLCELL_X2 FILLER_13_196 ();
 FILLCELL_X2 FILLER_13_215 ();
 FILLCELL_X2 FILLER_13_224 ();
 FILLCELL_X1 FILLER_13_226 ();
 FILLCELL_X1 FILLER_13_234 ();
 FILLCELL_X16 FILLER_13_257 ();
 FILLCELL_X8 FILLER_13_273 ();
 FILLCELL_X4 FILLER_13_281 ();
 FILLCELL_X2 FILLER_13_285 ();
 FILLCELL_X1 FILLER_13_287 ();
 FILLCELL_X2 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_3 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X16 FILLER_14_11 ();
 FILLCELL_X4 FILLER_14_27 ();
 FILLCELL_X1 FILLER_14_31 ();
 FILLCELL_X2 FILLER_14_49 ();
 FILLCELL_X1 FILLER_14_51 ();
 FILLCELL_X1 FILLER_14_75 ();
 FILLCELL_X4 FILLER_14_80 ();
 FILLCELL_X2 FILLER_14_104 ();
 FILLCELL_X4 FILLER_14_115 ();
 FILLCELL_X2 FILLER_14_119 ();
 FILLCELL_X2 FILLER_14_128 ();
 FILLCELL_X1 FILLER_14_130 ();
 FILLCELL_X2 FILLER_14_138 ();
 FILLCELL_X1 FILLER_14_140 ();
 FILLCELL_X16 FILLER_14_162 ();
 FILLCELL_X8 FILLER_14_178 ();
 FILLCELL_X4 FILLER_14_186 ();
 FILLCELL_X2 FILLER_14_190 ();
 FILLCELL_X8 FILLER_14_216 ();
 FILLCELL_X4 FILLER_14_224 ();
 FILLCELL_X4 FILLER_14_235 ();
 FILLCELL_X2 FILLER_14_239 ();
 FILLCELL_X16 FILLER_14_248 ();
 FILLCELL_X1 FILLER_14_264 ();
 FILLCELL_X4 FILLER_14_282 ();
 FILLCELL_X2 FILLER_14_286 ();
 FILLCELL_X2 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_3 ();
 FILLCELL_X1 FILLER_15_31 ();
 FILLCELL_X8 FILLER_15_57 ();
 FILLCELL_X2 FILLER_15_65 ();
 FILLCELL_X1 FILLER_15_67 ();
 FILLCELL_X8 FILLER_15_92 ();
 FILLCELL_X2 FILLER_15_100 ();
 FILLCELL_X2 FILLER_15_106 ();
 FILLCELL_X1 FILLER_15_108 ();
 FILLCELL_X4 FILLER_15_168 ();
 FILLCELL_X2 FILLER_15_172 ();
 FILLCELL_X1 FILLER_15_174 ();
 FILLCELL_X8 FILLER_15_178 ();
 FILLCELL_X4 FILLER_15_186 ();
 FILLCELL_X16 FILLER_15_221 ();
 FILLCELL_X2 FILLER_15_237 ();
 FILLCELL_X2 FILLER_15_264 ();
 FILLCELL_X1 FILLER_15_266 ();
 FILLCELL_X4 FILLER_15_275 ();
 FILLCELL_X2 FILLER_15_279 ();
 FILLCELL_X4 FILLER_15_284 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_9 ();
 FILLCELL_X1 FILLER_16_11 ();
 FILLCELL_X2 FILLER_16_19 ();
 FILLCELL_X4 FILLER_16_28 ();
 FILLCELL_X1 FILLER_16_32 ();
 FILLCELL_X16 FILLER_16_47 ();
 FILLCELL_X2 FILLER_16_63 ();
 FILLCELL_X1 FILLER_16_65 ();
 FILLCELL_X8 FILLER_16_90 ();
 FILLCELL_X4 FILLER_16_105 ();
 FILLCELL_X2 FILLER_16_109 ();
 FILLCELL_X1 FILLER_16_111 ();
 FILLCELL_X8 FILLER_16_139 ();
 FILLCELL_X2 FILLER_16_177 ();
 FILLCELL_X2 FILLER_16_182 ();
 FILLCELL_X1 FILLER_16_184 ();
 FILLCELL_X4 FILLER_16_188 ();
 FILLCELL_X1 FILLER_16_192 ();
 FILLCELL_X2 FILLER_16_198 ();
 FILLCELL_X4 FILLER_16_203 ();
 FILLCELL_X1 FILLER_16_213 ();
 FILLCELL_X2 FILLER_16_217 ();
 FILLCELL_X1 FILLER_16_219 ();
 FILLCELL_X4 FILLER_16_223 ();
 FILLCELL_X1 FILLER_16_233 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_43 ();
 FILLCELL_X1 FILLER_17_47 ();
 FILLCELL_X2 FILLER_17_51 ();
 FILLCELL_X16 FILLER_17_62 ();
 FILLCELL_X1 FILLER_17_92 ();
 FILLCELL_X8 FILLER_17_99 ();
 FILLCELL_X2 FILLER_17_107 ();
 FILLCELL_X4 FILLER_17_112 ();
 FILLCELL_X1 FILLER_17_116 ();
 FILLCELL_X8 FILLER_17_124 ();
 FILLCELL_X2 FILLER_17_132 ();
 FILLCELL_X2 FILLER_17_137 ();
 FILLCELL_X1 FILLER_17_139 ();
 FILLCELL_X16 FILLER_17_143 ();
 FILLCELL_X2 FILLER_17_159 ();
 FILLCELL_X1 FILLER_17_161 ();
 FILLCELL_X2 FILLER_17_178 ();
 FILLCELL_X2 FILLER_17_191 ();
 FILLCELL_X2 FILLER_17_199 ();
 FILLCELL_X1 FILLER_17_201 ();
 FILLCELL_X4 FILLER_17_205 ();
 FILLCELL_X1 FILLER_17_209 ();
 FILLCELL_X2 FILLER_17_213 ();
 FILLCELL_X4 FILLER_17_232 ();
 FILLCELL_X1 FILLER_17_236 ();
 FILLCELL_X8 FILLER_17_255 ();
 FILLCELL_X2 FILLER_17_263 ();
 FILLCELL_X4 FILLER_17_278 ();
 FILLCELL_X16 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_17 ();
 FILLCELL_X4 FILLER_18_25 ();
 FILLCELL_X1 FILLER_18_29 ();
 FILLCELL_X4 FILLER_18_44 ();
 FILLCELL_X2 FILLER_18_48 ();
 FILLCELL_X1 FILLER_18_53 ();
 FILLCELL_X1 FILLER_18_67 ();
 FILLCELL_X8 FILLER_18_71 ();
 FILLCELL_X4 FILLER_18_79 ();
 FILLCELL_X2 FILLER_18_89 ();
 FILLCELL_X1 FILLER_18_91 ();
 FILLCELL_X2 FILLER_18_99 ();
 FILLCELL_X1 FILLER_18_101 ();
 FILLCELL_X4 FILLER_18_109 ();
 FILLCELL_X2 FILLER_18_113 ();
 FILLCELL_X1 FILLER_18_115 ();
 FILLCELL_X4 FILLER_18_126 ();
 FILLCELL_X1 FILLER_18_130 ();
 FILLCELL_X1 FILLER_18_141 ();
 FILLCELL_X2 FILLER_18_147 ();
 FILLCELL_X8 FILLER_18_152 ();
 FILLCELL_X4 FILLER_18_160 ();
 FILLCELL_X2 FILLER_18_164 ();
 FILLCELL_X4 FILLER_18_202 ();
 FILLCELL_X2 FILLER_18_213 ();
 FILLCELL_X1 FILLER_18_215 ();
 FILLCELL_X2 FILLER_18_222 ();
 FILLCELL_X2 FILLER_18_255 ();
 FILLCELL_X1 FILLER_18_257 ();
 FILLCELL_X1 FILLER_18_287 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_17 ();
 FILLCELL_X1 FILLER_19_21 ();
 FILLCELL_X2 FILLER_19_29 ();
 FILLCELL_X1 FILLER_19_31 ();
 FILLCELL_X8 FILLER_19_39 ();
 FILLCELL_X8 FILLER_19_67 ();
 FILLCELL_X2 FILLER_19_75 ();
 FILLCELL_X4 FILLER_19_80 ();
 FILLCELL_X8 FILLER_19_87 ();
 FILLCELL_X8 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_106 ();
 FILLCELL_X16 FILLER_19_110 ();
 FILLCELL_X2 FILLER_19_126 ();
 FILLCELL_X1 FILLER_19_128 ();
 FILLCELL_X1 FILLER_19_144 ();
 FILLCELL_X2 FILLER_19_156 ();
 FILLCELL_X1 FILLER_19_158 ();
 FILLCELL_X8 FILLER_19_162 ();
 FILLCELL_X4 FILLER_19_170 ();
 FILLCELL_X2 FILLER_19_174 ();
 FILLCELL_X4 FILLER_19_196 ();
 FILLCELL_X2 FILLER_19_200 ();
 FILLCELL_X1 FILLER_19_202 ();
 FILLCELL_X8 FILLER_19_216 ();
 FILLCELL_X1 FILLER_19_224 ();
 FILLCELL_X16 FILLER_19_230 ();
 FILLCELL_X8 FILLER_19_246 ();
 FILLCELL_X4 FILLER_19_254 ();
 FILLCELL_X2 FILLER_19_262 ();
 FILLCELL_X1 FILLER_19_264 ();
 FILLCELL_X2 FILLER_19_274 ();
 FILLCELL_X2 FILLER_19_280 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_5 ();
 FILLCELL_X1 FILLER_20_7 ();
 FILLCELL_X4 FILLER_20_32 ();
 FILLCELL_X4 FILLER_20_43 ();
 FILLCELL_X1 FILLER_20_50 ();
 FILLCELL_X2 FILLER_20_60 ();
 FILLCELL_X2 FILLER_20_65 ();
 FILLCELL_X4 FILLER_20_70 ();
 FILLCELL_X2 FILLER_20_74 ();
 FILLCELL_X4 FILLER_20_93 ();
 FILLCELL_X2 FILLER_20_100 ();
 FILLCELL_X1 FILLER_20_105 ();
 FILLCELL_X4 FILLER_20_109 ();
 FILLCELL_X2 FILLER_20_113 ();
 FILLCELL_X1 FILLER_20_115 ();
 FILLCELL_X2 FILLER_20_136 ();
 FILLCELL_X16 FILLER_20_144 ();
 FILLCELL_X4 FILLER_20_160 ();
 FILLCELL_X1 FILLER_20_164 ();
 FILLCELL_X8 FILLER_20_168 ();
 FILLCELL_X4 FILLER_20_176 ();
 FILLCELL_X2 FILLER_20_183 ();
 FILLCELL_X1 FILLER_20_185 ();
 FILLCELL_X8 FILLER_20_197 ();
 FILLCELL_X4 FILLER_20_205 ();
 FILLCELL_X2 FILLER_20_212 ();
 FILLCELL_X1 FILLER_20_214 ();
 FILLCELL_X16 FILLER_20_235 ();
 FILLCELL_X1 FILLER_20_251 ();
 FILLCELL_X8 FILLER_20_269 ();
 FILLCELL_X2 FILLER_20_277 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_9 ();
 FILLCELL_X1 FILLER_21_11 ();
 FILLCELL_X32 FILLER_21_36 ();
 FILLCELL_X8 FILLER_21_68 ();
 FILLCELL_X16 FILLER_21_145 ();
 FILLCELL_X2 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_177 ();
 FILLCELL_X1 FILLER_21_181 ();
 FILLCELL_X8 FILLER_21_185 ();
 FILLCELL_X1 FILLER_21_193 ();
 FILLCELL_X4 FILLER_21_208 ();
 FILLCELL_X1 FILLER_21_212 ();
 FILLCELL_X2 FILLER_21_222 ();
 FILLCELL_X1 FILLER_21_224 ();
 FILLCELL_X2 FILLER_21_227 ();
 FILLCELL_X2 FILLER_21_242 ();
 FILLCELL_X4 FILLER_21_248 ();
 FILLCELL_X1 FILLER_21_252 ();
 FILLCELL_X8 FILLER_21_274 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_26 ();
 FILLCELL_X16 FILLER_22_34 ();
 FILLCELL_X1 FILLER_22_50 ();
 FILLCELL_X2 FILLER_22_77 ();
 FILLCELL_X1 FILLER_22_79 ();
 FILLCELL_X2 FILLER_22_94 ();
 FILLCELL_X4 FILLER_22_103 ();
 FILLCELL_X1 FILLER_22_107 ();
 FILLCELL_X8 FILLER_22_115 ();
 FILLCELL_X2 FILLER_22_123 ();
 FILLCELL_X16 FILLER_22_139 ();
 FILLCELL_X4 FILLER_22_155 ();
 FILLCELL_X4 FILLER_22_180 ();
 FILLCELL_X2 FILLER_22_184 ();
 FILLCELL_X1 FILLER_22_217 ();
 FILLCELL_X8 FILLER_22_241 ();
 FILLCELL_X4 FILLER_22_249 ();
 FILLCELL_X2 FILLER_22_253 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_5 ();
 FILLCELL_X1 FILLER_23_37 ();
 FILLCELL_X2 FILLER_23_46 ();
 FILLCELL_X1 FILLER_23_48 ();
 FILLCELL_X32 FILLER_23_88 ();
 FILLCELL_X8 FILLER_23_120 ();
 FILLCELL_X1 FILLER_23_135 ();
 FILLCELL_X2 FILLER_23_143 ();
 FILLCELL_X2 FILLER_23_162 ();
 FILLCELL_X1 FILLER_23_164 ();
 FILLCELL_X1 FILLER_23_174 ();
 FILLCELL_X1 FILLER_23_182 ();
 FILLCELL_X2 FILLER_23_190 ();
 FILLCELL_X1 FILLER_23_226 ();
 FILLCELL_X2 FILLER_23_240 ();
 FILLCELL_X1 FILLER_23_242 ();
 FILLCELL_X1 FILLER_23_261 ();
 FILLCELL_X16 FILLER_23_264 ();
 FILLCELL_X8 FILLER_23_280 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X8 FILLER_24_38 ();
 FILLCELL_X1 FILLER_24_46 ();
 FILLCELL_X2 FILLER_24_54 ();
 FILLCELL_X4 FILLER_24_70 ();
 FILLCELL_X2 FILLER_24_74 ();
 FILLCELL_X1 FILLER_24_76 ();
 FILLCELL_X4 FILLER_24_101 ();
 FILLCELL_X2 FILLER_24_105 ();
 FILLCELL_X2 FILLER_24_138 ();
 FILLCELL_X1 FILLER_24_140 ();
 FILLCELL_X2 FILLER_24_148 ();
 FILLCELL_X1 FILLER_24_150 ();
 FILLCELL_X8 FILLER_24_158 ();
 FILLCELL_X8 FILLER_24_176 ();
 FILLCELL_X2 FILLER_24_184 ();
 FILLCELL_X1 FILLER_24_186 ();
 FILLCELL_X4 FILLER_24_206 ();
 FILLCELL_X4 FILLER_24_213 ();
 FILLCELL_X4 FILLER_24_221 ();
 FILLCELL_X2 FILLER_24_225 ();
 FILLCELL_X4 FILLER_24_234 ();
 FILLCELL_X4 FILLER_24_271 ();
 FILLCELL_X1 FILLER_24_275 ();
 FILLCELL_X2 FILLER_24_283 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_5 ();
 FILLCELL_X2 FILLER_25_23 ();
 FILLCELL_X1 FILLER_25_25 ();
 FILLCELL_X2 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_59 ();
 FILLCELL_X4 FILLER_25_67 ();
 FILLCELL_X2 FILLER_25_71 ();
 FILLCELL_X4 FILLER_25_80 ();
 FILLCELL_X1 FILLER_25_84 ();
 FILLCELL_X2 FILLER_25_92 ();
 FILLCELL_X2 FILLER_25_101 ();
 FILLCELL_X1 FILLER_25_103 ();
 FILLCELL_X2 FILLER_25_111 ();
 FILLCELL_X1 FILLER_25_113 ();
 FILLCELL_X2 FILLER_25_131 ();
 FILLCELL_X1 FILLER_25_133 ();
 FILLCELL_X16 FILLER_25_172 ();
 FILLCELL_X2 FILLER_25_188 ();
 FILLCELL_X4 FILLER_25_216 ();
 FILLCELL_X2 FILLER_25_220 ();
 FILLCELL_X8 FILLER_25_238 ();
 FILLCELL_X8 FILLER_25_277 ();
 FILLCELL_X2 FILLER_25_285 ();
 FILLCELL_X1 FILLER_25_287 ();
 FILLCELL_X4 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_5 ();
 FILLCELL_X1 FILLER_26_7 ();
 FILLCELL_X4 FILLER_26_32 ();
 FILLCELL_X16 FILLER_26_64 ();
 FILLCELL_X4 FILLER_26_80 ();
 FILLCELL_X8 FILLER_26_101 ();
 FILLCELL_X2 FILLER_26_109 ();
 FILLCELL_X1 FILLER_26_111 ();
 FILLCELL_X4 FILLER_26_153 ();
 FILLCELL_X2 FILLER_26_157 ();
 FILLCELL_X1 FILLER_26_159 ();
 FILLCELL_X8 FILLER_26_177 ();
 FILLCELL_X4 FILLER_26_185 ();
 FILLCELL_X1 FILLER_26_189 ();
 FILLCELL_X8 FILLER_26_206 ();
 FILLCELL_X4 FILLER_26_214 ();
 FILLCELL_X2 FILLER_26_218 ();
 FILLCELL_X1 FILLER_26_220 ();
 FILLCELL_X4 FILLER_26_244 ();
 FILLCELL_X8 FILLER_26_257 ();
 FILLCELL_X1 FILLER_26_265 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X8 FILLER_27_33 ();
 FILLCELL_X4 FILLER_27_41 ();
 FILLCELL_X2 FILLER_27_45 ();
 FILLCELL_X8 FILLER_27_54 ();
 FILLCELL_X2 FILLER_27_62 ();
 FILLCELL_X1 FILLER_27_64 ();
 FILLCELL_X16 FILLER_27_69 ();
 FILLCELL_X8 FILLER_27_85 ();
 FILLCELL_X2 FILLER_27_93 ();
 FILLCELL_X8 FILLER_27_99 ();
 FILLCELL_X4 FILLER_27_107 ();
 FILLCELL_X4 FILLER_27_115 ();
 FILLCELL_X4 FILLER_27_126 ();
 FILLCELL_X1 FILLER_27_130 ();
 FILLCELL_X1 FILLER_27_142 ();
 FILLCELL_X4 FILLER_27_154 ();
 FILLCELL_X1 FILLER_27_158 ();
 FILLCELL_X2 FILLER_27_183 ();
 FILLCELL_X2 FILLER_27_211 ();
 FILLCELL_X4 FILLER_27_226 ();
 FILLCELL_X16 FILLER_27_250 ();
 FILLCELL_X4 FILLER_27_266 ();
 FILLCELL_X1 FILLER_27_270 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_29 ();
 FILLCELL_X8 FILLER_28_57 ();
 FILLCELL_X4 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_100 ();
 FILLCELL_X4 FILLER_28_132 ();
 FILLCELL_X16 FILLER_28_143 ();
 FILLCELL_X4 FILLER_28_159 ();
 FILLCELL_X8 FILLER_28_170 ();
 FILLCELL_X4 FILLER_28_178 ();
 FILLCELL_X2 FILLER_28_182 ();
 FILLCELL_X2 FILLER_28_226 ();
 FILLCELL_X2 FILLER_28_235 ();
 FILLCELL_X1 FILLER_28_237 ();
 FILLCELL_X2 FILLER_28_242 ();
 FILLCELL_X1 FILLER_28_244 ();
 FILLCELL_X16 FILLER_28_248 ();
 FILLCELL_X8 FILLER_28_264 ();
 FILLCELL_X2 FILLER_28_272 ();
 FILLCELL_X2 FILLER_28_278 ();
 FILLCELL_X4 FILLER_28_284 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_5 ();
 FILLCELL_X1 FILLER_29_30 ();
 FILLCELL_X8 FILLER_29_62 ();
 FILLCELL_X2 FILLER_29_70 ();
 FILLCELL_X1 FILLER_29_72 ();
 FILLCELL_X32 FILLER_29_104 ();
 FILLCELL_X16 FILLER_29_136 ();
 FILLCELL_X8 FILLER_29_152 ();
 FILLCELL_X4 FILLER_29_160 ();
 FILLCELL_X2 FILLER_29_164 ();
 FILLCELL_X1 FILLER_29_166 ();
 FILLCELL_X8 FILLER_29_174 ();
 FILLCELL_X1 FILLER_29_182 ();
 FILLCELL_X2 FILLER_29_275 ();
 FILLCELL_X8 FILLER_29_280 ();
 FILLCELL_X8 FILLER_30_1 ();
 FILLCELL_X2 FILLER_30_9 ();
 FILLCELL_X1 FILLER_30_11 ();
 FILLCELL_X8 FILLER_30_26 ();
 FILLCELL_X4 FILLER_30_34 ();
 FILLCELL_X8 FILLER_30_45 ();
 FILLCELL_X4 FILLER_30_60 ();
 FILLCELL_X2 FILLER_30_64 ();
 FILLCELL_X1 FILLER_30_90 ();
 FILLCELL_X8 FILLER_30_98 ();
 FILLCELL_X8 FILLER_30_130 ();
 FILLCELL_X8 FILLER_30_155 ();
 FILLCELL_X4 FILLER_30_187 ();
 FILLCELL_X2 FILLER_30_191 ();
 FILLCELL_X2 FILLER_30_251 ();
 FILLCELL_X4 FILLER_30_283 ();
 FILLCELL_X1 FILLER_30_287 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_33 ();
 FILLCELL_X4 FILLER_31_46 ();
 FILLCELL_X1 FILLER_31_50 ();
 FILLCELL_X4 FILLER_31_58 ();
 FILLCELL_X1 FILLER_31_62 ();
 FILLCELL_X4 FILLER_31_70 ();
 FILLCELL_X1 FILLER_31_74 ();
 FILLCELL_X4 FILLER_31_82 ();
 FILLCELL_X16 FILLER_31_93 ();
 FILLCELL_X2 FILLER_31_109 ();
 FILLCELL_X1 FILLER_31_118 ();
 FILLCELL_X1 FILLER_31_126 ();
 FILLCELL_X1 FILLER_31_134 ();
 FILLCELL_X1 FILLER_31_159 ();
 FILLCELL_X8 FILLER_31_177 ();
 FILLCELL_X4 FILLER_31_188 ();
 FILLCELL_X2 FILLER_31_192 ();
 FILLCELL_X1 FILLER_31_194 ();
 FILLCELL_X2 FILLER_31_202 ();
 FILLCELL_X1 FILLER_31_210 ();
 FILLCELL_X2 FILLER_31_216 ();
 FILLCELL_X1 FILLER_31_218 ();
 FILLCELL_X8 FILLER_31_226 ();
 FILLCELL_X2 FILLER_31_234 ();
 FILLCELL_X1 FILLER_31_236 ();
 FILLCELL_X8 FILLER_31_249 ();
 FILLCELL_X2 FILLER_31_264 ();
 FILLCELL_X1 FILLER_31_278 ();
 FILLCELL_X1 FILLER_31_281 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_3 ();
 FILLCELL_X1 FILLER_32_28 ();
 FILLCELL_X4 FILLER_32_56 ();
 FILLCELL_X2 FILLER_32_67 ();
 FILLCELL_X8 FILLER_32_91 ();
 FILLCELL_X4 FILLER_32_99 ();
 FILLCELL_X1 FILLER_32_103 ();
 FILLCELL_X4 FILLER_32_128 ();
 FILLCELL_X2 FILLER_32_132 ();
 FILLCELL_X32 FILLER_32_148 ();
 FILLCELL_X2 FILLER_32_180 ();
 FILLCELL_X4 FILLER_32_185 ();
 FILLCELL_X2 FILLER_32_189 ();
 FILLCELL_X4 FILLER_32_198 ();
 FILLCELL_X2 FILLER_32_202 ();
 FILLCELL_X1 FILLER_32_209 ();
 FILLCELL_X2 FILLER_32_215 ();
 FILLCELL_X8 FILLER_32_227 ();
 FILLCELL_X4 FILLER_32_235 ();
 FILLCELL_X8 FILLER_32_256 ();
 FILLCELL_X2 FILLER_32_264 ();
 FILLCELL_X1 FILLER_32_266 ();
 FILLCELL_X1 FILLER_32_284 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X1 FILLER_33_5 ();
 FILLCELL_X2 FILLER_33_30 ();
 FILLCELL_X1 FILLER_33_32 ();
 FILLCELL_X16 FILLER_33_64 ();
 FILLCELL_X4 FILLER_33_87 ();
 FILLCELL_X2 FILLER_33_91 ();
 FILLCELL_X1 FILLER_33_93 ();
 FILLCELL_X16 FILLER_33_101 ();
 FILLCELL_X4 FILLER_33_117 ();
 FILLCELL_X2 FILLER_33_121 ();
 FILLCELL_X16 FILLER_33_130 ();
 FILLCELL_X8 FILLER_33_146 ();
 FILLCELL_X4 FILLER_33_174 ();
 FILLCELL_X2 FILLER_33_178 ();
 FILLCELL_X4 FILLER_33_208 ();
 FILLCELL_X4 FILLER_33_215 ();
 FILLCELL_X2 FILLER_33_219 ();
 FILLCELL_X1 FILLER_33_240 ();
 FILLCELL_X2 FILLER_33_262 ();
 FILLCELL_X2 FILLER_33_286 ();
 FILLCELL_X8 FILLER_34_1 ();
 FILLCELL_X2 FILLER_34_9 ();
 FILLCELL_X1 FILLER_34_11 ();
 FILLCELL_X32 FILLER_34_19 ();
 FILLCELL_X16 FILLER_34_51 ();
 FILLCELL_X8 FILLER_34_67 ();
 FILLCELL_X2 FILLER_34_75 ();
 FILLCELL_X1 FILLER_34_108 ();
 FILLCELL_X4 FILLER_34_140 ();
 FILLCELL_X1 FILLER_34_144 ();
 FILLCELL_X8 FILLER_34_152 ();
 FILLCELL_X2 FILLER_34_160 ();
 FILLCELL_X1 FILLER_34_162 ();
 FILLCELL_X4 FILLER_34_176 ();
 FILLCELL_X8 FILLER_34_235 ();
 FILLCELL_X2 FILLER_34_243 ();
 FILLCELL_X2 FILLER_34_269 ();
 FILLCELL_X1 FILLER_34_271 ();
 FILLCELL_X2 FILLER_34_286 ();
 FILLCELL_X8 FILLER_35_1 ();
 FILLCELL_X1 FILLER_35_9 ();
 FILLCELL_X4 FILLER_35_41 ();
 FILLCELL_X2 FILLER_35_59 ();
 FILLCELL_X8 FILLER_35_68 ();
 FILLCELL_X2 FILLER_35_76 ();
 FILLCELL_X4 FILLER_35_95 ();
 FILLCELL_X2 FILLER_35_99 ();
 FILLCELL_X4 FILLER_35_108 ();
 FILLCELL_X4 FILLER_35_136 ();
 FILLCELL_X8 FILLER_35_147 ();
 FILLCELL_X4 FILLER_35_155 ();
 FILLCELL_X2 FILLER_35_159 ();
 FILLCELL_X1 FILLER_35_174 ();
 FILLCELL_X2 FILLER_35_185 ();
 FILLCELL_X1 FILLER_35_194 ();
 FILLCELL_X8 FILLER_35_203 ();
 FILLCELL_X4 FILLER_35_211 ();
 FILLCELL_X2 FILLER_35_215 ();
 FILLCELL_X4 FILLER_35_220 ();
 FILLCELL_X1 FILLER_35_224 ();
 FILLCELL_X2 FILLER_35_238 ();
 FILLCELL_X4 FILLER_35_271 ();
 FILLCELL_X16 FILLER_36_1 ();
 FILLCELL_X8 FILLER_36_17 ();
 FILLCELL_X4 FILLER_36_25 ();
 FILLCELL_X2 FILLER_36_29 ();
 FILLCELL_X1 FILLER_36_31 ();
 FILLCELL_X4 FILLER_36_115 ();
 FILLCELL_X1 FILLER_36_119 ();
 FILLCELL_X16 FILLER_36_151 ();
 FILLCELL_X1 FILLER_36_177 ();
 FILLCELL_X8 FILLER_36_203 ();
 FILLCELL_X2 FILLER_36_211 ();
 FILLCELL_X1 FILLER_36_224 ();
 FILLCELL_X16 FILLER_36_236 ();
 FILLCELL_X1 FILLER_36_252 ();
 FILLCELL_X8 FILLER_36_275 ();
 FILLCELL_X4 FILLER_36_283 ();
 FILLCELL_X1 FILLER_36_287 ();
 FILLCELL_X16 FILLER_37_1 ();
 FILLCELL_X4 FILLER_37_17 ();
 FILLCELL_X2 FILLER_37_21 ();
 FILLCELL_X8 FILLER_37_40 ();
 FILLCELL_X2 FILLER_37_48 ();
 FILLCELL_X1 FILLER_37_50 ();
 FILLCELL_X8 FILLER_37_68 ();
 FILLCELL_X4 FILLER_37_76 ();
 FILLCELL_X16 FILLER_37_104 ();
 FILLCELL_X4 FILLER_37_120 ();
 FILLCELL_X2 FILLER_37_124 ();
 FILLCELL_X8 FILLER_37_150 ();
 FILLCELL_X2 FILLER_37_158 ();
 FILLCELL_X1 FILLER_37_160 ();
 FILLCELL_X4 FILLER_37_180 ();
 FILLCELL_X2 FILLER_37_184 ();
 FILLCELL_X1 FILLER_37_186 ();
 FILLCELL_X1 FILLER_37_213 ();
 FILLCELL_X8 FILLER_37_248 ();
 FILLCELL_X4 FILLER_37_256 ();
 FILLCELL_X1 FILLER_37_260 ();
 FILLCELL_X16 FILLER_37_271 ();
 FILLCELL_X1 FILLER_37_287 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X16 FILLER_38_198 ();
 FILLCELL_X4 FILLER_38_214 ();
 FILLCELL_X2 FILLER_38_218 ();
 FILLCELL_X1 FILLER_38_220 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X16 FILLER_38_257 ();
 FILLCELL_X8 FILLER_38_273 ();
 FILLCELL_X4 FILLER_38_281 ();
 FILLCELL_X2 FILLER_38_285 ();
 FILLCELL_X1 FILLER_38_287 ();
endmodule
