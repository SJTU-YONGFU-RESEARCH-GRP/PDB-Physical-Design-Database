module parameterized_pwm (clk,
    enable,
    pwm_out,
    rst_n,
    div,
    duty);
 input clk;
 input enable;
 output pwm_out;
 input rst_n;
 input [15:0] div;
 input [7:0] duty;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \div_counter[0] ;
 wire \div_counter[10] ;
 wire \div_counter[11] ;
 wire \div_counter[12] ;
 wire \div_counter[13] ;
 wire \div_counter[14] ;
 wire \div_counter[15] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_counter[5] ;
 wire \div_counter[6] ;
 wire \div_counter[7] ;
 wire \div_counter[8] ;
 wire \div_counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _280_ (.A(net8),
    .ZN(_207_));
 INV_X1 _281_ (.A(net10),
    .ZN(_210_));
 INV_X1 _282_ (.A(net9),
    .ZN(_213_));
 INV_X1 _283_ (.A(net14),
    .ZN(_216_));
 INV_X1 _284_ (.A(net13),
    .ZN(_219_));
 INV_X1 _285_ (.A(net11),
    .ZN(_222_));
 INV_X1 _286_ (.A(net12),
    .ZN(_225_));
 INV_X1 _287_ (.A(net7),
    .ZN(_228_));
 INV_X1 _288_ (.A(net6),
    .ZN(_231_));
 INV_X1 _289_ (.A(net5),
    .ZN(_234_));
 INV_X1 _290_ (.A(net4),
    .ZN(_237_));
 INV_X1 _291_ (.A(net3),
    .ZN(_240_));
 INV_X1 _292_ (.A(net2),
    .ZN(_243_));
 INV_X1 _293_ (.A(net16),
    .ZN(_246_));
 INV_X1 _294_ (.A(net15),
    .ZN(_249_));
 INV_X1 _295_ (.A(net17),
    .ZN(_277_));
 BUF_X2 _296_ (.A(rst_n),
    .Z(_025_));
 INV_X1 _297_ (.A(_025_),
    .ZN(_026_));
 CLKBUF_X3 _298_ (.A(_026_),
    .Z(_027_));
 CLKBUF_X2 _299_ (.A(\counter[5] ),
    .Z(_028_));
 AND3_X1 _300_ (.A1(\counter[2] ),
    .A2(\counter[3] ),
    .A3(_252_),
    .ZN(_029_));
 AND3_X1 _301_ (.A1(_028_),
    .A2(\counter[4] ),
    .A3(_029_),
    .ZN(_030_));
 AND3_X1 _302_ (.A1(\counter[7] ),
    .A2(\counter[6] ),
    .A3(_030_),
    .ZN(_031_));
 NOR3_X1 _303_ (.A1(_027_),
    .A2(\counter[0] ),
    .A3(_031_),
    .ZN(_032_));
 AND2_X1 _304_ (.A1(_025_),
    .A2(\counter[0] ),
    .ZN(_033_));
 BUF_X2 _305_ (.A(enable),
    .Z(_034_));
 CLKBUF_X3 _306_ (.A(_034_),
    .Z(_035_));
 NOR4_X1 _307_ (.A1(net16),
    .A2(net15),
    .A3(net3),
    .A4(net6),
    .ZN(_036_));
 NOR4_X1 _308_ (.A1(net2),
    .A2(net5),
    .A3(net4),
    .A4(net7),
    .ZN(_037_));
 NOR4_X2 _309_ (.A1(net8),
    .A2(net1),
    .A3(net10),
    .A4(net13),
    .ZN(_038_));
 NOR4_X1 _310_ (.A1(net9),
    .A2(net12),
    .A3(net11),
    .A4(net14),
    .ZN(_039_));
 AND4_X2 _311_ (.A1(_036_),
    .A2(_037_),
    .A3(_038_),
    .A4(_039_),
    .ZN(_040_));
 AND4_X1 _312_ (.A1(_230_),
    .A2(_239_),
    .A3(_236_),
    .A4(_233_),
    .ZN(_041_));
 AND4_X1 _313_ (.A1(_242_),
    .A2(_251_),
    .A3(_248_),
    .A4(_245_),
    .ZN(_042_));
 AND2_X2 _314_ (.A1(_041_),
    .A2(_042_),
    .ZN(_043_));
 AOI21_X1 _315_ (.A(_217_),
    .B1(_220_),
    .B2(_218_),
    .ZN(_044_));
 AOI21_X1 _316_ (.A(_226_),
    .B1(_223_),
    .B2(_227_),
    .ZN(_045_));
 NAND2_X1 _317_ (.A1(_218_),
    .A2(_221_),
    .ZN(_046_));
 OAI21_X2 _318_ (.A(_044_),
    .B1(_045_),
    .B2(_046_),
    .ZN(_047_));
 NAND2_X1 _319_ (.A1(_043_),
    .A2(_047_),
    .ZN(_048_));
 OAI21_X2 _320_ (.A(_230_),
    .B1(_233_),
    .B2(_232_),
    .ZN(_049_));
 NOR2_X1 _321_ (.A1(_232_),
    .A2(_235_),
    .ZN(_050_));
 NAND2_X1 _322_ (.A1(_236_),
    .A2(_238_),
    .ZN(_051_));
 AOI21_X4 _323_ (.A(_049_),
    .B1(_050_),
    .B2(_051_),
    .ZN(_052_));
 AOI21_X1 _324_ (.A(_241_),
    .B1(_244_),
    .B2(_242_),
    .ZN(_053_));
 AOI21_X1 _325_ (.A(_247_),
    .B1(_250_),
    .B2(_248_),
    .ZN(_054_));
 NAND2_X1 _326_ (.A1(_242_),
    .A2(_245_),
    .ZN(_055_));
 OAI21_X1 _327_ (.A(_053_),
    .B1(_054_),
    .B2(_055_),
    .ZN(_056_));
 AOI211_X2 _328_ (.A(_229_),
    .B(_052_),
    .C1(_056_),
    .C2(_041_),
    .ZN(_057_));
 INV_X1 _329_ (.A(_212_),
    .ZN(_058_));
 INV_X1 _330_ (.A(_214_),
    .ZN(_059_));
 NAND3_X1 _331_ (.A1(_209_),
    .A2(_206_),
    .A3(_215_),
    .ZN(_060_));
 AOI21_X1 _332_ (.A(_058_),
    .B1(_059_),
    .B2(_060_),
    .ZN(_061_));
 NOR2_X1 _333_ (.A1(_208_),
    .A2(_211_),
    .ZN(_062_));
 INV_X1 _334_ (.A(_209_),
    .ZN(_063_));
 OAI21_X1 _335_ (.A(_062_),
    .B1(_205_),
    .B2(_063_),
    .ZN(_064_));
 INV_X1 _336_ (.A(_211_),
    .ZN(_065_));
 NAND2_X1 _337_ (.A1(_212_),
    .A2(_215_),
    .ZN(_066_));
 NAND2_X1 _338_ (.A1(_065_),
    .A2(_066_),
    .ZN(_067_));
 AOI21_X2 _339_ (.A(_061_),
    .B1(_064_),
    .B2(_067_),
    .ZN(_068_));
 AND2_X1 _340_ (.A1(_218_),
    .A2(_221_),
    .ZN(_069_));
 NAND4_X2 _341_ (.A1(_227_),
    .A2(_224_),
    .A3(_043_),
    .A4(_069_),
    .ZN(_070_));
 OAI211_X4 _342_ (.A(_048_),
    .B(_057_),
    .C1(_068_),
    .C2(_070_),
    .ZN(_071_));
 OAI21_X2 _343_ (.A(_035_),
    .B1(_040_),
    .B2(_071_),
    .ZN(_072_));
 MUX2_X1 _344_ (.A(_032_),
    .B(_033_),
    .S(_072_),
    .Z(_000_));
 AND2_X1 _345_ (.A1(_025_),
    .A2(_253_),
    .ZN(_073_));
 AND2_X1 _346_ (.A1(_025_),
    .A2(\counter[1] ),
    .ZN(_074_));
 MUX2_X1 _347_ (.A(_073_),
    .B(_074_),
    .S(_072_),
    .Z(_001_));
 AND2_X1 _348_ (.A1(_025_),
    .A2(\counter[2] ),
    .ZN(_075_));
 NOR2_X1 _349_ (.A1(_027_),
    .A2(\counter[2] ),
    .ZN(_076_));
 NAND2_X1 _350_ (.A1(_035_),
    .A2(_252_),
    .ZN(_077_));
 AND2_X1 _351_ (.A1(_041_),
    .A2(_056_),
    .ZN(_078_));
 NOR4_X4 _352_ (.A1(_229_),
    .A2(_078_),
    .A3(_040_),
    .A4(_052_),
    .ZN(_079_));
 INV_X1 _353_ (.A(_205_),
    .ZN(_080_));
 AOI21_X1 _354_ (.A(_208_),
    .B1(_080_),
    .B2(_209_),
    .ZN(_081_));
 AND2_X1 _355_ (.A1(_059_),
    .A2(_060_),
    .ZN(_082_));
 OAI221_X2 _356_ (.A(_065_),
    .B1(_066_),
    .B2(_081_),
    .C1(_082_),
    .C2(_058_),
    .ZN(_083_));
 AND4_X1 _357_ (.A1(_227_),
    .A2(_224_),
    .A3(_043_),
    .A4(_069_),
    .ZN(_084_));
 AOI22_X4 _358_ (.A1(_083_),
    .A2(_084_),
    .B1(_047_),
    .B2(_043_),
    .ZN(_085_));
 AOI21_X1 _359_ (.A(_077_),
    .B1(_079_),
    .B2(_085_),
    .ZN(_086_));
 MUX2_X1 _360_ (.A(_075_),
    .B(_076_),
    .S(_086_),
    .Z(_002_));
 INV_X1 _361_ (.A(\counter[3] ),
    .ZN(_087_));
 AND3_X1 _362_ (.A1(\counter[2] ),
    .A2(\counter[0] ),
    .A3(\counter[1] ),
    .ZN(_088_));
 INV_X1 _363_ (.A(_034_),
    .ZN(_089_));
 NOR2_X1 _364_ (.A1(_026_),
    .A2(_089_),
    .ZN(_090_));
 NAND3_X1 _365_ (.A1(_087_),
    .A2(_088_),
    .A3(_090_),
    .ZN(_091_));
 AOI21_X1 _366_ (.A(_091_),
    .B1(_079_),
    .B2(_085_),
    .ZN(_092_));
 NAND2_X1 _367_ (.A1(_025_),
    .A2(\counter[3] ),
    .ZN(_093_));
 NOR3_X1 _368_ (.A1(_040_),
    .A2(_071_),
    .A3(_093_),
    .ZN(_094_));
 NOR3_X1 _369_ (.A1(_031_),
    .A2(_088_),
    .A3(_093_),
    .ZN(_095_));
 NOR3_X1 _370_ (.A1(_027_),
    .A2(_035_),
    .A3(_087_),
    .ZN(_096_));
 OR4_X1 _371_ (.A1(_092_),
    .A2(_094_),
    .A3(_095_),
    .A4(_096_),
    .ZN(_003_));
 AND2_X1 _372_ (.A1(_025_),
    .A2(\counter[4] ),
    .ZN(_097_));
 NOR2_X1 _373_ (.A1(_027_),
    .A2(\counter[4] ),
    .ZN(_098_));
 NAND2_X1 _374_ (.A1(_035_),
    .A2(_029_),
    .ZN(_099_));
 AOI21_X1 _375_ (.A(_099_),
    .B1(_079_),
    .B2(_085_),
    .ZN(_100_));
 MUX2_X1 _376_ (.A(_097_),
    .B(_098_),
    .S(_100_),
    .Z(_004_));
 INV_X1 _377_ (.A(_028_),
    .ZN(_101_));
 AND3_X1 _378_ (.A1(\counter[4] ),
    .A2(\counter[3] ),
    .A3(_088_),
    .ZN(_102_));
 AND3_X1 _379_ (.A1(_101_),
    .A2(_090_),
    .A3(_102_),
    .ZN(_103_));
 OAI21_X1 _380_ (.A(_103_),
    .B1(_071_),
    .B2(_040_),
    .ZN(_104_));
 NAND2_X1 _381_ (.A1(_025_),
    .A2(_028_),
    .ZN(_105_));
 OR3_X1 _382_ (.A1(_040_),
    .A2(_071_),
    .A3(_105_),
    .ZN(_106_));
 NOR3_X1 _383_ (.A1(_031_),
    .A2(_102_),
    .A3(_105_),
    .ZN(_107_));
 NOR2_X1 _384_ (.A1(_027_),
    .A2(_035_),
    .ZN(_108_));
 AOI21_X1 _385_ (.A(_107_),
    .B1(_108_),
    .B2(_028_),
    .ZN(_109_));
 NAND3_X1 _386_ (.A1(_104_),
    .A2(_106_),
    .A3(_109_),
    .ZN(_005_));
 NOR2_X1 _387_ (.A1(_027_),
    .A2(\counter[6] ),
    .ZN(_110_));
 INV_X1 _388_ (.A(\counter[6] ),
    .ZN(_111_));
 NOR2_X1 _389_ (.A1(_027_),
    .A2(_111_),
    .ZN(_112_));
 AND2_X1 _390_ (.A1(_034_),
    .A2(_030_),
    .ZN(_113_));
 OAI21_X1 _391_ (.A(_113_),
    .B1(_071_),
    .B2(_040_),
    .ZN(_114_));
 MUX2_X1 _392_ (.A(_110_),
    .B(_112_),
    .S(_114_),
    .Z(_006_));
 INV_X1 _393_ (.A(\counter[7] ),
    .ZN(_115_));
 AOI21_X1 _394_ (.A(_030_),
    .B1(_102_),
    .B2(_028_),
    .ZN(_116_));
 OR3_X1 _395_ (.A1(_089_),
    .A2(_111_),
    .A3(_116_),
    .ZN(_117_));
 AOI21_X1 _396_ (.A(_117_),
    .B1(_079_),
    .B2(_085_),
    .ZN(_118_));
 NAND4_X1 _397_ (.A1(_025_),
    .A2(_115_),
    .A3(_028_),
    .A4(_102_),
    .ZN(_119_));
 OAI33_X1 _398_ (.A1(_027_),
    .A2(_115_),
    .A3(_118_),
    .B1(_119_),
    .B2(_111_),
    .B3(_072_),
    .ZN(_007_));
 OR3_X1 _399_ (.A1(_089_),
    .A2(\div_counter[0] ),
    .A3(_071_),
    .ZN(_120_));
 NAND2_X1 _400_ (.A1(_089_),
    .A2(\div_counter[0] ),
    .ZN(_121_));
 AOI21_X1 _401_ (.A(_027_),
    .B1(_120_),
    .B2(_121_),
    .ZN(_008_));
 AOI21_X2 _402_ (.A(_027_),
    .B1(_035_),
    .B2(_071_),
    .ZN(_122_));
 BUF_X2 _403_ (.A(_122_),
    .Z(_123_));
 BUF_X1 _404_ (.A(\div_counter[10] ),
    .Z(_124_));
 AND3_X1 _405_ (.A1(\div_counter[2] ),
    .A2(\div_counter[3] ),
    .A3(\div_counter[4] ),
    .ZN(_125_));
 NAND2_X1 _406_ (.A1(_254_),
    .A2(_125_),
    .ZN(_126_));
 INV_X1 _407_ (.A(\div_counter[8] ),
    .ZN(_127_));
 INV_X1 _408_ (.A(\div_counter[9] ),
    .ZN(_128_));
 CLKBUF_X2 _409_ (.A(\div_counter[5] ),
    .Z(_129_));
 NAND4_X2 _410_ (.A1(_034_),
    .A2(_129_),
    .A3(\div_counter[6] ),
    .A4(\div_counter[7] ),
    .ZN(_130_));
 OR3_X1 _411_ (.A1(_127_),
    .A2(_128_),
    .A3(_130_),
    .ZN(_131_));
 OR2_X1 _412_ (.A1(_126_),
    .A2(_131_),
    .ZN(_132_));
 XNOR2_X1 _413_ (.A(_124_),
    .B(_132_),
    .ZN(_133_));
 AND2_X1 _414_ (.A1(_123_),
    .A2(_133_),
    .ZN(_009_));
 BUF_X1 _415_ (.A(\div_counter[11] ),
    .Z(_134_));
 NAND3_X2 _416_ (.A1(\div_counter[0] ),
    .A2(\div_counter[1] ),
    .A3(_125_),
    .ZN(_135_));
 NOR2_X1 _417_ (.A1(_131_),
    .A2(_135_),
    .ZN(_136_));
 NAND2_X1 _418_ (.A1(_124_),
    .A2(_136_),
    .ZN(_137_));
 XNOR2_X1 _419_ (.A(_134_),
    .B(_137_),
    .ZN(_138_));
 AND2_X1 _420_ (.A1(_123_),
    .A2(_138_),
    .ZN(_010_));
 NAND2_X1 _421_ (.A1(_124_),
    .A2(_134_),
    .ZN(_139_));
 NOR2_X1 _422_ (.A1(_132_),
    .A2(_139_),
    .ZN(_140_));
 XOR2_X1 _423_ (.A(\div_counter[12] ),
    .B(_140_),
    .Z(_141_));
 AND2_X1 _424_ (.A1(_123_),
    .A2(_141_),
    .ZN(_011_));
 NAND4_X1 _425_ (.A1(_124_),
    .A2(_134_),
    .A3(\div_counter[12] ),
    .A4(_136_),
    .ZN(_142_));
 XNOR2_X1 _426_ (.A(\div_counter[13] ),
    .B(_142_),
    .ZN(_143_));
 AND2_X1 _427_ (.A1(_123_),
    .A2(_143_),
    .ZN(_012_));
 INV_X1 _428_ (.A(\div_counter[14] ),
    .ZN(_144_));
 NAND4_X1 _429_ (.A1(_124_),
    .A2(_134_),
    .A3(\div_counter[12] ),
    .A4(\div_counter[13] ),
    .ZN(_145_));
 NOR2_X1 _430_ (.A1(_132_),
    .A2(_145_),
    .ZN(_146_));
 XNOR2_X1 _431_ (.A(_144_),
    .B(_146_),
    .ZN(_147_));
 AND2_X1 _432_ (.A1(_123_),
    .A2(_147_),
    .ZN(_013_));
 OR4_X1 _433_ (.A1(_144_),
    .A2(_131_),
    .A3(_135_),
    .A4(_145_),
    .ZN(_148_));
 XNOR2_X1 _434_ (.A(\div_counter[15] ),
    .B(_148_),
    .ZN(_149_));
 AND2_X1 _435_ (.A1(_123_),
    .A2(_149_),
    .ZN(_014_));
 NAND2_X1 _436_ (.A1(_089_),
    .A2(\div_counter[1] ),
    .ZN(_150_));
 NAND2_X1 _437_ (.A1(_035_),
    .A2(_255_),
    .ZN(_151_));
 OAI21_X1 _438_ (.A(_150_),
    .B1(_151_),
    .B2(_071_),
    .ZN(_152_));
 AND2_X1 _439_ (.A1(_025_),
    .A2(_152_),
    .ZN(_015_));
 NAND2_X1 _440_ (.A1(_035_),
    .A2(_254_),
    .ZN(_153_));
 XNOR2_X1 _441_ (.A(\div_counter[2] ),
    .B(_153_),
    .ZN(_154_));
 AND2_X1 _442_ (.A1(_123_),
    .A2(_154_),
    .ZN(_016_));
 NAND4_X2 _443_ (.A1(_034_),
    .A2(\div_counter[0] ),
    .A3(\div_counter[2] ),
    .A4(\div_counter[1] ),
    .ZN(_155_));
 XNOR2_X1 _444_ (.A(\div_counter[3] ),
    .B(_155_),
    .ZN(_156_));
 AND2_X1 _445_ (.A1(_123_),
    .A2(_156_),
    .ZN(_017_));
 NAND4_X1 _446_ (.A1(_035_),
    .A2(_254_),
    .A3(\div_counter[2] ),
    .A4(\div_counter[3] ),
    .ZN(_157_));
 XNOR2_X1 _447_ (.A(\div_counter[4] ),
    .B(_157_),
    .ZN(_158_));
 AND2_X1 _448_ (.A1(_123_),
    .A2(_158_),
    .ZN(_018_));
 NAND2_X1 _449_ (.A1(\div_counter[3] ),
    .A2(\div_counter[4] ),
    .ZN(_159_));
 NOR2_X1 _450_ (.A1(_155_),
    .A2(_159_),
    .ZN(_160_));
 XOR2_X1 _451_ (.A(_129_),
    .B(_160_),
    .Z(_161_));
 AND2_X1 _452_ (.A1(_123_),
    .A2(_161_),
    .ZN(_019_));
 NAND4_X1 _453_ (.A1(_035_),
    .A2(_254_),
    .A3(_129_),
    .A4(_125_),
    .ZN(_162_));
 XNOR2_X1 _454_ (.A(\div_counter[6] ),
    .B(_162_),
    .ZN(_163_));
 AND2_X1 _455_ (.A1(_122_),
    .A2(_163_),
    .ZN(_020_));
 NAND3_X1 _456_ (.A1(_034_),
    .A2(_129_),
    .A3(\div_counter[6] ),
    .ZN(_164_));
 NOR2_X1 _457_ (.A1(_164_),
    .A2(_135_),
    .ZN(_165_));
 XOR2_X1 _458_ (.A(\div_counter[7] ),
    .B(_165_),
    .Z(_166_));
 AND2_X1 _459_ (.A1(_122_),
    .A2(_166_),
    .ZN(_021_));
 NOR2_X1 _460_ (.A1(_126_),
    .A2(_130_),
    .ZN(_167_));
 XNOR2_X1 _461_ (.A(_127_),
    .B(_167_),
    .ZN(_168_));
 AND2_X1 _462_ (.A1(_122_),
    .A2(_168_),
    .ZN(_022_));
 NOR3_X1 _463_ (.A1(_127_),
    .A2(_130_),
    .A3(_135_),
    .ZN(_169_));
 XNOR2_X1 _464_ (.A(_128_),
    .B(_169_),
    .ZN(_170_));
 AND2_X1 _465_ (.A1(_122_),
    .A2(_170_),
    .ZN(_023_));
 AND3_X1 _466_ (.A1(_258_),
    .A2(_261_),
    .A3(_264_),
    .ZN(_171_));
 INV_X1 _467_ (.A(_257_),
    .ZN(_172_));
 AOI21_X1 _468_ (.A(_260_),
    .B1(_263_),
    .B2(_261_),
    .ZN(_173_));
 INV_X1 _469_ (.A(_258_),
    .ZN(_174_));
 OAI21_X1 _470_ (.A(_172_),
    .B1(_173_),
    .B2(_174_),
    .ZN(_175_));
 AND2_X1 _471_ (.A1(_276_),
    .A2(_279_),
    .ZN(_176_));
 NAND4_X1 _472_ (.A1(_267_),
    .A2(_273_),
    .A3(_171_),
    .A4(_176_),
    .ZN(_177_));
 INV_X1 _473_ (.A(_270_),
    .ZN(_178_));
 OAI221_X1 _474_ (.A(_090_),
    .B1(_171_),
    .B2(_175_),
    .C1(_177_),
    .C2(_178_),
    .ZN(_179_));
 NOR2_X1 _475_ (.A1(_266_),
    .A2(_175_),
    .ZN(_180_));
 INV_X1 _476_ (.A(_275_),
    .ZN(_181_));
 INV_X1 _477_ (.A(_276_),
    .ZN(_182_));
 OAI21_X1 _478_ (.A(_181_),
    .B1(_278_),
    .B2(_182_),
    .ZN(_183_));
 AOI21_X1 _479_ (.A(_272_),
    .B1(_183_),
    .B2(_273_),
    .ZN(_184_));
 NOR2_X1 _480_ (.A1(_178_),
    .A2(_184_),
    .ZN(_185_));
 OAI21_X1 _481_ (.A(_267_),
    .B1(_269_),
    .B2(_185_),
    .ZN(_186_));
 AOI21_X1 _482_ (.A(_179_),
    .B1(_180_),
    .B2(_186_),
    .ZN(_024_));
 HA_X1 _483_ (.A(net1),
    .B(_204_),
    .CO(_205_),
    .S(_206_));
 HA_X1 _484_ (.A(_207_),
    .B(\div_counter[1] ),
    .CO(_208_),
    .S(_209_));
 HA_X1 _485_ (.A(_210_),
    .B(\div_counter[3] ),
    .CO(_211_),
    .S(_212_));
 HA_X1 _486_ (.A(_213_),
    .B(\div_counter[2] ),
    .CO(_214_),
    .S(_215_));
 HA_X1 _487_ (.A(_216_),
    .B(\div_counter[7] ),
    .CO(_217_),
    .S(_218_));
 HA_X1 _488_ (.A(_219_),
    .B(\div_counter[6] ),
    .CO(_220_),
    .S(_221_));
 HA_X1 _489_ (.A(_222_),
    .B(\div_counter[4] ),
    .CO(_223_),
    .S(_224_));
 HA_X1 _490_ (.A(_225_),
    .B(\div_counter[5] ),
    .CO(_226_),
    .S(_227_));
 HA_X1 _491_ (.A(_228_),
    .B(\div_counter[15] ),
    .CO(_229_),
    .S(_230_));
 HA_X1 _492_ (.A(_231_),
    .B(\div_counter[14] ),
    .CO(_232_),
    .S(_233_));
 HA_X1 _493_ (.A(_234_),
    .B(\div_counter[13] ),
    .CO(_235_),
    .S(_236_));
 HA_X1 _494_ (.A(_237_),
    .B(\div_counter[12] ),
    .CO(_238_),
    .S(_239_));
 HA_X1 _495_ (.A(_240_),
    .B(\div_counter[11] ),
    .CO(_241_),
    .S(_242_));
 HA_X1 _496_ (.A(_243_),
    .B(\div_counter[10] ),
    .CO(_244_),
    .S(_245_));
 HA_X1 _497_ (.A(_246_),
    .B(\div_counter[9] ),
    .CO(_247_),
    .S(_248_));
 HA_X1 _498_ (.A(_249_),
    .B(\div_counter[8] ),
    .CO(_250_),
    .S(_251_));
 HA_X1 _499_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_252_),
    .S(_253_));
 HA_X1 _500_ (.A(\div_counter[0] ),
    .B(\div_counter[1] ),
    .CO(_254_),
    .S(_255_));
 HA_X1 _501_ (.A(_256_),
    .B(net24),
    .CO(_257_),
    .S(_258_));
 HA_X1 _502_ (.A(_259_),
    .B(net23),
    .CO(_260_),
    .S(_261_));
 HA_X1 _503_ (.A(_262_),
    .B(net22),
    .CO(_263_),
    .S(_264_));
 HA_X1 _504_ (.A(_265_),
    .B(net21),
    .CO(_266_),
    .S(_267_));
 HA_X1 _505_ (.A(_268_),
    .B(net20),
    .CO(_269_),
    .S(_270_));
 HA_X1 _506_ (.A(_271_),
    .B(net19),
    .CO(_272_),
    .S(_273_));
 HA_X1 _507_ (.A(_274_),
    .B(net18),
    .CO(_275_),
    .S(_276_));
 HA_X1 _508_ (.A(\counter[0] ),
    .B(_277_),
    .CO(_278_),
    .S(_279_));
 DFF_X2 \counter[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[0] ),
    .QN(_203_));
 DFF_X1 \counter[1]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[1] ),
    .QN(_274_));
 DFF_X1 \counter[2]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[2] ),
    .QN(_271_));
 DFF_X1 \counter[3]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[3] ),
    .QN(_268_));
 DFF_X1 \counter[4]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[4] ),
    .QN(_265_));
 DFF_X1 \counter[5]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[5] ),
    .QN(_262_));
 DFF_X1 \counter[6]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[6] ),
    .QN(_259_));
 DFF_X1 \counter[7]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[7] ),
    .QN(_256_));
 DFF_X2 \div_counter[0]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\div_counter[0] ),
    .QN(_204_));
 DFF_X1 \div_counter[10]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[10] ),
    .QN(_202_));
 DFF_X1 \div_counter[11]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[11] ),
    .QN(_201_));
 DFF_X2 \div_counter[12]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[12] ),
    .QN(_200_));
 DFF_X1 \div_counter[13]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[13] ),
    .QN(_199_));
 DFF_X1 \div_counter[14]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[14] ),
    .QN(_198_));
 DFF_X1 \div_counter[15]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[15] ),
    .QN(_197_));
 DFF_X2 \div_counter[1]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\div_counter[1] ),
    .QN(_196_));
 DFF_X2 \div_counter[2]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[2] ),
    .QN(_195_));
 DFF_X2 \div_counter[3]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[3] ),
    .QN(_194_));
 DFF_X2 \div_counter[4]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[4] ),
    .QN(_193_));
 DFF_X1 \div_counter[5]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[5] ),
    .QN(_192_));
 DFF_X2 \div_counter[6]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[6] ),
    .QN(_191_));
 DFF_X2 \div_counter[7]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[7] ),
    .QN(_190_));
 DFF_X1 \div_counter[8]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[8] ),
    .QN(_189_));
 DFF_X1 \div_counter[9]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\div_counter[9] ),
    .QN(_188_));
 DFF_X1 \pwm_reg$_SDFF_PN0_  (.D(_024_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net25),
    .QN(_187_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_89 ();
 BUF_X1 input1 (.A(div[0]),
    .Z(net1));
 BUF_X1 input2 (.A(div[10]),
    .Z(net2));
 BUF_X1 input3 (.A(div[11]),
    .Z(net3));
 BUF_X1 input4 (.A(div[12]),
    .Z(net4));
 BUF_X1 input5 (.A(div[13]),
    .Z(net5));
 BUF_X1 input6 (.A(div[14]),
    .Z(net6));
 BUF_X1 input7 (.A(div[15]),
    .Z(net7));
 BUF_X1 input8 (.A(div[1]),
    .Z(net8));
 BUF_X1 input9 (.A(div[2]),
    .Z(net9));
 BUF_X1 input10 (.A(div[3]),
    .Z(net10));
 BUF_X1 input11 (.A(div[4]),
    .Z(net11));
 BUF_X1 input12 (.A(div[5]),
    .Z(net12));
 BUF_X1 input13 (.A(div[6]),
    .Z(net13));
 BUF_X1 input14 (.A(div[7]),
    .Z(net14));
 BUF_X1 input15 (.A(div[8]),
    .Z(net15));
 BUF_X1 input16 (.A(div[9]),
    .Z(net16));
 BUF_X1 input17 (.A(duty[0]),
    .Z(net17));
 BUF_X1 input18 (.A(duty[1]),
    .Z(net18));
 BUF_X1 input19 (.A(duty[2]),
    .Z(net19));
 BUF_X1 input20 (.A(duty[3]),
    .Z(net20));
 BUF_X1 input21 (.A(duty[4]),
    .Z(net21));
 BUF_X1 input22 (.A(duty[5]),
    .Z(net22));
 BUF_X1 input23 (.A(duty[6]),
    .Z(net23));
 BUF_X1 input24 (.A(duty[7]),
    .Z(net24));
 BUF_X1 output25 (.A(net25),
    .Z(pwm_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X2 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X16 FILLER_0_129 ();
 FILLCELL_X8 FILLER_0_148 ();
 FILLCELL_X4 FILLER_0_156 ();
 FILLCELL_X2 FILLER_0_160 ();
 FILLCELL_X2 FILLER_0_165 ();
 FILLCELL_X1 FILLER_0_167 ();
 FILLCELL_X2 FILLER_0_171 ();
 FILLCELL_X32 FILLER_0_176 ();
 FILLCELL_X32 FILLER_0_208 ();
 FILLCELL_X32 FILLER_0_240 ();
 FILLCELL_X32 FILLER_0_272 ();
 FILLCELL_X32 FILLER_0_304 ();
 FILLCELL_X2 FILLER_0_336 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_161 ();
 FILLCELL_X1 FILLER_1_165 ();
 FILLCELL_X32 FILLER_1_169 ();
 FILLCELL_X32 FILLER_1_201 ();
 FILLCELL_X32 FILLER_1_233 ();
 FILLCELL_X32 FILLER_1_265 ();
 FILLCELL_X32 FILLER_1_297 ();
 FILLCELL_X8 FILLER_1_329 ();
 FILLCELL_X1 FILLER_1_337 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X16 FILLER_2_321 ();
 FILLCELL_X1 FILLER_2_337 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X16 FILLER_3_321 ();
 FILLCELL_X1 FILLER_3_337 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X16 FILLER_4_321 ();
 FILLCELL_X1 FILLER_4_337 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X16 FILLER_5_321 ();
 FILLCELL_X1 FILLER_5_337 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X16 FILLER_6_321 ();
 FILLCELL_X1 FILLER_6_337 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X16 FILLER_7_321 ();
 FILLCELL_X1 FILLER_7_337 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X2 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_172 ();
 FILLCELL_X32 FILLER_8_204 ();
 FILLCELL_X32 FILLER_8_236 ();
 FILLCELL_X32 FILLER_8_268 ();
 FILLCELL_X32 FILLER_8_300 ();
 FILLCELL_X4 FILLER_8_332 ();
 FILLCELL_X2 FILLER_8_336 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X16 FILLER_9_129 ();
 FILLCELL_X8 FILLER_9_145 ();
 FILLCELL_X4 FILLER_9_153 ();
 FILLCELL_X2 FILLER_9_163 ();
 FILLCELL_X1 FILLER_9_165 ();
 FILLCELL_X4 FILLER_9_168 ();
 FILLCELL_X32 FILLER_9_182 ();
 FILLCELL_X32 FILLER_9_214 ();
 FILLCELL_X32 FILLER_9_246 ();
 FILLCELL_X32 FILLER_9_278 ();
 FILLCELL_X16 FILLER_9_310 ();
 FILLCELL_X8 FILLER_9_326 ();
 FILLCELL_X4 FILLER_9_334 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X8 FILLER_10_129 ();
 FILLCELL_X4 FILLER_10_137 ();
 FILLCELL_X2 FILLER_10_141 ();
 FILLCELL_X1 FILLER_10_143 ();
 FILLCELL_X2 FILLER_10_146 ();
 FILLCELL_X1 FILLER_10_148 ();
 FILLCELL_X32 FILLER_10_180 ();
 FILLCELL_X32 FILLER_10_212 ();
 FILLCELL_X32 FILLER_10_244 ();
 FILLCELL_X32 FILLER_10_276 ();
 FILLCELL_X16 FILLER_10_308 ();
 FILLCELL_X8 FILLER_10_324 ();
 FILLCELL_X4 FILLER_10_332 ();
 FILLCELL_X2 FILLER_10_336 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X8 FILLER_11_129 ();
 FILLCELL_X4 FILLER_11_137 ();
 FILLCELL_X1 FILLER_11_141 ();
 FILLCELL_X4 FILLER_11_152 ();
 FILLCELL_X32 FILLER_11_181 ();
 FILLCELL_X1 FILLER_11_213 ();
 FILLCELL_X32 FILLER_11_218 ();
 FILLCELL_X32 FILLER_11_250 ();
 FILLCELL_X32 FILLER_11_282 ();
 FILLCELL_X16 FILLER_11_314 ();
 FILLCELL_X8 FILLER_11_330 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X16 FILLER_12_140 ();
 FILLCELL_X32 FILLER_12_173 ();
 FILLCELL_X32 FILLER_12_205 ();
 FILLCELL_X32 FILLER_12_237 ();
 FILLCELL_X32 FILLER_12_269 ();
 FILLCELL_X32 FILLER_12_301 ();
 FILLCELL_X4 FILLER_12_333 ();
 FILLCELL_X1 FILLER_12_337 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_9 ();
 FILLCELL_X2 FILLER_13_13 ();
 FILLCELL_X32 FILLER_13_34 ();
 FILLCELL_X32 FILLER_13_66 ();
 FILLCELL_X16 FILLER_13_98 ();
 FILLCELL_X4 FILLER_13_114 ();
 FILLCELL_X2 FILLER_13_118 ();
 FILLCELL_X32 FILLER_13_139 ();
 FILLCELL_X32 FILLER_13_171 ();
 FILLCELL_X32 FILLER_13_203 ();
 FILLCELL_X8 FILLER_13_235 ();
 FILLCELL_X1 FILLER_13_243 ();
 FILLCELL_X32 FILLER_13_261 ();
 FILLCELL_X16 FILLER_13_293 ();
 FILLCELL_X4 FILLER_13_309 ();
 FILLCELL_X2 FILLER_13_313 ();
 FILLCELL_X1 FILLER_13_315 ();
 FILLCELL_X2 FILLER_13_329 ();
 FILLCELL_X1 FILLER_13_331 ();
 FILLCELL_X2 FILLER_13_335 ();
 FILLCELL_X1 FILLER_13_337 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X32 FILLER_14_34 ();
 FILLCELL_X32 FILLER_14_66 ();
 FILLCELL_X16 FILLER_14_98 ();
 FILLCELL_X2 FILLER_14_114 ();
 FILLCELL_X1 FILLER_14_116 ();
 FILLCELL_X32 FILLER_14_137 ();
 FILLCELL_X32 FILLER_14_169 ();
 FILLCELL_X8 FILLER_14_201 ();
 FILLCELL_X4 FILLER_14_209 ();
 FILLCELL_X1 FILLER_14_213 ();
 FILLCELL_X8 FILLER_14_233 ();
 FILLCELL_X1 FILLER_14_241 ();
 FILLCELL_X32 FILLER_14_253 ();
 FILLCELL_X16 FILLER_14_285 ();
 FILLCELL_X8 FILLER_14_301 ();
 FILLCELL_X4 FILLER_14_309 ();
 FILLCELL_X2 FILLER_14_313 ();
 FILLCELL_X1 FILLER_14_327 ();
 FILLCELL_X8 FILLER_14_330 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X16 FILLER_15_27 ();
 FILLCELL_X1 FILLER_15_43 ();
 FILLCELL_X32 FILLER_15_61 ();
 FILLCELL_X32 FILLER_15_93 ();
 FILLCELL_X1 FILLER_15_125 ();
 FILLCELL_X2 FILLER_15_129 ();
 FILLCELL_X2 FILLER_15_136 ();
 FILLCELL_X1 FILLER_15_138 ();
 FILLCELL_X16 FILLER_15_148 ();
 FILLCELL_X4 FILLER_15_164 ();
 FILLCELL_X2 FILLER_15_168 ();
 FILLCELL_X1 FILLER_15_170 ();
 FILLCELL_X8 FILLER_15_209 ();
 FILLCELL_X2 FILLER_15_217 ();
 FILLCELL_X1 FILLER_15_219 ();
 FILLCELL_X8 FILLER_15_231 ();
 FILLCELL_X1 FILLER_15_239 ();
 FILLCELL_X32 FILLER_15_254 ();
 FILLCELL_X16 FILLER_15_286 ();
 FILLCELL_X8 FILLER_15_302 ();
 FILLCELL_X2 FILLER_15_310 ();
 FILLCELL_X2 FILLER_15_316 ();
 FILLCELL_X1 FILLER_15_318 ();
 FILLCELL_X1 FILLER_15_321 ();
 FILLCELL_X8 FILLER_15_326 ();
 FILLCELL_X4 FILLER_15_334 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X1 FILLER_16_21 ();
 FILLCELL_X2 FILLER_16_25 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X1 FILLER_16_49 ();
 FILLCELL_X2 FILLER_16_65 ();
 FILLCELL_X1 FILLER_16_73 ();
 FILLCELL_X4 FILLER_16_101 ();
 FILLCELL_X2 FILLER_16_105 ();
 FILLCELL_X1 FILLER_16_107 ();
 FILLCELL_X4 FILLER_16_112 ();
 FILLCELL_X2 FILLER_16_116 ();
 FILLCELL_X1 FILLER_16_118 ();
 FILLCELL_X1 FILLER_16_125 ();
 FILLCELL_X1 FILLER_16_129 ();
 FILLCELL_X1 FILLER_16_135 ();
 FILLCELL_X1 FILLER_16_139 ();
 FILLCELL_X8 FILLER_16_147 ();
 FILLCELL_X4 FILLER_16_155 ();
 FILLCELL_X1 FILLER_16_159 ();
 FILLCELL_X2 FILLER_16_170 ();
 FILLCELL_X1 FILLER_16_188 ();
 FILLCELL_X16 FILLER_16_196 ();
 FILLCELL_X8 FILLER_16_212 ();
 FILLCELL_X4 FILLER_16_220 ();
 FILLCELL_X1 FILLER_16_224 ();
 FILLCELL_X16 FILLER_16_229 ();
 FILLCELL_X8 FILLER_16_245 ();
 FILLCELL_X2 FILLER_16_253 ();
 FILLCELL_X4 FILLER_16_263 ();
 FILLCELL_X2 FILLER_16_267 ();
 FILLCELL_X2 FILLER_16_283 ();
 FILLCELL_X8 FILLER_16_302 ();
 FILLCELL_X4 FILLER_16_310 ();
 FILLCELL_X2 FILLER_16_324 ();
 FILLCELL_X1 FILLER_16_326 ();
 FILLCELL_X8 FILLER_16_330 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_17 ();
 FILLCELL_X2 FILLER_17_29 ();
 FILLCELL_X16 FILLER_17_36 ();
 FILLCELL_X8 FILLER_17_52 ();
 FILLCELL_X4 FILLER_17_60 ();
 FILLCELL_X2 FILLER_17_64 ();
 FILLCELL_X1 FILLER_17_66 ();
 FILLCELL_X32 FILLER_17_70 ();
 FILLCELL_X2 FILLER_17_102 ();
 FILLCELL_X32 FILLER_17_123 ();
 FILLCELL_X16 FILLER_17_155 ();
 FILLCELL_X4 FILLER_17_171 ();
 FILLCELL_X2 FILLER_17_175 ();
 FILLCELL_X4 FILLER_17_180 ();
 FILLCELL_X2 FILLER_17_184 ();
 FILLCELL_X32 FILLER_17_188 ();
 FILLCELL_X16 FILLER_17_220 ();
 FILLCELL_X8 FILLER_17_236 ();
 FILLCELL_X4 FILLER_17_244 ();
 FILLCELL_X2 FILLER_17_248 ();
 FILLCELL_X1 FILLER_17_250 ();
 FILLCELL_X2 FILLER_17_254 ();
 FILLCELL_X32 FILLER_17_265 ();
 FILLCELL_X16 FILLER_17_297 ();
 FILLCELL_X16 FILLER_17_322 ();
 FILLCELL_X16 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_17 ();
 FILLCELL_X1 FILLER_18_21 ();
 FILLCELL_X32 FILLER_18_25 ();
 FILLCELL_X8 FILLER_18_57 ();
 FILLCELL_X2 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_71 ();
 FILLCELL_X16 FILLER_18_103 ();
 FILLCELL_X4 FILLER_18_119 ();
 FILLCELL_X2 FILLER_18_123 ();
 FILLCELL_X1 FILLER_18_131 ();
 FILLCELL_X2 FILLER_18_135 ();
 FILLCELL_X1 FILLER_18_137 ();
 FILLCELL_X32 FILLER_18_143 ();
 FILLCELL_X16 FILLER_18_175 ();
 FILLCELL_X8 FILLER_18_191 ();
 FILLCELL_X8 FILLER_18_204 ();
 FILLCELL_X1 FILLER_18_212 ();
 FILLCELL_X32 FILLER_18_215 ();
 FILLCELL_X1 FILLER_18_251 ();
 FILLCELL_X1 FILLER_18_270 ();
 FILLCELL_X16 FILLER_18_288 ();
 FILLCELL_X4 FILLER_18_304 ();
 FILLCELL_X1 FILLER_18_308 ();
 FILLCELL_X8 FILLER_18_327 ();
 FILLCELL_X2 FILLER_18_335 ();
 FILLCELL_X1 FILLER_18_337 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X1 FILLER_19_13 ();
 FILLCELL_X1 FILLER_19_26 ();
 FILLCELL_X1 FILLER_19_37 ();
 FILLCELL_X1 FILLER_19_41 ();
 FILLCELL_X1 FILLER_19_49 ();
 FILLCELL_X1 FILLER_19_53 ();
 FILLCELL_X32 FILLER_19_64 ();
 FILLCELL_X8 FILLER_19_96 ();
 FILLCELL_X2 FILLER_19_104 ();
 FILLCELL_X1 FILLER_19_106 ();
 FILLCELL_X32 FILLER_19_111 ();
 FILLCELL_X8 FILLER_19_143 ();
 FILLCELL_X4 FILLER_19_151 ();
 FILLCELL_X2 FILLER_19_155 ();
 FILLCELL_X32 FILLER_19_174 ();
 FILLCELL_X4 FILLER_19_206 ();
 FILLCELL_X1 FILLER_19_213 ();
 FILLCELL_X2 FILLER_19_219 ();
 FILLCELL_X8 FILLER_19_228 ();
 FILLCELL_X8 FILLER_19_244 ();
 FILLCELL_X4 FILLER_19_252 ();
 FILLCELL_X32 FILLER_19_267 ();
 FILLCELL_X8 FILLER_19_299 ();
 FILLCELL_X4 FILLER_19_307 ();
 FILLCELL_X2 FILLER_19_311 ();
 FILLCELL_X8 FILLER_19_323 ();
 FILLCELL_X4 FILLER_19_331 ();
 FILLCELL_X2 FILLER_19_335 ();
 FILLCELL_X1 FILLER_19_337 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_9 ();
 FILLCELL_X2 FILLER_20_13 ();
 FILLCELL_X1 FILLER_20_15 ();
 FILLCELL_X2 FILLER_20_24 ();
 FILLCELL_X1 FILLER_20_26 ();
 FILLCELL_X1 FILLER_20_39 ();
 FILLCELL_X1 FILLER_20_46 ();
 FILLCELL_X2 FILLER_20_60 ();
 FILLCELL_X1 FILLER_20_62 ();
 FILLCELL_X2 FILLER_20_94 ();
 FILLCELL_X4 FILLER_20_122 ();
 FILLCELL_X8 FILLER_20_140 ();
 FILLCELL_X2 FILLER_20_148 ();
 FILLCELL_X1 FILLER_20_159 ();
 FILLCELL_X4 FILLER_20_163 ();
 FILLCELL_X2 FILLER_20_167 ();
 FILLCELL_X32 FILLER_20_181 ();
 FILLCELL_X4 FILLER_20_218 ();
 FILLCELL_X2 FILLER_20_222 ();
 FILLCELL_X8 FILLER_20_228 ();
 FILLCELL_X1 FILLER_20_236 ();
 FILLCELL_X1 FILLER_20_242 ();
 FILLCELL_X2 FILLER_20_248 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X2 FILLER_20_260 ();
 FILLCELL_X4 FILLER_20_265 ();
 FILLCELL_X2 FILLER_20_269 ();
 FILLCELL_X4 FILLER_20_278 ();
 FILLCELL_X1 FILLER_20_282 ();
 FILLCELL_X8 FILLER_20_300 ();
 FILLCELL_X4 FILLER_20_308 ();
 FILLCELL_X2 FILLER_20_312 ();
 FILLCELL_X2 FILLER_20_321 ();
 FILLCELL_X1 FILLER_20_323 ();
 FILLCELL_X4 FILLER_20_334 ();
 FILLCELL_X4 FILLER_21_4 ();
 FILLCELL_X4 FILLER_21_11 ();
 FILLCELL_X2 FILLER_21_18 ();
 FILLCELL_X1 FILLER_21_20 ();
 FILLCELL_X4 FILLER_21_26 ();
 FILLCELL_X8 FILLER_21_32 ();
 FILLCELL_X2 FILLER_21_40 ();
 FILLCELL_X8 FILLER_21_56 ();
 FILLCELL_X4 FILLER_21_64 ();
 FILLCELL_X1 FILLER_21_68 ();
 FILLCELL_X8 FILLER_21_74 ();
 FILLCELL_X2 FILLER_21_82 ();
 FILLCELL_X1 FILLER_21_84 ();
 FILLCELL_X1 FILLER_21_92 ();
 FILLCELL_X16 FILLER_21_100 ();
 FILLCELL_X4 FILLER_21_116 ();
 FILLCELL_X2 FILLER_21_120 ();
 FILLCELL_X4 FILLER_21_134 ();
 FILLCELL_X1 FILLER_21_138 ();
 FILLCELL_X8 FILLER_21_143 ();
 FILLCELL_X2 FILLER_21_151 ();
 FILLCELL_X16 FILLER_21_176 ();
 FILLCELL_X4 FILLER_21_192 ();
 FILLCELL_X1 FILLER_21_196 ();
 FILLCELL_X8 FILLER_21_205 ();
 FILLCELL_X1 FILLER_21_213 ();
 FILLCELL_X4 FILLER_21_230 ();
 FILLCELL_X2 FILLER_21_234 ();
 FILLCELL_X1 FILLER_21_236 ();
 FILLCELL_X8 FILLER_21_254 ();
 FILLCELL_X8 FILLER_21_266 ();
 FILLCELL_X32 FILLER_21_281 ();
 FILLCELL_X2 FILLER_21_333 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_21 ();
 FILLCELL_X8 FILLER_22_25 ();
 FILLCELL_X4 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_40 ();
 FILLCELL_X32 FILLER_22_72 ();
 FILLCELL_X32 FILLER_22_104 ();
 FILLCELL_X16 FILLER_22_136 ();
 FILLCELL_X4 FILLER_22_152 ();
 FILLCELL_X2 FILLER_22_156 ();
 FILLCELL_X1 FILLER_22_158 ();
 FILLCELL_X16 FILLER_22_168 ();
 FILLCELL_X8 FILLER_22_184 ();
 FILLCELL_X4 FILLER_22_192 ();
 FILLCELL_X2 FILLER_22_196 ();
 FILLCELL_X4 FILLER_22_211 ();
 FILLCELL_X2 FILLER_22_215 ();
 FILLCELL_X2 FILLER_22_219 ();
 FILLCELL_X1 FILLER_22_221 ();
 FILLCELL_X16 FILLER_22_229 ();
 FILLCELL_X1 FILLER_22_245 ();
 FILLCELL_X4 FILLER_22_250 ();
 FILLCELL_X2 FILLER_22_254 ();
 FILLCELL_X1 FILLER_22_256 ();
 FILLCELL_X32 FILLER_22_261 ();
 FILLCELL_X32 FILLER_22_293 ();
 FILLCELL_X8 FILLER_22_325 ();
 FILLCELL_X4 FILLER_22_333 ();
 FILLCELL_X1 FILLER_22_337 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_5 ();
 FILLCELL_X2 FILLER_23_32 ();
 FILLCELL_X32 FILLER_23_37 ();
 FILLCELL_X32 FILLER_23_69 ();
 FILLCELL_X16 FILLER_23_101 ();
 FILLCELL_X2 FILLER_23_117 ();
 FILLCELL_X16 FILLER_23_121 ();
 FILLCELL_X4 FILLER_23_137 ();
 FILLCELL_X2 FILLER_23_141 ();
 FILLCELL_X32 FILLER_23_164 ();
 FILLCELL_X4 FILLER_23_196 ();
 FILLCELL_X2 FILLER_23_200 ();
 FILLCELL_X1 FILLER_23_202 ();
 FILLCELL_X4 FILLER_23_237 ();
 FILLCELL_X2 FILLER_23_241 ();
 FILLCELL_X1 FILLER_23_243 ();
 FILLCELL_X32 FILLER_23_261 ();
 FILLCELL_X32 FILLER_23_293 ();
 FILLCELL_X8 FILLER_23_325 ();
 FILLCELL_X4 FILLER_23_333 ();
 FILLCELL_X1 FILLER_23_337 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_12 ();
 FILLCELL_X1 FILLER_24_14 ();
 FILLCELL_X4 FILLER_24_18 ();
 FILLCELL_X1 FILLER_24_25 ();
 FILLCELL_X1 FILLER_24_40 ();
 FILLCELL_X1 FILLER_24_46 ();
 FILLCELL_X2 FILLER_24_50 ();
 FILLCELL_X16 FILLER_24_62 ();
 FILLCELL_X4 FILLER_24_78 ();
 FILLCELL_X2 FILLER_24_82 ();
 FILLCELL_X1 FILLER_24_84 ();
 FILLCELL_X2 FILLER_24_94 ();
 FILLCELL_X16 FILLER_24_99 ();
 FILLCELL_X8 FILLER_24_115 ();
 FILLCELL_X4 FILLER_24_123 ();
 FILLCELL_X2 FILLER_24_127 ();
 FILLCELL_X1 FILLER_24_129 ();
 FILLCELL_X2 FILLER_24_139 ();
 FILLCELL_X1 FILLER_24_141 ();
 FILLCELL_X4 FILLER_24_152 ();
 FILLCELL_X2 FILLER_24_156 ();
 FILLCELL_X1 FILLER_24_158 ();
 FILLCELL_X32 FILLER_24_169 ();
 FILLCELL_X32 FILLER_24_201 ();
 FILLCELL_X32 FILLER_24_233 ();
 FILLCELL_X32 FILLER_24_265 ();
 FILLCELL_X8 FILLER_24_297 ();
 FILLCELL_X2 FILLER_24_305 ();
 FILLCELL_X8 FILLER_24_330 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_9 ();
 FILLCELL_X4 FILLER_25_27 ();
 FILLCELL_X2 FILLER_25_31 ();
 FILLCELL_X1 FILLER_25_33 ();
 FILLCELL_X1 FILLER_25_51 ();
 FILLCELL_X16 FILLER_25_66 ();
 FILLCELL_X2 FILLER_25_82 ();
 FILLCELL_X1 FILLER_25_84 ();
 FILLCELL_X16 FILLER_25_103 ();
 FILLCELL_X8 FILLER_25_119 ();
 FILLCELL_X4 FILLER_25_127 ();
 FILLCELL_X4 FILLER_25_138 ();
 FILLCELL_X2 FILLER_25_142 ();
 FILLCELL_X32 FILLER_25_163 ();
 FILLCELL_X32 FILLER_25_195 ();
 FILLCELL_X32 FILLER_25_227 ();
 FILLCELL_X32 FILLER_25_259 ();
 FILLCELL_X16 FILLER_25_291 ();
 FILLCELL_X4 FILLER_25_307 ();
 FILLCELL_X1 FILLER_25_311 ();
 FILLCELL_X4 FILLER_25_332 ();
 FILLCELL_X2 FILLER_25_336 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X16 FILLER_26_33 ();
 FILLCELL_X1 FILLER_26_49 ();
 FILLCELL_X2 FILLER_26_64 ();
 FILLCELL_X1 FILLER_26_83 ();
 FILLCELL_X1 FILLER_26_90 ();
 FILLCELL_X16 FILLER_26_108 ();
 FILLCELL_X2 FILLER_26_124 ();
 FILLCELL_X32 FILLER_26_136 ();
 FILLCELL_X16 FILLER_26_168 ();
 FILLCELL_X8 FILLER_26_184 ();
 FILLCELL_X4 FILLER_26_192 ();
 FILLCELL_X2 FILLER_26_196 ();
 FILLCELL_X1 FILLER_26_198 ();
 FILLCELL_X32 FILLER_26_203 ();
 FILLCELL_X32 FILLER_26_235 ();
 FILLCELL_X32 FILLER_26_267 ();
 FILLCELL_X16 FILLER_26_299 ();
 FILLCELL_X2 FILLER_26_315 ();
 FILLCELL_X1 FILLER_26_317 ();
 FILLCELL_X8 FILLER_26_328 ();
 FILLCELL_X2 FILLER_26_336 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_97 ();
 FILLCELL_X8 FILLER_27_113 ();
 FILLCELL_X2 FILLER_27_121 ();
 FILLCELL_X1 FILLER_27_123 ();
 FILLCELL_X32 FILLER_27_143 ();
 FILLCELL_X32 FILLER_27_175 ();
 FILLCELL_X32 FILLER_27_207 ();
 FILLCELL_X32 FILLER_27_239 ();
 FILLCELL_X32 FILLER_27_271 ();
 FILLCELL_X32 FILLER_27_303 ();
 FILLCELL_X2 FILLER_27_335 ();
 FILLCELL_X1 FILLER_27_337 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X2 FILLER_28_321 ();
 FILLCELL_X8 FILLER_28_326 ();
 FILLCELL_X4 FILLER_28_334 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X16 FILLER_29_321 ();
 FILLCELL_X1 FILLER_29_337 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X16 FILLER_30_321 ();
 FILLCELL_X1 FILLER_30_337 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X16 FILLER_31_321 ();
 FILLCELL_X1 FILLER_31_337 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X16 FILLER_32_321 ();
 FILLCELL_X1 FILLER_32_337 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X16 FILLER_33_321 ();
 FILLCELL_X1 FILLER_33_337 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X16 FILLER_34_321 ();
 FILLCELL_X1 FILLER_34_337 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X16 FILLER_35_321 ();
 FILLCELL_X1 FILLER_35_337 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X16 FILLER_36_321 ();
 FILLCELL_X1 FILLER_36_337 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X16 FILLER_37_321 ();
 FILLCELL_X1 FILLER_37_337 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X16 FILLER_38_321 ();
 FILLCELL_X1 FILLER_38_337 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X16 FILLER_39_321 ();
 FILLCELL_X1 FILLER_39_337 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X16 FILLER_40_321 ();
 FILLCELL_X1 FILLER_40_337 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X16 FILLER_41_321 ();
 FILLCELL_X1 FILLER_41_337 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X16 FILLER_42_321 ();
 FILLCELL_X1 FILLER_42_337 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X16 FILLER_43_321 ();
 FILLCELL_X1 FILLER_43_337 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X16 FILLER_44_321 ();
 FILLCELL_X1 FILLER_44_337 ();
endmodule
