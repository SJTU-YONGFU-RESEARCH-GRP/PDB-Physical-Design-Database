module configurable_mult (sign_mode,
    a,
    b,
    product);
 input sign_mode;
 input [7:0] a;
 input [7:0] b;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _022_;
 wire net1;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire net5;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire _494_;
 wire _495_;
 wire _496_;
 wire _497_;
 wire _498_;
 wire _499_;
 wire _500_;
 wire _501_;
 wire _502_;
 wire _503_;
 wire _504_;
 wire _505_;
 wire _506_;
 wire _507_;
 wire _508_;
 wire _509_;
 wire _510_;
 wire _511_;
 wire _512_;
 wire _513_;
 wire _514_;
 wire _515_;
 wire _516_;
 wire _517_;
 wire _518_;
 wire _519_;
 wire _520_;
 wire _521_;
 wire _522_;
 wire _523_;
 wire _524_;
 wire _525_;
 wire _526_;
 wire _527_;
 wire _528_;
 wire _529_;
 wire _530_;
 wire _531_;
 wire _532_;
 wire _533_;
 wire _534_;
 wire _535_;
 wire _536_;
 wire _537_;
 wire net2;
 wire net3;
 wire net4;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net44;
 wire net50;

 BUF_X8 _538_ (.A(b[0]),
    .Z(_000_));
 BUF_X8 _539_ (.A(a[1]),
    .Z(_001_));
 AND2_X1 _540_ (.A1(net5),
    .A2(_001_),
    .ZN(_415_));
 BUF_X16 _541_ (.A(a[0]),
    .Z(_002_));
 BUF_X16 _542_ (.A(b[1]),
    .Z(_003_));
 AND2_X1 _543_ (.A1(_002_),
    .A2(_003_),
    .ZN(_414_));
 BUF_X8 _544_ (.A(b[2]),
    .Z(_004_));
 NAND2_X1 _545_ (.A1(_002_),
    .A2(_004_),
    .ZN(_139_));
 BUF_X16 _546_ (.A(a[3]),
    .Z(_005_));
 NAND2_X1 _547_ (.A1(net5),
    .A2(_005_),
    .ZN(_144_));
 BUF_X16 _548_ (.A(a[2]),
    .Z(_006_));
 NAND2_X1 _549_ (.A1(_003_),
    .A2(_006_),
    .ZN(_145_));
 NAND2_X1 _550_ (.A1(_001_),
    .A2(_004_),
    .ZN(_146_));
 BUF_X8 _551_ (.A(b[3]),
    .Z(_007_));
 NAND2_X1 _552_ (.A1(_002_),
    .A2(_007_),
    .ZN(_149_));
 BUF_X8 _553_ (.A(a[4]),
    .Z(_008_));
 NAND2_X1 _554_ (.A1(_000_),
    .A2(_008_),
    .ZN(_153_));
 NAND2_X1 _555_ (.A1(_003_),
    .A2(_005_),
    .ZN(_152_));
 NAND2_X1 _556_ (.A1(_006_),
    .A2(_004_),
    .ZN(_154_));
 AND2_X1 _557_ (.A1(_001_),
    .A2(_007_),
    .ZN(_424_));
 BUF_X8 _558_ (.A(b[4]),
    .Z(_009_));
 AND2_X1 _559_ (.A1(_002_),
    .A2(_009_),
    .ZN(_425_));
 BUF_X8 _560_ (.A(a[5]),
    .Z(_010_));
 NAND2_X1 _561_ (.A1(_000_),
    .A2(_010_),
    .ZN(_162_));
 NAND2_X1 _562_ (.A1(_003_),
    .A2(_008_),
    .ZN(_160_));
 NAND2_X1 _563_ (.A1(_004_),
    .A2(_005_),
    .ZN(_161_));
 BUF_X16 _564_ (.A(b[5]),
    .Z(_011_));
 NAND2_X4 _565_ (.A1(_011_),
    .A2(_002_),
    .ZN(_167_));
 BUF_X4 _566_ (.A(a[6]),
    .Z(_012_));
 NAND2_X1 _567_ (.A1(_000_),
    .A2(_012_),
    .ZN(_179_));
 NAND2_X1 _568_ (.A1(_003_),
    .A2(_010_),
    .ZN(_178_));
 NAND2_X1 _569_ (.A1(_004_),
    .A2(_008_),
    .ZN(_177_));
 NAND2_X1 _570_ (.A1(_001_),
    .A2(_011_),
    .ZN(_182_));
 BUF_X2 _571_ (.A(b[6]),
    .Z(_013_));
 AND2_X1 _572_ (.A1(_002_),
    .A2(_013_),
    .ZN(_436_));
 NAND2_X1 _573_ (.A1(_003_),
    .A2(_012_),
    .ZN(_201_));
 INV_X1 _574_ (.A(_201_),
    .ZN(_442_));
 NAND2_X1 _575_ (.A1(_004_),
    .A2(_010_),
    .ZN(_202_));
 NAND2_X2 _576_ (.A1(_006_),
    .A2(_011_),
    .ZN(_205_));
 BUF_X16 _577_ (.A(net1),
    .Z(_014_));
 AND2_X1 _578_ (.A1(_003_),
    .A2(net47),
    .ZN(_453_));
 AND2_X1 _579_ (.A1(_004_),
    .A2(_012_),
    .ZN(_454_));
 AND2_X2 _580_ (.A1(_007_),
    .A2(_010_),
    .ZN(_237_));
 AND2_X2 _581_ (.A1(_008_),
    .A2(_009_),
    .ZN(_238_));
 AND2_X4 _582_ (.A1(_011_),
    .A2(_005_),
    .ZN(_239_));
 NAND2_X1 _583_ (.A1(_006_),
    .A2(_013_),
    .ZN(_247_));
 INV_X1 _584_ (.A(_247_),
    .ZN(_457_));
 BUF_X8 _585_ (.A(b[7]),
    .Z(_015_));
 INV_X4 _586_ (.A(_015_),
    .ZN(_016_));
 NOR2_X1 _587_ (.A1(_001_),
    .A2(_016_),
    .ZN(_460_));
 INV_X1 _588_ (.A(_267_),
    .ZN(_264_));
 NAND2_X1 _589_ (.A1(_004_),
    .A2(net47),
    .ZN(_274_));
 INV_X1 _590_ (.A(_274_),
    .ZN(_462_));
 AND2_X1 _591_ (.A1(_007_),
    .A2(_012_),
    .ZN(_268_));
 AND2_X2 _592_ (.A1(_009_),
    .A2(_010_),
    .ZN(_269_));
 AND2_X2 _593_ (.A1(_008_),
    .A2(_011_),
    .ZN(_270_));
 NAND2_X1 _594_ (.A1(_005_),
    .A2(_013_),
    .ZN(_278_));
 INV_X1 _595_ (.A(_278_),
    .ZN(_463_));
 NOR2_X1 _596_ (.A1(_006_),
    .A2(_016_),
    .ZN(_468_));
 NAND2_X4 _597_ (.A1(_007_),
    .A2(_014_),
    .ZN(_304_));
 INV_X2 _598_ (.A(_304_),
    .ZN(_343_));
 NAND2_X1 _599_ (.A1(_008_),
    .A2(_013_),
    .ZN(_309_));
 INV_X1 _600_ (.A(_309_),
    .ZN(_472_));
 INV_X2 _601_ (.A(_199_),
    .ZN(_194_));
 AND3_X1 _602_ (.A1(net5),
    .A2(_003_),
    .A3(net1),
    .ZN(_017_));
 OR2_X1 _603_ (.A1(_467_),
    .A2(_017_),
    .ZN(_320_));
 INV_X2 _604_ (.A(_320_),
    .ZN(_348_));
 NOR2_X1 _605_ (.A1(_005_),
    .A2(_016_),
    .ZN(_481_));
 AND2_X4 _606_ (.A1(_009_),
    .A2(_014_),
    .ZN(_344_));
 AND2_X1 _607_ (.A1(_011_),
    .A2(_012_),
    .ZN(_345_));
 NAND2_X1 _608_ (.A1(_010_),
    .A2(_013_),
    .ZN(_336_));
 INV_X1 _609_ (.A(_336_),
    .ZN(_491_));
 NOR2_X1 _610_ (.A1(_008_),
    .A2(_016_),
    .ZN(_498_));
 AND2_X4 _611_ (.A1(_014_),
    .A2(_011_),
    .ZN(_374_));
 AND2_X1 _612_ (.A1(_012_),
    .A2(_013_),
    .ZN(_365_));
 AND2_X1 _613_ (.A1(_010_),
    .A2(_015_),
    .ZN(_366_));
 NOR2_X1 _614_ (.A1(_010_),
    .A2(_016_),
    .ZN(_507_));
 AND2_X1 _615_ (.A1(_013_),
    .A2(net47),
    .ZN(_513_));
 AND2_X1 _616_ (.A1(_012_),
    .A2(_015_),
    .ZN(_512_));
 NOR2_X1 _617_ (.A1(_012_),
    .A2(_016_),
    .ZN(_520_));
 AND2_X1 _618_ (.A1(net47),
    .A2(_015_),
    .ZN(_525_));
 NAND2_X4 _619_ (.A1(_006_),
    .A2(_007_),
    .ZN(_165_));
 NAND2_X4 _620_ (.A1(_000_),
    .A2(_014_),
    .ZN(_200_));
 NAND2_X1 _621_ (.A1(_002_),
    .A2(_015_),
    .ZN(_212_));
 NAND2_X1 _622_ (.A1(_005_),
    .A2(_009_),
    .ZN(_206_));
 NAND2_X1 _623_ (.A1(_001_),
    .A2(_015_),
    .ZN(_246_));
 INV_X1 _624_ (.A(_455_),
    .ZN(_273_));
 NAND2_X1 _625_ (.A1(_010_),
    .A2(_011_),
    .ZN(_303_));
 NAND2_X1 _626_ (.A1(_008_),
    .A2(_015_),
    .ZN(_335_));
 NAND2_X1 _627_ (.A1(_001_),
    .A2(_003_),
    .ZN(_140_));
 NAND2_X2 _628_ (.A1(_001_),
    .A2(_009_),
    .ZN(_166_));
 NAND2_X1 _629_ (.A1(_006_),
    .A2(_009_),
    .ZN(_183_));
 INV_X1 _630_ (.A(_198_),
    .ZN(_193_));
 NAND2_X1 _631_ (.A1(_007_),
    .A2(_008_),
    .ZN(_207_));
 OR2_X1 _632_ (.A1(_002_),
    .A2(_016_),
    .ZN(_228_));
 NAND2_X1 _633_ (.A1(net5),
    .A2(_006_),
    .ZN(_141_));
 NAND2_X1 _634_ (.A1(_005_),
    .A2(_007_),
    .ZN(_184_));
 NAND2_X1 _635_ (.A1(_001_),
    .A2(_013_),
    .ZN(_213_));
 NAND2_X1 _636_ (.A1(_006_),
    .A2(_015_),
    .ZN(_280_));
 NAND2_X1 _637_ (.A1(_009_),
    .A2(_012_),
    .ZN(_305_));
 NAND2_X1 _638_ (.A1(_005_),
    .A2(_015_),
    .ZN(_310_));
 INV_X2 _639_ (.A(net16),
    .ZN(_243_));
 INV_X2 _640_ (.A(_257_),
    .ZN(_261_));
 INV_X1 _641_ (.A(_272_),
    .ZN(_275_));
 INV_X1 _642_ (.A(_290_),
    .ZN(_296_));
 INV_X1 _643_ (.A(_295_),
    .ZN(_298_));
 INV_X1 _644_ (.A(_316_),
    .ZN(_317_));
 INV_X1 _645_ (.A(_322_),
    .ZN(_328_));
 INV_X1 _646_ (.A(_326_),
    .ZN(_329_));
 INV_X1 _647_ (.A(_347_),
    .ZN(_349_));
 INV_X1 _648_ (.A(_356_),
    .ZN(_358_));
 INV_X2 _649_ (.A(_376_),
    .ZN(_377_));
 INV_X1 _650_ (.A(_383_),
    .ZN(_384_));
 INV_X1 _651_ (.A(_397_),
    .ZN(_398_));
 INV_X1 _652_ (.A(_407_),
    .ZN(_408_));
 INV_X1 _653_ (.A(_240_),
    .ZN(_279_));
 INV_X1 _654_ (.A(_256_),
    .ZN(_297_));
 INV_X1 _655_ (.A(_271_),
    .ZN(_308_));
 INV_X1 _656_ (.A(_289_),
    .ZN(_327_));
 INV_X1 _657_ (.A(_294_),
    .ZN(_332_));
 INV_X1 _658_ (.A(_315_),
    .ZN(_339_));
 INV_X1 _659_ (.A(_321_),
    .ZN(_357_));
 INV_X1 _660_ (.A(_325_),
    .ZN(_361_));
 INV_X1 _661_ (.A(_355_),
    .ZN(_387_));
 INV_X1 _662_ (.A(_382_),
    .ZN(_401_));
 INV_X1 _663_ (.A(_396_),
    .ZN(_411_));
 INV_X1 _664_ (.A(_151_),
    .ZN(_421_));
 INV_X1 _665_ (.A(_150_),
    .ZN(_427_));
 INV_X1 _666_ (.A(_158_),
    .ZN(_173_));
 INV_X1 _667_ (.A(_168_),
    .ZN(_435_));
 INV_X2 _668_ (.A(_230_),
    .ZN(_449_));
 INV_X1 _669_ (.A(_190_),
    .ZN(_218_));
 XOR2_X2 _670_ (.A(_000_),
    .B(_003_),
    .Z(_018_));
 AND2_X4 _671_ (.A1(_018_),
    .A2(_014_),
    .ZN(_458_));
 INV_X1 _672_ (.A(_319_),
    .ZN(_473_));
 INV_X2 _673_ (.A(_252_),
    .ZN(_477_));
 INV_X1 _674_ (.A(_301_),
    .ZN(_482_));
 INV_X1 _675_ (.A(_265_),
    .ZN(_486_));
 INV_X1 _676_ (.A(_342_),
    .ZN(_494_));
 INV_X1 _677_ (.A(_306_),
    .ZN(_352_));
 INV_X1 _678_ (.A(_333_),
    .ZN(_499_));
 INV_X1 _679_ (.A(_337_),
    .ZN(_369_));
 INV_X1 _680_ (.A(_362_),
    .ZN(_508_));
 INV_X1 _681_ (.A(_378_),
    .ZN(_517_));
 INV_X1 _682_ (.A(_388_),
    .ZN(_521_));
 NOR2_X1 _683_ (.A1(net47),
    .A2(_016_),
    .ZN(_530_));
 INV_X1 _684_ (.A(_413_),
    .ZN(_534_));
 INV_X1 _685_ (.A(_143_),
    .ZN(_418_));
 INV_X1 _686_ (.A(_159_),
    .ZN(_428_));
 INV_X2 _687_ (.A(_171_),
    .ZN(_174_));
 INV_X1 _688_ (.A(_191_),
    .ZN(_438_));
 INV_X1 _689_ (.A(_217_),
    .ZN(_220_));
 XNOR2_X2 _690_ (.A(_015_),
    .B(_200_),
    .ZN(_446_));
 INV_X1 _691_ (.A(_185_),
    .ZN(_443_));
 INV_X2 _692_ (.A(_233_),
    .ZN(_234_));
 INV_X1 _693_ (.A(_447_),
    .ZN(_019_));
 OAI21_X1 _694_ (.A(_019_),
    .B1(_200_),
    .B2(_016_),
    .ZN(_255_));
 INV_X2 _695_ (.A(_253_),
    .ZN(_464_));
 OR2_X2 _696_ (.A1(_459_),
    .A2(_017_),
    .ZN(_288_));
 INV_X2 _697_ (.A(_266_),
    .ZN(_469_));
 INV_X1 _698_ (.A(_276_),
    .ZN(_313_));
 INV_X1 _699_ (.A(_312_),
    .ZN(_314_));
 INV_X1 _700_ (.A(_285_),
    .ZN(_474_));
 INV_X2 _701_ (.A(_286_),
    .ZN(_478_));
 INV_X1 _702_ (.A(_334_),
    .ZN(_483_));
 INV_X2 _703_ (.A(_302_),
    .ZN(_487_));
 INV_X1 _704_ (.A(_338_),
    .ZN(_492_));
 INV_X1 _705_ (.A(_318_),
    .ZN(_495_));
 INV_X1 _706_ (.A(_363_),
    .ZN(_500_));
 INV_X1 _707_ (.A(_341_),
    .ZN(_503_));
 INV_X1 _708_ (.A(net25),
    .ZN(_506_));
 INV_X2 _709_ (.A(_389_),
    .ZN(_509_));
 INV_X1 _710_ (.A(_403_),
    .ZN(_522_));
 INV_X1 _711_ (.A(_402_),
    .ZN(_535_));
 INV_X1 _712_ (.A(_437_),
    .ZN(_189_));
 INV_X1 _713_ (.A(_448_),
    .ZN(_225_));
 INV_X2 _714_ (.A(net20),
    .ZN(_291_));
 INV_X1 _715_ (.A(_426_),
    .ZN(_157_));
 INV_X1 _716_ (.A(_197_),
    .ZN(_192_));
 INV_X1 _717_ (.A(_450_),
    .ZN(_231_));
 INV_X1 _718_ (.A(_456_),
    .ZN(_242_));
 INV_X1 _719_ (.A(_461_),
    .ZN(_258_));
 INV_X1 _720_ (.A(_493_),
    .ZN(_340_));
 AND2_X2 _721_ (.A1(net5),
    .A2(_002_),
    .ZN(net3));
 BUF_X4 _722_ (.A(net2),
    .Z(_020_));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 NAND2_X1 _724_ (.A1(net31),
    .A2(_465_),
    .ZN(_022_));
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 NAND3_X1 _726_ (.A1(_445_),
    .A2(_466_),
    .A3(_480_),
    .ZN(_024_));
 AOI21_X4 _727_ (.A(_440_),
    .B1(net43),
    .B2(_441_),
    .ZN(_025_));
 INV_X1 _728_ (.A(_444_),
    .ZN(_026_));
 NAND2_X1 _729_ (.A1(_466_),
    .A2(_480_),
    .ZN(_027_));
 OAI221_X2 _730_ (.A(_022_),
    .B1(_024_),
    .B2(_025_),
    .C1(_026_),
    .C2(_027_),
    .ZN(_028_));
 OAI21_X4 _731_ (.A(_476_),
    .B1(_028_),
    .B2(_479_),
    .ZN(_029_));
 OR3_X2 _732_ (.A1(_476_),
    .A2(_028_),
    .A3(_479_),
    .ZN(_030_));
 AOI21_X4 _733_ (.A(_020_),
    .B1(_030_),
    .B2(_029_),
    .ZN(_031_));
 INV_X1 _734_ (.A(_485_),
    .ZN(_032_));
 BUF_X4 _735_ (.A(_489_),
    .Z(_033_));
 NAND2_X4 _736_ (.A1(_033_),
    .A2(_470_),
    .ZN(_034_));
 BUF_X2 _737_ (.A(_471_),
    .Z(_035_));
 NAND3_X2 _738_ (.A1(_035_),
    .A2(_033_),
    .A3(net40),
    .ZN(_036_));
 INV_X1 _739_ (.A(_451_),
    .ZN(_037_));
 NAND2_X1 _740_ (.A1(_035_),
    .A2(_033_),
    .ZN(_038_));
 OAI221_X2 _741_ (.A(_034_),
    .B1(_036_),
    .B2(_025_),
    .C1(_037_),
    .C2(_038_),
    .ZN(_039_));
 NOR2_X4 _742_ (.A1(_488_),
    .A2(net35),
    .ZN(_040_));
 XNOR2_X2 _743_ (.A(_032_),
    .B(_040_),
    .ZN(_041_));
 AOI21_X4 _744_ (.A(_031_),
    .B1(_041_),
    .B2(_020_),
    .ZN(net4));
 BUF_X2 _745_ (.A(_502_),
    .Z(_042_));
 INV_X1 _746_ (.A(_484_),
    .ZN(_043_));
 AND2_X2 _747_ (.A1(_035_),
    .A2(_033_),
    .ZN(_044_));
 INV_X2 _748_ (.A(net39),
    .ZN(_045_));
 OAI21_X4 _749_ (.A(_037_),
    .B1(net49),
    .B2(_045_),
    .ZN(_046_));
 AOI221_X2 _750_ (.A(_488_),
    .B1(_044_),
    .B2(_046_),
    .C1(_470_),
    .C2(_033_),
    .ZN(_047_));
 OAI21_X2 _751_ (.A(_043_),
    .B1(_047_),
    .B2(_032_),
    .ZN(_048_));
 XOR2_X1 _752_ (.A(_048_),
    .B(_042_),
    .Z(_049_));
 BUF_X1 _753_ (.A(_497_),
    .Z(_050_));
 INV_X1 _754_ (.A(_475_),
    .ZN(_051_));
 OAI21_X4 _755_ (.A(net32),
    .B1(net33),
    .B2(_465_),
    .ZN(_052_));
 NOR2_X1 _756_ (.A1(_444_),
    .A2(_465_),
    .ZN(_053_));
 INV_X1 _757_ (.A(net44),
    .ZN(_054_));
 OR2_X2 _758_ (.A1(_054_),
    .A2(_195_),
    .ZN(_055_));
 AOI21_X4 _759_ (.A(_052_),
    .B1(_055_),
    .B2(_053_),
    .ZN(_056_));
 OAI21_X2 _760_ (.A(_476_),
    .B1(_056_),
    .B2(_479_),
    .ZN(_057_));
 NAND2_X1 _761_ (.A1(_057_),
    .A2(_051_),
    .ZN(_058_));
 XOR2_X1 _762_ (.A(_058_),
    .B(_050_),
    .Z(_059_));
 INV_X4 _763_ (.A(_020_),
    .ZN(_060_));
 MUX2_X2 _764_ (.A(_049_),
    .B(_059_),
    .S(_060_),
    .Z(net6));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 OAI21_X4 _766_ (.A(_043_),
    .B1(_040_),
    .B2(_032_),
    .ZN(_062_));
 AOI21_X2 _767_ (.A(_501_),
    .B1(_062_),
    .B2(_042_),
    .ZN(_063_));
 XNOR2_X1 _768_ (.A(_063_),
    .B(net23),
    .ZN(_064_));
 BUF_X1 _769_ (.A(_505_),
    .Z(_065_));
 NAND2_X1 _770_ (.A1(_051_),
    .A2(_029_),
    .ZN(_066_));
 AOI21_X1 _771_ (.A(_496_),
    .B1(_066_),
    .B2(_050_),
    .ZN(_067_));
 XNOR2_X1 _772_ (.A(_065_),
    .B(_067_),
    .ZN(_068_));
 MUX2_X2 _773_ (.A(_064_),
    .B(_068_),
    .S(_060_),
    .Z(net7));
 BUF_X1 _774_ (.A(_516_),
    .Z(_069_));
 AOI21_X1 _775_ (.A(_504_),
    .B1(_496_),
    .B2(_065_),
    .ZN(_070_));
 NAND2_X1 _776_ (.A1(_050_),
    .A2(_065_),
    .ZN(_071_));
 NOR2_X1 _777_ (.A1(_476_),
    .A2(_475_),
    .ZN(_072_));
 OAI21_X1 _778_ (.A(_070_),
    .B1(_071_),
    .B2(_072_),
    .ZN(_073_));
 INV_X1 _779_ (.A(_479_),
    .ZN(_074_));
 NAND3_X1 _780_ (.A1(_051_),
    .A2(_074_),
    .A3(_070_),
    .ZN(_075_));
 OAI21_X4 _781_ (.A(_073_),
    .B1(net41),
    .B2(_075_),
    .ZN(_076_));
 XNOR2_X2 _782_ (.A(_076_),
    .B(_069_),
    .ZN(_077_));
 NAND2_X2 _783_ (.A1(_077_),
    .A2(_060_),
    .ZN(_078_));
 BUF_X8 clone5 (.A(b[0]),
    .Z(net5));
 NOR2_X1 _785_ (.A1(_501_),
    .A2(_510_),
    .ZN(_080_));
 OAI21_X1 _786_ (.A(_042_),
    .B1(_484_),
    .B2(_485_),
    .ZN(_081_));
 INV_X1 _787_ (.A(_488_),
    .ZN(_082_));
 NAND3_X2 _788_ (.A1(_043_),
    .A2(_082_),
    .A3(_034_),
    .ZN(_083_));
 AOI21_X4 _789_ (.A(_083_),
    .B1(_046_),
    .B2(_044_),
    .ZN(_084_));
 OAI21_X2 _790_ (.A(_080_),
    .B1(_084_),
    .B2(_081_),
    .ZN(_085_));
 OAI21_X2 _791_ (.A(_085_),
    .B1(_510_),
    .B2(net21),
    .ZN(_086_));
 XOR2_X2 _792_ (.A(_086_),
    .B(net46),
    .Z(_087_));
 OAI21_X4 _793_ (.A(_078_),
    .B1(_087_),
    .B2(_060_),
    .ZN(net8));
 INV_X1 _794_ (.A(_537_),
    .ZN(_088_));
 NOR3_X1 _795_ (.A1(_524_),
    .A2(_088_),
    .A3(_523_),
    .ZN(_089_));
 INV_X1 _796_ (.A(_523_),
    .ZN(_090_));
 NOR2_X1 _797_ (.A1(_537_),
    .A2(_090_),
    .ZN(_091_));
 OAI21_X1 _798_ (.A(_020_),
    .B1(_089_),
    .B2(_091_),
    .ZN(_092_));
 INV_X1 _799_ (.A(_529_),
    .ZN(_093_));
 NAND2_X1 _800_ (.A1(_093_),
    .A2(_515_),
    .ZN(_094_));
 OR3_X1 _801_ (.A1(_020_),
    .A2(_093_),
    .A3(_515_),
    .ZN(_095_));
 OAI221_X2 _802_ (.A(_092_),
    .B1(_094_),
    .B2(_020_),
    .C1(_069_),
    .C2(_095_),
    .ZN(_096_));
 OR2_X2 _803_ (.A1(_039_),
    .A2(_488_),
    .ZN(_097_));
 AND3_X1 _804_ (.A1(_485_),
    .A2(_042_),
    .A3(net21),
    .ZN(_098_));
 AOI21_X1 _805_ (.A(_501_),
    .B1(_484_),
    .B2(_042_),
    .ZN(_099_));
 INV_X1 _806_ (.A(_099_),
    .ZN(_100_));
 AOI221_X2 _807_ (.A(_510_),
    .B1(_098_),
    .B2(_097_),
    .C1(_100_),
    .C2(net21),
    .ZN(_101_));
 AND2_X1 _808_ (.A1(net2),
    .A2(net45),
    .ZN(_102_));
 AOI21_X2 _809_ (.A(_101_),
    .B1(_102_),
    .B2(_088_),
    .ZN(_103_));
 NAND3_X1 _810_ (.A1(_020_),
    .A2(_537_),
    .A3(_090_),
    .ZN(_104_));
 AOI21_X2 _811_ (.A(_103_),
    .B1(_104_),
    .B2(_101_),
    .ZN(_105_));
 AOI21_X1 _812_ (.A(_496_),
    .B1(_475_),
    .B2(_050_),
    .ZN(_106_));
 INV_X1 _813_ (.A(_106_),
    .ZN(_107_));
 AOI21_X1 _814_ (.A(_504_),
    .B1(_107_),
    .B2(_065_),
    .ZN(_108_));
 OAI21_X1 _815_ (.A(_108_),
    .B1(_071_),
    .B2(_029_),
    .ZN(_109_));
 NAND4_X1 _816_ (.A1(_060_),
    .A2(_069_),
    .A3(_093_),
    .A4(_109_),
    .ZN(_110_));
 OAI21_X1 _817_ (.A(_110_),
    .B1(_109_),
    .B2(_095_),
    .ZN(_111_));
 OR3_X4 _818_ (.A1(_105_),
    .A2(_096_),
    .A3(_111_),
    .ZN(net9));
 OAI21_X4 _819_ (.A(_524_),
    .B1(_510_),
    .B2(net22),
    .ZN(_112_));
 AOI21_X4 _820_ (.A(_088_),
    .B1(_090_),
    .B2(_112_),
    .ZN(_113_));
 OR2_X4 _821_ (.A1(_536_),
    .A2(_113_),
    .ZN(_114_));
 NOR4_X2 _822_ (.A1(_501_),
    .A2(_510_),
    .A3(_523_),
    .A4(_536_),
    .ZN(_115_));
 OAI21_X2 _823_ (.A(_115_),
    .B1(_081_),
    .B2(_084_),
    .ZN(_116_));
 XNOR2_X1 _824_ (.A(_406_),
    .B(_533_),
    .ZN(_117_));
 XNOR2_X1 _825_ (.A(_409_),
    .B(_412_),
    .ZN(_118_));
 XNOR2_X1 _826_ (.A(_117_),
    .B(_118_),
    .ZN(_119_));
 XNOR2_X1 _827_ (.A(_531_),
    .B(_519_),
    .ZN(_120_));
 XNOR2_X1 _828_ (.A(_119_),
    .B(_120_),
    .ZN(_121_));
 AND3_X4 _829_ (.A1(_114_),
    .A2(_116_),
    .A3(_121_),
    .ZN(_122_));
 AOI21_X4 _830_ (.A(_121_),
    .B1(_114_),
    .B2(_116_),
    .ZN(_123_));
 OAI21_X4 _831_ (.A(_020_),
    .B1(_123_),
    .B2(_122_),
    .ZN(_124_));
 AOI21_X1 _832_ (.A(_528_),
    .B1(_515_),
    .B2(_529_),
    .ZN(_125_));
 NAND2_X1 _833_ (.A1(_069_),
    .A2(_529_),
    .ZN(_126_));
 OAI21_X4 _834_ (.A(_125_),
    .B1(_076_),
    .B2(_126_),
    .ZN(_127_));
 XNOR2_X2 _835_ (.A(_127_),
    .B(_526_),
    .ZN(_128_));
 OAI21_X4 _836_ (.A(_124_),
    .B1(_020_),
    .B2(_128_),
    .ZN(net10));
 BUF_X2 _837_ (.A(_417_),
    .Z(net11));
 BUF_X2 _838_ (.A(_420_),
    .Z(net12));
 BUF_X2 _839_ (.A(_423_),
    .Z(net13));
 BUF_X2 _840_ (.A(_432_),
    .Z(net14));
 BUF_X2 _841_ (.A(_434_),
    .Z(net15));
 BUF_X2 rebuffer7 (.A(_241_),
    .Z(net16));
 MUX2_X1 _843_ (.A(net50),
    .B(net40),
    .S(_020_),
    .Z(_129_));
 XNOR2_X2 _844_ (.A(_129_),
    .B(net49),
    .ZN(net17));
 OAI21_X1 _845_ (.A(_037_),
    .B1(_025_),
    .B2(_045_),
    .ZN(_130_));
 XOR2_X1 _846_ (.A(_035_),
    .B(_130_),
    .Z(_131_));
 OAI21_X1 _847_ (.A(_026_),
    .B1(_025_),
    .B2(_054_),
    .ZN(_132_));
 XOR2_X1 _848_ (.A(net34),
    .B(_132_),
    .Z(_133_));
 MUX2_X2 _849_ (.A(_131_),
    .B(_133_),
    .S(_060_),
    .Z(net18));
 AOI21_X1 _850_ (.A(_470_),
    .B1(_046_),
    .B2(_035_),
    .ZN(_134_));
 XNOR2_X1 _851_ (.A(_033_),
    .B(_134_),
    .ZN(_135_));
 NAND2_X2 _852_ (.A1(_055_),
    .A2(_026_),
    .ZN(_136_));
 AOI21_X2 _853_ (.A(_465_),
    .B1(_136_),
    .B2(net34),
    .ZN(_137_));
 XNOR2_X1 _854_ (.A(_137_),
    .B(net42),
    .ZN(_138_));
 MUX2_X2 _855_ (.A(_135_),
    .B(_138_),
    .S(_060_),
    .Z(net19));
 FA_X1 _856_ (.A(_139_),
    .B(_140_),
    .CI(_141_),
    .CO(_142_),
    .S(_143_));
 FA_X1 _857_ (.A(_144_),
    .B(_145_),
    .CI(_146_),
    .CO(_147_),
    .S(_148_));
 FA_X1 _858_ (.A(_149_),
    .B(_142_),
    .CI(_148_),
    .CO(_150_),
    .S(_151_));
 FA_X1 _859_ (.A(_152_),
    .B(_153_),
    .CI(_154_),
    .CO(_155_),
    .S(_156_));
 FA_X1 _860_ (.A(_156_),
    .B(_147_),
    .CI(_157_),
    .CO(_158_),
    .S(_159_));
 FA_X1 _861_ (.A(_160_),
    .B(_161_),
    .CI(_162_),
    .CO(_163_),
    .S(_164_));
 FA_X1 _862_ (.A(_165_),
    .B(_166_),
    .CI(_167_),
    .CO(_168_),
    .S(_169_));
 FA_X1 _863_ (.A(_164_),
    .B(_169_),
    .CI(_155_),
    .CO(_170_),
    .S(_171_));
 FA_X1 _864_ (.A(_172_),
    .B(_173_),
    .CI(_174_),
    .CO(_175_),
    .S(_176_));
 FA_X1 _865_ (.A(_177_),
    .B(_178_),
    .CI(_179_),
    .CO(_180_),
    .S(_181_));
 FA_X1 _866_ (.A(_182_),
    .B(_183_),
    .CI(_184_),
    .CO(_185_),
    .S(_186_));
 FA_X1 _867_ (.A(_181_),
    .B(_186_),
    .CI(_163_),
    .CO(_187_),
    .S(_188_));
 FA_X1 _868_ (.A(_189_),
    .B(_170_),
    .CI(_188_),
    .CO(_190_),
    .S(_191_));
 FA_X1 _869_ (.A(_194_),
    .B(_193_),
    .CI(_192_),
    .CO(_195_),
    .S(_196_));
 FA_X1 _870_ (.A(_202_),
    .B(_201_),
    .CI(_200_),
    .CO(_203_),
    .S(_204_));
 FA_X1 _871_ (.A(_205_),
    .B(_206_),
    .CI(_207_),
    .CO(_208_),
    .S(_209_));
 FA_X1 _872_ (.A(_180_),
    .B(_204_),
    .CI(_209_),
    .CO(_210_),
    .S(_211_));
 FA_X1 _873_ (.A(_212_),
    .B(_213_),
    .CI(_185_),
    .CO(_214_),
    .S(_215_));
 FA_X1 _874_ (.A(_215_),
    .B(_187_),
    .CI(_211_),
    .CO(_216_),
    .S(_217_));
 FA_X1 _875_ (.A(_218_),
    .B(_219_),
    .CI(_220_),
    .CO(_221_),
    .S(_222_));
 FA_X1 _876_ (.A(_206_),
    .B(_202_),
    .CI(_207_),
    .CO(_223_),
    .S(_224_));
 FA_X1 _877_ (.A(_180_),
    .B(_224_),
    .CI(_225_),
    .CO(_226_),
    .S(_227_));
 FA_X1 _878_ (.A(_205_),
    .B(_228_),
    .CI(_213_),
    .CO(_229_),
    .S(_230_));
 FA_X1 _879_ (.A(_227_),
    .B(_187_),
    .CI(_231_),
    .CO(_232_),
    .S(_233_));
 FA_X1 _880_ (.A(_218_),
    .B(_219_),
    .CI(_234_),
    .CO(_235_),
    .S(_236_));
 FA_X1 _881_ (.A(_238_),
    .B(_239_),
    .CI(_237_),
    .CO(_240_),
    .S(_241_));
 FA_X1 _882_ (.A(_203_),
    .B(_242_),
    .CI(_243_),
    .CO(_244_),
    .S(_245_));
 FA_X1 _883_ (.A(_246_),
    .B(_208_),
    .CI(_247_),
    .CO(_248_),
    .S(_249_));
 FA_X1 _884_ (.A(_210_),
    .B(_245_),
    .CI(_249_),
    .CO(_250_),
    .S(_251_));
 FA_X1 _885_ (.A(_214_),
    .B(_251_),
    .CI(_216_),
    .CO(_252_),
    .S(_253_));
 FA_X1 _886_ (.A(_254_),
    .B(_255_),
    .CI(_241_),
    .CO(_256_),
    .S(_257_));
 FA_X1 _887_ (.A(_258_),
    .B(_223_),
    .CI(_229_),
    .CO(_259_),
    .S(_260_));
 FA_X1 _888_ (.A(_226_),
    .B(_261_),
    .CI(_260_),
    .CO(_262_),
    .S(_263_));
 FA_X1 _889_ (.A(_264_),
    .B(_232_),
    .CI(_263_),
    .CO(_265_),
    .S(_266_));
 FA_X1 _890_ (.A(_270_),
    .B(_269_),
    .CI(_268_),
    .CO(_271_),
    .S(_272_));
 FA_X1 _891_ (.A(_273_),
    .B(_274_),
    .CI(_275_),
    .CO(_276_),
    .S(_277_));
 FA_X1 _892_ (.A(_278_),
    .B(_279_),
    .CI(_280_),
    .CO(_281_),
    .S(_282_));
 FA_X1 _893_ (.A(_244_),
    .B(_282_),
    .CI(_277_),
    .CO(_283_),
    .S(_284_));
 FA_X1 _894_ (.A(_250_),
    .B(_248_),
    .CI(_284_),
    .CO(_285_),
    .S(_286_));
 FA_X1 _895_ (.A(_288_),
    .B(_272_),
    .CI(_287_),
    .CO(_289_),
    .S(_290_));
 FA_X1 _896_ (.A(_240_),
    .B(_292_),
    .CI(_293_),
    .CO(_294_),
    .S(_295_));
 FA_X1 _897_ (.A(_298_),
    .B(_297_),
    .CI(_296_),
    .CO(_299_),
    .S(_300_));
 FA_X1 _898_ (.A(_262_),
    .B(_259_),
    .CI(_300_),
    .CO(_301_),
    .S(_302_));
 FA_X1 _899_ (.A(_303_),
    .B(_304_),
    .CI(_305_),
    .CO(_306_),
    .S(_307_));
 FA_X1 _900_ (.A(_308_),
    .B(_309_),
    .CI(_310_),
    .CO(_311_),
    .S(_312_));
 FA_X1 _901_ (.A(_307_),
    .B(_313_),
    .CI(_314_),
    .CO(_315_),
    .S(_316_));
 FA_X1 _902_ (.A(_283_),
    .B(_317_),
    .CI(_281_),
    .CO(_318_),
    .S(_319_));
 FA_X1 _903_ (.A(_307_),
    .B(net20),
    .CI(_320_),
    .CO(_321_),
    .S(_322_));
 FA_X1 _904_ (.A(_271_),
    .B(_323_),
    .CI(_324_),
    .CO(_325_),
    .S(_326_));
 FA_X1 _905_ (.A(_327_),
    .B(_328_),
    .CI(_329_),
    .CO(_330_),
    .S(_331_));
 FA_X1 _906_ (.A(_331_),
    .B(_299_),
    .CI(_332_),
    .CO(_333_),
    .S(_334_));
 FA_X1 _907_ (.A(_335_),
    .B(_306_),
    .CI(_336_),
    .CO(_337_),
    .S(_338_));
 FA_X1 _908_ (.A(_311_),
    .B(_339_),
    .CI(_340_),
    .CO(_341_),
    .S(_342_));
 FA_X1 _909_ (.A(_343_),
    .B(_344_),
    .CI(_345_),
    .CO(_346_),
    .S(_347_));
 FA_X1 _910_ (.A(_291_),
    .B(_348_),
    .CI(_349_),
    .CO(_350_),
    .S(_351_));
 FA_X1 _911_ (.A(_352_),
    .B(_353_),
    .CI(_354_),
    .CO(_355_),
    .S(_356_));
 FA_X1 _912_ (.A(_351_),
    .B(_357_),
    .CI(_358_),
    .CO(_359_),
    .S(_360_));
 FA_X1 _913_ (.A(_361_),
    .B(_330_),
    .CI(_360_),
    .CO(_362_),
    .S(_363_));
 FA_X1 _914_ (.A(_364_),
    .B(_365_),
    .CI(_366_),
    .CO(_367_),
    .S(_368_));
 FA_X1 _915_ (.A(_369_),
    .B(_370_),
    .CI(_371_),
    .CO(_372_),
    .S(_373_));
 FA_X1 _916_ (.A(_343_),
    .B(_374_),
    .CI(_344_),
    .CO(_375_),
    .S(_376_));
 FA_X1 _917_ (.A(_348_),
    .B(_377_),
    .CI(_291_),
    .CO(_378_),
    .S(_379_));
 FA_X1 _918_ (.A(_380_),
    .B(_381_),
    .CI(_346_),
    .CO(_382_),
    .S(_383_));
 FA_X1 _919_ (.A(_384_),
    .B(_350_),
    .CI(_379_),
    .CO(_385_),
    .S(_386_));
 FA_X1 _920_ (.A(_387_),
    .B(_359_),
    .CI(_386_),
    .CO(_388_),
    .S(_389_));
 FA_X1 _921_ (.A(_390_),
    .B(_391_),
    .CI(_367_),
    .CO(_392_),
    .S(_393_));
 FA_X1 _922_ (.A(_394_),
    .B(_375_),
    .CI(_395_),
    .CO(_396_),
    .S(_397_));
 FA_X1 _923_ (.A(_378_),
    .B(net24),
    .CI(_398_),
    .CO(_399_),
    .S(_400_));
 FA_X1 _924_ (.A(_385_),
    .B(_401_),
    .CI(_400_),
    .CO(_402_),
    .S(_403_));
 FA_X1 _925_ (.A(_375_),
    .B(_404_),
    .CI(_405_),
    .CO(_406_),
    .S(_407_));
 FA_X1 _926_ (.A(_378_),
    .B(_408_),
    .CI(net24),
    .CO(_409_),
    .S(_410_));
 FA_X1 _927_ (.A(_411_),
    .B(_410_),
    .CI(_399_),
    .CO(_412_),
    .S(_413_));
 HA_X1 _928_ (.A(_414_),
    .B(_415_),
    .CO(_416_),
    .S(_417_));
 HA_X1 _929_ (.A(_416_),
    .B(_418_),
    .CO(_419_),
    .S(_420_));
 HA_X1 _930_ (.A(_421_),
    .B(_419_),
    .CO(_422_),
    .S(_423_));
 HA_X1 _931_ (.A(_424_),
    .B(_425_),
    .CO(_172_),
    .S(_426_));
 HA_X1 _932_ (.A(_427_),
    .B(_428_),
    .CO(_429_),
    .S(_430_));
 HA_X1 _933_ (.A(_430_),
    .B(_422_),
    .CO(_431_),
    .S(_432_));
 HA_X1 _934_ (.A(_429_),
    .B(_176_),
    .CO(_198_),
    .S(_433_));
 HA_X1 _935_ (.A(_433_),
    .B(_431_),
    .CO(_199_),
    .S(_434_));
 HA_X1 _936_ (.A(_435_),
    .B(_436_),
    .CO(_219_),
    .S(_437_));
 HA_X1 _937_ (.A(_175_),
    .B(_438_),
    .CO(_439_),
    .S(_197_));
 HA_X1 _938_ (.A(_197_),
    .B(_198_),
    .CO(_440_),
    .S(_441_));
 HA_X1 _939_ (.A(_439_),
    .B(_222_),
    .CO(_444_),
    .S(_445_));
 HA_X1 _940_ (.A(_442_),
    .B(_446_),
    .CO(_447_),
    .S(_448_));
 HA_X1 _941_ (.A(_449_),
    .B(_443_),
    .CO(_267_),
    .S(_450_));
 HA_X1 _942_ (.A(_236_),
    .B(_439_),
    .CO(_451_),
    .S(_452_));
 HA_X1 _943_ (.A(_453_),
    .B(_454_),
    .CO(_455_),
    .S(_456_));
 HA_X1 _944_ (.A(_454_),
    .B(_458_),
    .CO(_459_),
    .S(_254_));
 HA_X1 _945_ (.A(_457_),
    .B(_460_),
    .CO(_293_),
    .S(_461_));
 HA_X1 _946_ (.A(_221_),
    .B(_464_),
    .CO(_465_),
    .S(_466_));
 HA_X1 _947_ (.A(_458_),
    .B(_462_),
    .CO(_467_),
    .S(_287_));
 HA_X1 _948_ (.A(_463_),
    .B(_468_),
    .CO(_323_),
    .S(_292_));
 HA_X1 _949_ (.A(_235_),
    .B(_469_),
    .CO(_470_),
    .S(_471_));
 HA_X1 _950_ (.A(_473_),
    .B(_474_),
    .CO(_475_),
    .S(_476_));
 HA_X1 _951_ (.A(_478_),
    .B(_477_),
    .CO(_479_),
    .S(_480_));
 HA_X1 _952_ (.A(_472_),
    .B(_481_),
    .CO(_354_),
    .S(_324_));
 HA_X1 _953_ (.A(_482_),
    .B(_483_),
    .CO(_484_),
    .S(_485_));
 HA_X1 _954_ (.A(_486_),
    .B(_487_),
    .CO(_488_),
    .S(_489_));
 HA_X1 _955_ (.A(_344_),
    .B(_345_),
    .CO(_364_),
    .S(_490_));
 HA_X1 _956_ (.A(_490_),
    .B(_492_),
    .CO(_371_),
    .S(_493_));
 HA_X1 _957_ (.A(_494_),
    .B(_495_),
    .CO(_496_),
    .S(_497_));
 HA_X1 _958_ (.A(_491_),
    .B(_498_),
    .CO(_380_),
    .S(_353_));
 HA_X1 _959_ (.A(_499_),
    .B(_500_),
    .CO(_501_),
    .S(_502_));
 HA_X1 _960_ (.A(_368_),
    .B(net48),
    .CO(_390_),
    .S(_370_));
 HA_X1 _961_ (.A(_373_),
    .B(_503_),
    .CO(_504_),
    .S(_505_));
 HA_X1 _962_ (.A(_507_),
    .B(_365_),
    .CO(_395_),
    .S(_381_));
 HA_X1 _963_ (.A(_508_),
    .B(_509_),
    .CO(_510_),
    .S(_511_));
 HA_X1 _964_ (.A(_512_),
    .B(_513_),
    .CO(_514_),
    .S(_391_));
 HA_X1 _965_ (.A(_393_),
    .B(_372_),
    .CO(_515_),
    .S(_516_));
 HA_X1 _966_ (.A(_517_),
    .B(_506_),
    .CO(_518_),
    .S(_519_));
 HA_X1 _967_ (.A(_520_),
    .B(_513_),
    .CO(_405_),
    .S(_394_));
 HA_X1 _968_ (.A(_521_),
    .B(_522_),
    .CO(_523_),
    .S(_524_));
 HA_X1 _969_ (.A(_514_),
    .B(_525_),
    .CO(_526_),
    .S(_527_));
 HA_X1 _970_ (.A(_527_),
    .B(_392_),
    .CO(_528_),
    .S(_529_));
 HA_X1 _971_ (.A(_530_),
    .B(_513_),
    .CO(_531_),
    .S(_404_));
 HA_X1 _972_ (.A(_375_),
    .B(_404_),
    .CO(_532_),
    .S(_533_));
 HA_X1 _973_ (.A(_534_),
    .B(_535_),
    .CO(_536_),
    .S(_537_));
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Left_513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_901 ();
 BUF_X32 input1 (.A(a[7]),
    .Z(net1));
 CLKBUF_X3 input2 (.A(sign_mode),
    .Z(net2));
 BUF_X1 output3 (.A(net3),
    .Z(product[0]));
 BUF_X1 output4 (.A(net4),
    .Z(product[10]));
 BUF_X2 output5 (.A(net6),
    .Z(product[11]));
 BUF_X2 output6 (.A(net7),
    .Z(product[12]));
 BUF_X1 output7 (.A(net8),
    .Z(product[13]));
 BUF_X1 output8 (.A(net9),
    .Z(product[14]));
 BUF_X2 output9 (.A(net10),
    .Z(product[15]));
 BUF_X1 output10 (.A(net11),
    .Z(product[1]));
 BUF_X1 output11 (.A(net12),
    .Z(product[2]));
 BUF_X1 output12 (.A(net13),
    .Z(product[3]));
 BUF_X1 output13 (.A(net14),
    .Z(product[4]));
 BUF_X1 output14 (.A(net15),
    .Z(product[5]));
 BUF_X2 output15 (.A(_196_),
    .Z(product[6]));
 BUF_X1 output16 (.A(net17),
    .Z(product[7]));
 BUF_X2 output17 (.A(net18),
    .Z(product[8]));
 BUF_X1 output18 (.A(net19),
    .Z(product[9]));
 BUF_X2 rebuffer1 (.A(_287_),
    .Z(net20));
 BUF_X4 rebuffer2 (.A(_511_),
    .Z(net21));
 BUF_X4 rebuffer3 (.A(net21),
    .Z(net22));
 BUF_X1 rebuffer4 (.A(net21),
    .Z(net23));
 BUF_X2 rebuffer5 (.A(_379_),
    .Z(net24));
 BUF_X1 rebuffer6 (.A(net24),
    .Z(net25));
 BUF_X2 rebuffer12 (.A(_480_),
    .Z(net31));
 BUF_X4 rebuffer13 (.A(net31),
    .Z(net32));
 BUF_X2 rebuffer14 (.A(_466_),
    .Z(net33));
 BUF_X4 rebuffer15 (.A(net33),
    .Z(net34));
 BUF_X2 rebuffer16 (.A(_039_),
    .Z(net35));
 BUF_X1 rebuffer20 (.A(_452_),
    .Z(net39));
 BUF_X2 rebuffer21 (.A(_452_),
    .Z(net40));
 BUF_X4 rebuffer22 (.A(_056_),
    .Z(net41));
 BUF_X1 rebuffer23 (.A(_480_),
    .Z(net42));
 BUF_X1 rebuffer24 (.A(_199_),
    .Z(net43));
 BUF_X1 rebuffer26 (.A(_524_),
    .Z(net45));
 BUF_X1 rebuffer27 (.A(net45),
    .Z(net46));
 BUF_X4 clone28 (.A(net1),
    .Z(net47));
 BUF_X1 rebuffer29 (.A(_374_),
    .Z(net48));
 BUF_X2 rebuffer30 (.A(_195_),
    .Z(net49));
 BUF_X1 rebuffer17 (.A(_445_),
    .Z(net44));
 BUF_X1 rebuffer18 (.A(net44),
    .Z(net50));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X32 FILLER_0_856 ();
 FILLCELL_X32 FILLER_0_888 ();
 FILLCELL_X32 FILLER_0_920 ();
 FILLCELL_X16 FILLER_0_952 ();
 FILLCELL_X4 FILLER_0_968 ();
 FILLCELL_X2 FILLER_0_972 ();
 FILLCELL_X1 FILLER_0_974 ();
 FILLCELL_X32 FILLER_0_1024 ();
 FILLCELL_X32 FILLER_0_1056 ();
 FILLCELL_X32 FILLER_0_1088 ();
 FILLCELL_X32 FILLER_0_1120 ();
 FILLCELL_X32 FILLER_0_1152 ();
 FILLCELL_X32 FILLER_0_1184 ();
 FILLCELL_X32 FILLER_0_1216 ();
 FILLCELL_X8 FILLER_0_1248 ();
 FILLCELL_X4 FILLER_0_1256 ();
 FILLCELL_X2 FILLER_0_1260 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X32 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_0_1679 ();
 FILLCELL_X32 FILLER_0_1711 ();
 FILLCELL_X32 FILLER_0_1743 ();
 FILLCELL_X32 FILLER_0_1775 ();
 FILLCELL_X32 FILLER_0_1807 ();
 FILLCELL_X32 FILLER_0_1839 ();
 FILLCELL_X16 FILLER_0_1871 ();
 FILLCELL_X4 FILLER_0_1887 ();
 FILLCELL_X2 FILLER_0_1891 ();
 FILLCELL_X2 FILLER_0_1894 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X32 FILLER_1_801 ();
 FILLCELL_X32 FILLER_1_833 ();
 FILLCELL_X32 FILLER_1_865 ();
 FILLCELL_X32 FILLER_1_897 ();
 FILLCELL_X32 FILLER_1_929 ();
 FILLCELL_X32 FILLER_1_961 ();
 FILLCELL_X32 FILLER_1_993 ();
 FILLCELL_X32 FILLER_1_1025 ();
 FILLCELL_X32 FILLER_1_1057 ();
 FILLCELL_X32 FILLER_1_1089 ();
 FILLCELL_X32 FILLER_1_1121 ();
 FILLCELL_X32 FILLER_1_1153 ();
 FILLCELL_X32 FILLER_1_1185 ();
 FILLCELL_X32 FILLER_1_1217 ();
 FILLCELL_X8 FILLER_1_1249 ();
 FILLCELL_X4 FILLER_1_1257 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X32 FILLER_1_1648 ();
 FILLCELL_X32 FILLER_1_1680 ();
 FILLCELL_X32 FILLER_1_1712 ();
 FILLCELL_X32 FILLER_1_1744 ();
 FILLCELL_X32 FILLER_1_1776 ();
 FILLCELL_X32 FILLER_1_1808 ();
 FILLCELL_X32 FILLER_1_1840 ();
 FILLCELL_X16 FILLER_1_1872 ();
 FILLCELL_X8 FILLER_1_1888 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X32 FILLER_2_952 ();
 FILLCELL_X32 FILLER_2_984 ();
 FILLCELL_X32 FILLER_2_1016 ();
 FILLCELL_X32 FILLER_2_1048 ();
 FILLCELL_X32 FILLER_2_1080 ();
 FILLCELL_X32 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1144 ();
 FILLCELL_X32 FILLER_2_1176 ();
 FILLCELL_X32 FILLER_2_1208 ();
 FILLCELL_X32 FILLER_2_1240 ();
 FILLCELL_X32 FILLER_2_1272 ();
 FILLCELL_X32 FILLER_2_1304 ();
 FILLCELL_X32 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1368 ();
 FILLCELL_X32 FILLER_2_1400 ();
 FILLCELL_X32 FILLER_2_1432 ();
 FILLCELL_X32 FILLER_2_1464 ();
 FILLCELL_X32 FILLER_2_1496 ();
 FILLCELL_X32 FILLER_2_1528 ();
 FILLCELL_X32 FILLER_2_1560 ();
 FILLCELL_X32 FILLER_2_1592 ();
 FILLCELL_X32 FILLER_2_1624 ();
 FILLCELL_X32 FILLER_2_1656 ();
 FILLCELL_X32 FILLER_2_1688 ();
 FILLCELL_X32 FILLER_2_1720 ();
 FILLCELL_X32 FILLER_2_1752 ();
 FILLCELL_X32 FILLER_2_1784 ();
 FILLCELL_X32 FILLER_2_1816 ();
 FILLCELL_X32 FILLER_2_1848 ();
 FILLCELL_X8 FILLER_2_1880 ();
 FILLCELL_X4 FILLER_2_1888 ();
 FILLCELL_X2 FILLER_2_1892 ();
 FILLCELL_X1 FILLER_2_1895 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X32 FILLER_3_1648 ();
 FILLCELL_X32 FILLER_3_1680 ();
 FILLCELL_X32 FILLER_3_1712 ();
 FILLCELL_X32 FILLER_3_1744 ();
 FILLCELL_X32 FILLER_3_1776 ();
 FILLCELL_X32 FILLER_3_1808 ();
 FILLCELL_X32 FILLER_3_1840 ();
 FILLCELL_X16 FILLER_3_1872 ();
 FILLCELL_X8 FILLER_3_1888 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X32 FILLER_4_1304 ();
 FILLCELL_X32 FILLER_4_1336 ();
 FILLCELL_X32 FILLER_4_1368 ();
 FILLCELL_X32 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1432 ();
 FILLCELL_X32 FILLER_4_1464 ();
 FILLCELL_X32 FILLER_4_1496 ();
 FILLCELL_X32 FILLER_4_1528 ();
 FILLCELL_X32 FILLER_4_1560 ();
 FILLCELL_X32 FILLER_4_1592 ();
 FILLCELL_X32 FILLER_4_1624 ();
 FILLCELL_X32 FILLER_4_1656 ();
 FILLCELL_X32 FILLER_4_1688 ();
 FILLCELL_X32 FILLER_4_1720 ();
 FILLCELL_X32 FILLER_4_1752 ();
 FILLCELL_X32 FILLER_4_1784 ();
 FILLCELL_X32 FILLER_4_1816 ();
 FILLCELL_X32 FILLER_4_1848 ();
 FILLCELL_X8 FILLER_4_1880 ();
 FILLCELL_X4 FILLER_4_1888 ();
 FILLCELL_X2 FILLER_4_1892 ();
 FILLCELL_X1 FILLER_4_1895 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X32 FILLER_5_1648 ();
 FILLCELL_X32 FILLER_5_1680 ();
 FILLCELL_X32 FILLER_5_1712 ();
 FILLCELL_X32 FILLER_5_1744 ();
 FILLCELL_X32 FILLER_5_1776 ();
 FILLCELL_X32 FILLER_5_1808 ();
 FILLCELL_X32 FILLER_5_1840 ();
 FILLCELL_X16 FILLER_5_1872 ();
 FILLCELL_X8 FILLER_5_1888 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X32 FILLER_6_1304 ();
 FILLCELL_X32 FILLER_6_1336 ();
 FILLCELL_X32 FILLER_6_1368 ();
 FILLCELL_X32 FILLER_6_1400 ();
 FILLCELL_X32 FILLER_6_1432 ();
 FILLCELL_X32 FILLER_6_1464 ();
 FILLCELL_X32 FILLER_6_1496 ();
 FILLCELL_X32 FILLER_6_1528 ();
 FILLCELL_X32 FILLER_6_1560 ();
 FILLCELL_X32 FILLER_6_1592 ();
 FILLCELL_X32 FILLER_6_1624 ();
 FILLCELL_X32 FILLER_6_1656 ();
 FILLCELL_X32 FILLER_6_1688 ();
 FILLCELL_X32 FILLER_6_1720 ();
 FILLCELL_X32 FILLER_6_1752 ();
 FILLCELL_X32 FILLER_6_1784 ();
 FILLCELL_X32 FILLER_6_1816 ();
 FILLCELL_X32 FILLER_6_1848 ();
 FILLCELL_X8 FILLER_6_1880 ();
 FILLCELL_X4 FILLER_6_1888 ();
 FILLCELL_X2 FILLER_6_1892 ();
 FILLCELL_X1 FILLER_6_1895 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X32 FILLER_7_1648 ();
 FILLCELL_X32 FILLER_7_1680 ();
 FILLCELL_X32 FILLER_7_1712 ();
 FILLCELL_X32 FILLER_7_1744 ();
 FILLCELL_X32 FILLER_7_1776 ();
 FILLCELL_X32 FILLER_7_1808 ();
 FILLCELL_X32 FILLER_7_1840 ();
 FILLCELL_X16 FILLER_7_1872 ();
 FILLCELL_X8 FILLER_7_1888 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X32 FILLER_8_1304 ();
 FILLCELL_X32 FILLER_8_1336 ();
 FILLCELL_X32 FILLER_8_1368 ();
 FILLCELL_X32 FILLER_8_1400 ();
 FILLCELL_X32 FILLER_8_1432 ();
 FILLCELL_X32 FILLER_8_1464 ();
 FILLCELL_X32 FILLER_8_1496 ();
 FILLCELL_X32 FILLER_8_1528 ();
 FILLCELL_X32 FILLER_8_1560 ();
 FILLCELL_X32 FILLER_8_1592 ();
 FILLCELL_X32 FILLER_8_1624 ();
 FILLCELL_X32 FILLER_8_1656 ();
 FILLCELL_X32 FILLER_8_1688 ();
 FILLCELL_X32 FILLER_8_1720 ();
 FILLCELL_X32 FILLER_8_1752 ();
 FILLCELL_X32 FILLER_8_1784 ();
 FILLCELL_X32 FILLER_8_1816 ();
 FILLCELL_X32 FILLER_8_1848 ();
 FILLCELL_X8 FILLER_8_1880 ();
 FILLCELL_X4 FILLER_8_1888 ();
 FILLCELL_X2 FILLER_8_1892 ();
 FILLCELL_X1 FILLER_8_1895 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X32 FILLER_9_1648 ();
 FILLCELL_X32 FILLER_9_1680 ();
 FILLCELL_X32 FILLER_9_1712 ();
 FILLCELL_X32 FILLER_9_1744 ();
 FILLCELL_X32 FILLER_9_1776 ();
 FILLCELL_X32 FILLER_9_1808 ();
 FILLCELL_X32 FILLER_9_1840 ();
 FILLCELL_X16 FILLER_9_1872 ();
 FILLCELL_X8 FILLER_9_1888 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X32 FILLER_10_1304 ();
 FILLCELL_X32 FILLER_10_1336 ();
 FILLCELL_X32 FILLER_10_1368 ();
 FILLCELL_X32 FILLER_10_1400 ();
 FILLCELL_X32 FILLER_10_1432 ();
 FILLCELL_X32 FILLER_10_1464 ();
 FILLCELL_X32 FILLER_10_1496 ();
 FILLCELL_X32 FILLER_10_1528 ();
 FILLCELL_X32 FILLER_10_1560 ();
 FILLCELL_X32 FILLER_10_1592 ();
 FILLCELL_X32 FILLER_10_1624 ();
 FILLCELL_X32 FILLER_10_1656 ();
 FILLCELL_X32 FILLER_10_1688 ();
 FILLCELL_X32 FILLER_10_1720 ();
 FILLCELL_X32 FILLER_10_1752 ();
 FILLCELL_X32 FILLER_10_1784 ();
 FILLCELL_X32 FILLER_10_1816 ();
 FILLCELL_X32 FILLER_10_1848 ();
 FILLCELL_X8 FILLER_10_1880 ();
 FILLCELL_X4 FILLER_10_1888 ();
 FILLCELL_X2 FILLER_10_1892 ();
 FILLCELL_X1 FILLER_10_1895 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X32 FILLER_11_1648 ();
 FILLCELL_X32 FILLER_11_1680 ();
 FILLCELL_X32 FILLER_11_1712 ();
 FILLCELL_X32 FILLER_11_1744 ();
 FILLCELL_X32 FILLER_11_1776 ();
 FILLCELL_X32 FILLER_11_1808 ();
 FILLCELL_X32 FILLER_11_1840 ();
 FILLCELL_X16 FILLER_11_1872 ();
 FILLCELL_X8 FILLER_11_1888 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X32 FILLER_12_1592 ();
 FILLCELL_X32 FILLER_12_1624 ();
 FILLCELL_X32 FILLER_12_1656 ();
 FILLCELL_X32 FILLER_12_1688 ();
 FILLCELL_X32 FILLER_12_1720 ();
 FILLCELL_X32 FILLER_12_1752 ();
 FILLCELL_X32 FILLER_12_1784 ();
 FILLCELL_X32 FILLER_12_1816 ();
 FILLCELL_X32 FILLER_12_1848 ();
 FILLCELL_X8 FILLER_12_1880 ();
 FILLCELL_X4 FILLER_12_1888 ();
 FILLCELL_X2 FILLER_12_1892 ();
 FILLCELL_X1 FILLER_12_1895 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X32 FILLER_13_1648 ();
 FILLCELL_X32 FILLER_13_1680 ();
 FILLCELL_X32 FILLER_13_1712 ();
 FILLCELL_X32 FILLER_13_1744 ();
 FILLCELL_X32 FILLER_13_1776 ();
 FILLCELL_X32 FILLER_13_1808 ();
 FILLCELL_X32 FILLER_13_1840 ();
 FILLCELL_X16 FILLER_13_1872 ();
 FILLCELL_X8 FILLER_13_1888 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X32 FILLER_14_1688 ();
 FILLCELL_X32 FILLER_14_1720 ();
 FILLCELL_X32 FILLER_14_1752 ();
 FILLCELL_X32 FILLER_14_1784 ();
 FILLCELL_X32 FILLER_14_1816 ();
 FILLCELL_X32 FILLER_14_1848 ();
 FILLCELL_X8 FILLER_14_1880 ();
 FILLCELL_X4 FILLER_14_1888 ();
 FILLCELL_X2 FILLER_14_1892 ();
 FILLCELL_X1 FILLER_14_1895 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X32 FILLER_15_1584 ();
 FILLCELL_X32 FILLER_15_1616 ();
 FILLCELL_X32 FILLER_15_1648 ();
 FILLCELL_X32 FILLER_15_1680 ();
 FILLCELL_X32 FILLER_15_1712 ();
 FILLCELL_X32 FILLER_15_1744 ();
 FILLCELL_X32 FILLER_15_1776 ();
 FILLCELL_X32 FILLER_15_1808 ();
 FILLCELL_X32 FILLER_15_1840 ();
 FILLCELL_X16 FILLER_15_1872 ();
 FILLCELL_X8 FILLER_15_1888 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X32 FILLER_16_1592 ();
 FILLCELL_X32 FILLER_16_1624 ();
 FILLCELL_X32 FILLER_16_1656 ();
 FILLCELL_X32 FILLER_16_1688 ();
 FILLCELL_X32 FILLER_16_1720 ();
 FILLCELL_X32 FILLER_16_1752 ();
 FILLCELL_X32 FILLER_16_1784 ();
 FILLCELL_X32 FILLER_16_1816 ();
 FILLCELL_X32 FILLER_16_1848 ();
 FILLCELL_X8 FILLER_16_1880 ();
 FILLCELL_X4 FILLER_16_1888 ();
 FILLCELL_X2 FILLER_16_1892 ();
 FILLCELL_X1 FILLER_16_1895 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X32 FILLER_17_1584 ();
 FILLCELL_X32 FILLER_17_1616 ();
 FILLCELL_X32 FILLER_17_1648 ();
 FILLCELL_X32 FILLER_17_1680 ();
 FILLCELL_X32 FILLER_17_1712 ();
 FILLCELL_X32 FILLER_17_1744 ();
 FILLCELL_X32 FILLER_17_1776 ();
 FILLCELL_X32 FILLER_17_1808 ();
 FILLCELL_X32 FILLER_17_1840 ();
 FILLCELL_X16 FILLER_17_1872 ();
 FILLCELL_X8 FILLER_17_1888 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X32 FILLER_18_1752 ();
 FILLCELL_X32 FILLER_18_1784 ();
 FILLCELL_X32 FILLER_18_1816 ();
 FILLCELL_X32 FILLER_18_1848 ();
 FILLCELL_X8 FILLER_18_1880 ();
 FILLCELL_X4 FILLER_18_1888 ();
 FILLCELL_X2 FILLER_18_1892 ();
 FILLCELL_X1 FILLER_18_1895 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X32 FILLER_19_1584 ();
 FILLCELL_X32 FILLER_19_1616 ();
 FILLCELL_X32 FILLER_19_1648 ();
 FILLCELL_X32 FILLER_19_1680 ();
 FILLCELL_X32 FILLER_19_1712 ();
 FILLCELL_X32 FILLER_19_1744 ();
 FILLCELL_X32 FILLER_19_1776 ();
 FILLCELL_X32 FILLER_19_1808 ();
 FILLCELL_X32 FILLER_19_1840 ();
 FILLCELL_X16 FILLER_19_1872 ();
 FILLCELL_X8 FILLER_19_1888 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X32 FILLER_20_1592 ();
 FILLCELL_X32 FILLER_20_1624 ();
 FILLCELL_X32 FILLER_20_1656 ();
 FILLCELL_X32 FILLER_20_1688 ();
 FILLCELL_X32 FILLER_20_1720 ();
 FILLCELL_X32 FILLER_20_1752 ();
 FILLCELL_X32 FILLER_20_1784 ();
 FILLCELL_X32 FILLER_20_1816 ();
 FILLCELL_X32 FILLER_20_1848 ();
 FILLCELL_X8 FILLER_20_1880 ();
 FILLCELL_X4 FILLER_20_1888 ();
 FILLCELL_X2 FILLER_20_1892 ();
 FILLCELL_X1 FILLER_20_1895 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X32 FILLER_21_1744 ();
 FILLCELL_X32 FILLER_21_1776 ();
 FILLCELL_X32 FILLER_21_1808 ();
 FILLCELL_X32 FILLER_21_1840 ();
 FILLCELL_X16 FILLER_21_1872 ();
 FILLCELL_X8 FILLER_21_1888 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X32 FILLER_22_1752 ();
 FILLCELL_X32 FILLER_22_1784 ();
 FILLCELL_X32 FILLER_22_1816 ();
 FILLCELL_X32 FILLER_22_1848 ();
 FILLCELL_X8 FILLER_22_1880 ();
 FILLCELL_X4 FILLER_22_1888 ();
 FILLCELL_X2 FILLER_22_1892 ();
 FILLCELL_X1 FILLER_22_1895 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X32 FILLER_23_1584 ();
 FILLCELL_X32 FILLER_23_1616 ();
 FILLCELL_X32 FILLER_23_1648 ();
 FILLCELL_X32 FILLER_23_1680 ();
 FILLCELL_X32 FILLER_23_1712 ();
 FILLCELL_X32 FILLER_23_1744 ();
 FILLCELL_X32 FILLER_23_1776 ();
 FILLCELL_X32 FILLER_23_1808 ();
 FILLCELL_X32 FILLER_23_1840 ();
 FILLCELL_X16 FILLER_23_1872 ();
 FILLCELL_X8 FILLER_23_1888 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X32 FILLER_24_1592 ();
 FILLCELL_X32 FILLER_24_1624 ();
 FILLCELL_X32 FILLER_24_1656 ();
 FILLCELL_X32 FILLER_24_1688 ();
 FILLCELL_X32 FILLER_24_1720 ();
 FILLCELL_X32 FILLER_24_1752 ();
 FILLCELL_X32 FILLER_24_1784 ();
 FILLCELL_X32 FILLER_24_1816 ();
 FILLCELL_X32 FILLER_24_1848 ();
 FILLCELL_X8 FILLER_24_1880 ();
 FILLCELL_X4 FILLER_24_1888 ();
 FILLCELL_X2 FILLER_24_1892 ();
 FILLCELL_X1 FILLER_24_1895 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X32 FILLER_25_1584 ();
 FILLCELL_X32 FILLER_25_1616 ();
 FILLCELL_X32 FILLER_25_1648 ();
 FILLCELL_X32 FILLER_25_1680 ();
 FILLCELL_X32 FILLER_25_1712 ();
 FILLCELL_X32 FILLER_25_1744 ();
 FILLCELL_X32 FILLER_25_1776 ();
 FILLCELL_X32 FILLER_25_1808 ();
 FILLCELL_X32 FILLER_25_1840 ();
 FILLCELL_X16 FILLER_25_1872 ();
 FILLCELL_X8 FILLER_25_1888 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X32 FILLER_26_1592 ();
 FILLCELL_X32 FILLER_26_1624 ();
 FILLCELL_X32 FILLER_26_1656 ();
 FILLCELL_X32 FILLER_26_1688 ();
 FILLCELL_X32 FILLER_26_1720 ();
 FILLCELL_X32 FILLER_26_1752 ();
 FILLCELL_X32 FILLER_26_1784 ();
 FILLCELL_X32 FILLER_26_1816 ();
 FILLCELL_X32 FILLER_26_1848 ();
 FILLCELL_X8 FILLER_26_1880 ();
 FILLCELL_X4 FILLER_26_1888 ();
 FILLCELL_X2 FILLER_26_1892 ();
 FILLCELL_X1 FILLER_26_1895 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X32 FILLER_27_1584 ();
 FILLCELL_X32 FILLER_27_1616 ();
 FILLCELL_X32 FILLER_27_1648 ();
 FILLCELL_X32 FILLER_27_1680 ();
 FILLCELL_X32 FILLER_27_1712 ();
 FILLCELL_X32 FILLER_27_1744 ();
 FILLCELL_X32 FILLER_27_1776 ();
 FILLCELL_X32 FILLER_27_1808 ();
 FILLCELL_X32 FILLER_27_1840 ();
 FILLCELL_X16 FILLER_27_1872 ();
 FILLCELL_X8 FILLER_27_1888 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X32 FILLER_28_1592 ();
 FILLCELL_X32 FILLER_28_1624 ();
 FILLCELL_X32 FILLER_28_1656 ();
 FILLCELL_X32 FILLER_28_1688 ();
 FILLCELL_X32 FILLER_28_1720 ();
 FILLCELL_X32 FILLER_28_1752 ();
 FILLCELL_X32 FILLER_28_1784 ();
 FILLCELL_X32 FILLER_28_1816 ();
 FILLCELL_X32 FILLER_28_1848 ();
 FILLCELL_X8 FILLER_28_1880 ();
 FILLCELL_X4 FILLER_28_1888 ();
 FILLCELL_X2 FILLER_28_1892 ();
 FILLCELL_X1 FILLER_28_1895 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X32 FILLER_29_1584 ();
 FILLCELL_X32 FILLER_29_1616 ();
 FILLCELL_X32 FILLER_29_1648 ();
 FILLCELL_X32 FILLER_29_1680 ();
 FILLCELL_X32 FILLER_29_1712 ();
 FILLCELL_X32 FILLER_29_1744 ();
 FILLCELL_X32 FILLER_29_1776 ();
 FILLCELL_X32 FILLER_29_1808 ();
 FILLCELL_X32 FILLER_29_1840 ();
 FILLCELL_X16 FILLER_29_1872 ();
 FILLCELL_X8 FILLER_29_1888 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X32 FILLER_30_1592 ();
 FILLCELL_X32 FILLER_30_1624 ();
 FILLCELL_X32 FILLER_30_1656 ();
 FILLCELL_X32 FILLER_30_1688 ();
 FILLCELL_X32 FILLER_30_1720 ();
 FILLCELL_X32 FILLER_30_1752 ();
 FILLCELL_X32 FILLER_30_1784 ();
 FILLCELL_X32 FILLER_30_1816 ();
 FILLCELL_X32 FILLER_30_1848 ();
 FILLCELL_X8 FILLER_30_1880 ();
 FILLCELL_X4 FILLER_30_1888 ();
 FILLCELL_X2 FILLER_30_1892 ();
 FILLCELL_X1 FILLER_30_1895 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X32 FILLER_31_1584 ();
 FILLCELL_X32 FILLER_31_1616 ();
 FILLCELL_X32 FILLER_31_1648 ();
 FILLCELL_X32 FILLER_31_1680 ();
 FILLCELL_X32 FILLER_31_1712 ();
 FILLCELL_X32 FILLER_31_1744 ();
 FILLCELL_X32 FILLER_31_1776 ();
 FILLCELL_X32 FILLER_31_1808 ();
 FILLCELL_X32 FILLER_31_1840 ();
 FILLCELL_X16 FILLER_31_1872 ();
 FILLCELL_X8 FILLER_31_1888 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X32 FILLER_32_1592 ();
 FILLCELL_X32 FILLER_32_1624 ();
 FILLCELL_X32 FILLER_32_1656 ();
 FILLCELL_X32 FILLER_32_1688 ();
 FILLCELL_X32 FILLER_32_1720 ();
 FILLCELL_X32 FILLER_32_1752 ();
 FILLCELL_X32 FILLER_32_1784 ();
 FILLCELL_X32 FILLER_32_1816 ();
 FILLCELL_X32 FILLER_32_1848 ();
 FILLCELL_X8 FILLER_32_1880 ();
 FILLCELL_X4 FILLER_32_1888 ();
 FILLCELL_X2 FILLER_32_1892 ();
 FILLCELL_X1 FILLER_32_1895 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X32 FILLER_33_1584 ();
 FILLCELL_X32 FILLER_33_1616 ();
 FILLCELL_X32 FILLER_33_1648 ();
 FILLCELL_X32 FILLER_33_1680 ();
 FILLCELL_X32 FILLER_33_1712 ();
 FILLCELL_X32 FILLER_33_1744 ();
 FILLCELL_X32 FILLER_33_1776 ();
 FILLCELL_X32 FILLER_33_1808 ();
 FILLCELL_X32 FILLER_33_1840 ();
 FILLCELL_X16 FILLER_33_1872 ();
 FILLCELL_X8 FILLER_33_1888 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X32 FILLER_34_1592 ();
 FILLCELL_X32 FILLER_34_1624 ();
 FILLCELL_X32 FILLER_34_1656 ();
 FILLCELL_X32 FILLER_34_1688 ();
 FILLCELL_X32 FILLER_34_1720 ();
 FILLCELL_X32 FILLER_34_1752 ();
 FILLCELL_X32 FILLER_34_1784 ();
 FILLCELL_X32 FILLER_34_1816 ();
 FILLCELL_X32 FILLER_34_1848 ();
 FILLCELL_X8 FILLER_34_1880 ();
 FILLCELL_X4 FILLER_34_1888 ();
 FILLCELL_X2 FILLER_34_1892 ();
 FILLCELL_X1 FILLER_34_1895 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X32 FILLER_35_1584 ();
 FILLCELL_X32 FILLER_35_1616 ();
 FILLCELL_X32 FILLER_35_1648 ();
 FILLCELL_X32 FILLER_35_1680 ();
 FILLCELL_X32 FILLER_35_1712 ();
 FILLCELL_X32 FILLER_35_1744 ();
 FILLCELL_X32 FILLER_35_1776 ();
 FILLCELL_X32 FILLER_35_1808 ();
 FILLCELL_X32 FILLER_35_1840 ();
 FILLCELL_X16 FILLER_35_1872 ();
 FILLCELL_X8 FILLER_35_1888 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X32 FILLER_36_1592 ();
 FILLCELL_X32 FILLER_36_1624 ();
 FILLCELL_X32 FILLER_36_1656 ();
 FILLCELL_X32 FILLER_36_1688 ();
 FILLCELL_X32 FILLER_36_1720 ();
 FILLCELL_X32 FILLER_36_1752 ();
 FILLCELL_X32 FILLER_36_1784 ();
 FILLCELL_X32 FILLER_36_1816 ();
 FILLCELL_X32 FILLER_36_1848 ();
 FILLCELL_X8 FILLER_36_1880 ();
 FILLCELL_X4 FILLER_36_1888 ();
 FILLCELL_X2 FILLER_36_1892 ();
 FILLCELL_X1 FILLER_36_1895 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X32 FILLER_37_1584 ();
 FILLCELL_X32 FILLER_37_1616 ();
 FILLCELL_X32 FILLER_37_1648 ();
 FILLCELL_X32 FILLER_37_1680 ();
 FILLCELL_X32 FILLER_37_1712 ();
 FILLCELL_X32 FILLER_37_1744 ();
 FILLCELL_X32 FILLER_37_1776 ();
 FILLCELL_X32 FILLER_37_1808 ();
 FILLCELL_X32 FILLER_37_1840 ();
 FILLCELL_X16 FILLER_37_1872 ();
 FILLCELL_X8 FILLER_37_1888 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X32 FILLER_38_1592 ();
 FILLCELL_X32 FILLER_38_1624 ();
 FILLCELL_X32 FILLER_38_1656 ();
 FILLCELL_X32 FILLER_38_1688 ();
 FILLCELL_X32 FILLER_38_1720 ();
 FILLCELL_X32 FILLER_38_1752 ();
 FILLCELL_X32 FILLER_38_1784 ();
 FILLCELL_X32 FILLER_38_1816 ();
 FILLCELL_X32 FILLER_38_1848 ();
 FILLCELL_X8 FILLER_38_1880 ();
 FILLCELL_X4 FILLER_38_1888 ();
 FILLCELL_X2 FILLER_38_1892 ();
 FILLCELL_X1 FILLER_38_1895 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X32 FILLER_39_1584 ();
 FILLCELL_X32 FILLER_39_1616 ();
 FILLCELL_X32 FILLER_39_1648 ();
 FILLCELL_X32 FILLER_39_1680 ();
 FILLCELL_X32 FILLER_39_1712 ();
 FILLCELL_X32 FILLER_39_1744 ();
 FILLCELL_X32 FILLER_39_1776 ();
 FILLCELL_X32 FILLER_39_1808 ();
 FILLCELL_X32 FILLER_39_1840 ();
 FILLCELL_X16 FILLER_39_1872 ();
 FILLCELL_X8 FILLER_39_1888 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X32 FILLER_40_1592 ();
 FILLCELL_X32 FILLER_40_1624 ();
 FILLCELL_X32 FILLER_40_1656 ();
 FILLCELL_X32 FILLER_40_1688 ();
 FILLCELL_X32 FILLER_40_1720 ();
 FILLCELL_X32 FILLER_40_1752 ();
 FILLCELL_X32 FILLER_40_1784 ();
 FILLCELL_X32 FILLER_40_1816 ();
 FILLCELL_X32 FILLER_40_1848 ();
 FILLCELL_X8 FILLER_40_1880 ();
 FILLCELL_X4 FILLER_40_1888 ();
 FILLCELL_X2 FILLER_40_1892 ();
 FILLCELL_X1 FILLER_40_1895 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X32 FILLER_41_1584 ();
 FILLCELL_X32 FILLER_41_1616 ();
 FILLCELL_X32 FILLER_41_1648 ();
 FILLCELL_X32 FILLER_41_1680 ();
 FILLCELL_X32 FILLER_41_1712 ();
 FILLCELL_X32 FILLER_41_1744 ();
 FILLCELL_X32 FILLER_41_1776 ();
 FILLCELL_X32 FILLER_41_1808 ();
 FILLCELL_X32 FILLER_41_1840 ();
 FILLCELL_X16 FILLER_41_1872 ();
 FILLCELL_X8 FILLER_41_1888 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X32 FILLER_42_1592 ();
 FILLCELL_X32 FILLER_42_1624 ();
 FILLCELL_X32 FILLER_42_1656 ();
 FILLCELL_X32 FILLER_42_1688 ();
 FILLCELL_X32 FILLER_42_1720 ();
 FILLCELL_X32 FILLER_42_1752 ();
 FILLCELL_X32 FILLER_42_1784 ();
 FILLCELL_X32 FILLER_42_1816 ();
 FILLCELL_X32 FILLER_42_1848 ();
 FILLCELL_X8 FILLER_42_1880 ();
 FILLCELL_X4 FILLER_42_1888 ();
 FILLCELL_X2 FILLER_42_1892 ();
 FILLCELL_X1 FILLER_42_1895 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X32 FILLER_43_1584 ();
 FILLCELL_X32 FILLER_43_1616 ();
 FILLCELL_X32 FILLER_43_1648 ();
 FILLCELL_X32 FILLER_43_1680 ();
 FILLCELL_X32 FILLER_43_1712 ();
 FILLCELL_X32 FILLER_43_1744 ();
 FILLCELL_X32 FILLER_43_1776 ();
 FILLCELL_X32 FILLER_43_1808 ();
 FILLCELL_X32 FILLER_43_1840 ();
 FILLCELL_X16 FILLER_43_1872 ();
 FILLCELL_X8 FILLER_43_1888 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X32 FILLER_44_1592 ();
 FILLCELL_X32 FILLER_44_1624 ();
 FILLCELL_X32 FILLER_44_1656 ();
 FILLCELL_X32 FILLER_44_1688 ();
 FILLCELL_X32 FILLER_44_1720 ();
 FILLCELL_X32 FILLER_44_1752 ();
 FILLCELL_X32 FILLER_44_1784 ();
 FILLCELL_X32 FILLER_44_1816 ();
 FILLCELL_X32 FILLER_44_1848 ();
 FILLCELL_X8 FILLER_44_1880 ();
 FILLCELL_X4 FILLER_44_1888 ();
 FILLCELL_X2 FILLER_44_1892 ();
 FILLCELL_X1 FILLER_44_1895 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X32 FILLER_45_1584 ();
 FILLCELL_X32 FILLER_45_1616 ();
 FILLCELL_X32 FILLER_45_1648 ();
 FILLCELL_X32 FILLER_45_1680 ();
 FILLCELL_X32 FILLER_45_1712 ();
 FILLCELL_X32 FILLER_45_1744 ();
 FILLCELL_X32 FILLER_45_1776 ();
 FILLCELL_X32 FILLER_45_1808 ();
 FILLCELL_X32 FILLER_45_1840 ();
 FILLCELL_X16 FILLER_45_1872 ();
 FILLCELL_X8 FILLER_45_1888 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X32 FILLER_46_1592 ();
 FILLCELL_X32 FILLER_46_1624 ();
 FILLCELL_X32 FILLER_46_1656 ();
 FILLCELL_X32 FILLER_46_1688 ();
 FILLCELL_X32 FILLER_46_1720 ();
 FILLCELL_X32 FILLER_46_1752 ();
 FILLCELL_X32 FILLER_46_1784 ();
 FILLCELL_X32 FILLER_46_1816 ();
 FILLCELL_X32 FILLER_46_1848 ();
 FILLCELL_X8 FILLER_46_1880 ();
 FILLCELL_X4 FILLER_46_1888 ();
 FILLCELL_X2 FILLER_46_1892 ();
 FILLCELL_X1 FILLER_46_1895 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X32 FILLER_47_1584 ();
 FILLCELL_X32 FILLER_47_1616 ();
 FILLCELL_X32 FILLER_47_1648 ();
 FILLCELL_X32 FILLER_47_1680 ();
 FILLCELL_X32 FILLER_47_1712 ();
 FILLCELL_X32 FILLER_47_1744 ();
 FILLCELL_X32 FILLER_47_1776 ();
 FILLCELL_X32 FILLER_47_1808 ();
 FILLCELL_X32 FILLER_47_1840 ();
 FILLCELL_X16 FILLER_47_1872 ();
 FILLCELL_X8 FILLER_47_1888 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X32 FILLER_48_1592 ();
 FILLCELL_X32 FILLER_48_1624 ();
 FILLCELL_X32 FILLER_48_1656 ();
 FILLCELL_X32 FILLER_48_1688 ();
 FILLCELL_X32 FILLER_48_1720 ();
 FILLCELL_X32 FILLER_48_1752 ();
 FILLCELL_X32 FILLER_48_1784 ();
 FILLCELL_X32 FILLER_48_1816 ();
 FILLCELL_X32 FILLER_48_1848 ();
 FILLCELL_X8 FILLER_48_1880 ();
 FILLCELL_X4 FILLER_48_1888 ();
 FILLCELL_X2 FILLER_48_1892 ();
 FILLCELL_X1 FILLER_48_1895 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X32 FILLER_49_1584 ();
 FILLCELL_X32 FILLER_49_1616 ();
 FILLCELL_X32 FILLER_49_1648 ();
 FILLCELL_X32 FILLER_49_1680 ();
 FILLCELL_X32 FILLER_49_1712 ();
 FILLCELL_X32 FILLER_49_1744 ();
 FILLCELL_X32 FILLER_49_1776 ();
 FILLCELL_X32 FILLER_49_1808 ();
 FILLCELL_X32 FILLER_49_1840 ();
 FILLCELL_X16 FILLER_49_1872 ();
 FILLCELL_X8 FILLER_49_1888 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X32 FILLER_50_1592 ();
 FILLCELL_X32 FILLER_50_1624 ();
 FILLCELL_X32 FILLER_50_1656 ();
 FILLCELL_X32 FILLER_50_1688 ();
 FILLCELL_X32 FILLER_50_1720 ();
 FILLCELL_X32 FILLER_50_1752 ();
 FILLCELL_X32 FILLER_50_1784 ();
 FILLCELL_X32 FILLER_50_1816 ();
 FILLCELL_X32 FILLER_50_1848 ();
 FILLCELL_X8 FILLER_50_1880 ();
 FILLCELL_X4 FILLER_50_1888 ();
 FILLCELL_X2 FILLER_50_1892 ();
 FILLCELL_X1 FILLER_50_1895 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X32 FILLER_51_1584 ();
 FILLCELL_X32 FILLER_51_1616 ();
 FILLCELL_X32 FILLER_51_1648 ();
 FILLCELL_X32 FILLER_51_1680 ();
 FILLCELL_X32 FILLER_51_1712 ();
 FILLCELL_X32 FILLER_51_1744 ();
 FILLCELL_X32 FILLER_51_1776 ();
 FILLCELL_X32 FILLER_51_1808 ();
 FILLCELL_X32 FILLER_51_1840 ();
 FILLCELL_X16 FILLER_51_1872 ();
 FILLCELL_X8 FILLER_51_1888 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X32 FILLER_52_1592 ();
 FILLCELL_X32 FILLER_52_1624 ();
 FILLCELL_X32 FILLER_52_1656 ();
 FILLCELL_X32 FILLER_52_1688 ();
 FILLCELL_X32 FILLER_52_1720 ();
 FILLCELL_X32 FILLER_52_1752 ();
 FILLCELL_X32 FILLER_52_1784 ();
 FILLCELL_X32 FILLER_52_1816 ();
 FILLCELL_X32 FILLER_52_1848 ();
 FILLCELL_X8 FILLER_52_1880 ();
 FILLCELL_X4 FILLER_52_1888 ();
 FILLCELL_X2 FILLER_52_1892 ();
 FILLCELL_X1 FILLER_52_1895 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X32 FILLER_53_1584 ();
 FILLCELL_X32 FILLER_53_1616 ();
 FILLCELL_X32 FILLER_53_1648 ();
 FILLCELL_X32 FILLER_53_1680 ();
 FILLCELL_X32 FILLER_53_1712 ();
 FILLCELL_X32 FILLER_53_1744 ();
 FILLCELL_X32 FILLER_53_1776 ();
 FILLCELL_X32 FILLER_53_1808 ();
 FILLCELL_X32 FILLER_53_1840 ();
 FILLCELL_X16 FILLER_53_1872 ();
 FILLCELL_X8 FILLER_53_1888 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X32 FILLER_54_1592 ();
 FILLCELL_X32 FILLER_54_1624 ();
 FILLCELL_X32 FILLER_54_1656 ();
 FILLCELL_X32 FILLER_54_1688 ();
 FILLCELL_X32 FILLER_54_1720 ();
 FILLCELL_X32 FILLER_54_1752 ();
 FILLCELL_X32 FILLER_54_1784 ();
 FILLCELL_X32 FILLER_54_1816 ();
 FILLCELL_X32 FILLER_54_1848 ();
 FILLCELL_X8 FILLER_54_1880 ();
 FILLCELL_X4 FILLER_54_1888 ();
 FILLCELL_X2 FILLER_54_1892 ();
 FILLCELL_X1 FILLER_54_1895 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X32 FILLER_55_1584 ();
 FILLCELL_X32 FILLER_55_1616 ();
 FILLCELL_X32 FILLER_55_1648 ();
 FILLCELL_X32 FILLER_55_1680 ();
 FILLCELL_X32 FILLER_55_1712 ();
 FILLCELL_X32 FILLER_55_1744 ();
 FILLCELL_X32 FILLER_55_1776 ();
 FILLCELL_X32 FILLER_55_1808 ();
 FILLCELL_X32 FILLER_55_1840 ();
 FILLCELL_X16 FILLER_55_1872 ();
 FILLCELL_X8 FILLER_55_1888 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X32 FILLER_56_1592 ();
 FILLCELL_X32 FILLER_56_1624 ();
 FILLCELL_X32 FILLER_56_1656 ();
 FILLCELL_X32 FILLER_56_1688 ();
 FILLCELL_X32 FILLER_56_1720 ();
 FILLCELL_X32 FILLER_56_1752 ();
 FILLCELL_X32 FILLER_56_1784 ();
 FILLCELL_X32 FILLER_56_1816 ();
 FILLCELL_X32 FILLER_56_1848 ();
 FILLCELL_X8 FILLER_56_1880 ();
 FILLCELL_X4 FILLER_56_1888 ();
 FILLCELL_X2 FILLER_56_1892 ();
 FILLCELL_X1 FILLER_56_1895 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X32 FILLER_57_1584 ();
 FILLCELL_X32 FILLER_57_1616 ();
 FILLCELL_X32 FILLER_57_1648 ();
 FILLCELL_X32 FILLER_57_1680 ();
 FILLCELL_X32 FILLER_57_1712 ();
 FILLCELL_X32 FILLER_57_1744 ();
 FILLCELL_X32 FILLER_57_1776 ();
 FILLCELL_X32 FILLER_57_1808 ();
 FILLCELL_X32 FILLER_57_1840 ();
 FILLCELL_X16 FILLER_57_1872 ();
 FILLCELL_X8 FILLER_57_1888 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X32 FILLER_58_1592 ();
 FILLCELL_X32 FILLER_58_1624 ();
 FILLCELL_X32 FILLER_58_1656 ();
 FILLCELL_X32 FILLER_58_1688 ();
 FILLCELL_X32 FILLER_58_1720 ();
 FILLCELL_X32 FILLER_58_1752 ();
 FILLCELL_X32 FILLER_58_1784 ();
 FILLCELL_X32 FILLER_58_1816 ();
 FILLCELL_X32 FILLER_58_1848 ();
 FILLCELL_X8 FILLER_58_1880 ();
 FILLCELL_X4 FILLER_58_1888 ();
 FILLCELL_X2 FILLER_58_1892 ();
 FILLCELL_X1 FILLER_58_1895 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X32 FILLER_59_1584 ();
 FILLCELL_X32 FILLER_59_1616 ();
 FILLCELL_X32 FILLER_59_1648 ();
 FILLCELL_X32 FILLER_59_1680 ();
 FILLCELL_X32 FILLER_59_1712 ();
 FILLCELL_X32 FILLER_59_1744 ();
 FILLCELL_X32 FILLER_59_1776 ();
 FILLCELL_X32 FILLER_59_1808 ();
 FILLCELL_X32 FILLER_59_1840 ();
 FILLCELL_X16 FILLER_59_1872 ();
 FILLCELL_X8 FILLER_59_1888 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X32 FILLER_60_1592 ();
 FILLCELL_X32 FILLER_60_1624 ();
 FILLCELL_X32 FILLER_60_1656 ();
 FILLCELL_X32 FILLER_60_1688 ();
 FILLCELL_X32 FILLER_60_1720 ();
 FILLCELL_X32 FILLER_60_1752 ();
 FILLCELL_X32 FILLER_60_1784 ();
 FILLCELL_X32 FILLER_60_1816 ();
 FILLCELL_X32 FILLER_60_1848 ();
 FILLCELL_X8 FILLER_60_1880 ();
 FILLCELL_X4 FILLER_60_1888 ();
 FILLCELL_X2 FILLER_60_1892 ();
 FILLCELL_X1 FILLER_60_1895 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X32 FILLER_61_1584 ();
 FILLCELL_X32 FILLER_61_1616 ();
 FILLCELL_X32 FILLER_61_1648 ();
 FILLCELL_X32 FILLER_61_1680 ();
 FILLCELL_X32 FILLER_61_1712 ();
 FILLCELL_X32 FILLER_61_1744 ();
 FILLCELL_X32 FILLER_61_1776 ();
 FILLCELL_X32 FILLER_61_1808 ();
 FILLCELL_X32 FILLER_61_1840 ();
 FILLCELL_X16 FILLER_61_1872 ();
 FILLCELL_X8 FILLER_61_1888 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X32 FILLER_62_1592 ();
 FILLCELL_X32 FILLER_62_1624 ();
 FILLCELL_X32 FILLER_62_1656 ();
 FILLCELL_X32 FILLER_62_1688 ();
 FILLCELL_X32 FILLER_62_1720 ();
 FILLCELL_X32 FILLER_62_1752 ();
 FILLCELL_X32 FILLER_62_1784 ();
 FILLCELL_X32 FILLER_62_1816 ();
 FILLCELL_X32 FILLER_62_1848 ();
 FILLCELL_X8 FILLER_62_1880 ();
 FILLCELL_X4 FILLER_62_1888 ();
 FILLCELL_X2 FILLER_62_1892 ();
 FILLCELL_X1 FILLER_62_1895 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X32 FILLER_63_1584 ();
 FILLCELL_X32 FILLER_63_1616 ();
 FILLCELL_X32 FILLER_63_1648 ();
 FILLCELL_X32 FILLER_63_1680 ();
 FILLCELL_X32 FILLER_63_1712 ();
 FILLCELL_X32 FILLER_63_1744 ();
 FILLCELL_X32 FILLER_63_1776 ();
 FILLCELL_X32 FILLER_63_1808 ();
 FILLCELL_X32 FILLER_63_1840 ();
 FILLCELL_X16 FILLER_63_1872 ();
 FILLCELL_X8 FILLER_63_1888 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X32 FILLER_64_1592 ();
 FILLCELL_X32 FILLER_64_1624 ();
 FILLCELL_X32 FILLER_64_1656 ();
 FILLCELL_X32 FILLER_64_1688 ();
 FILLCELL_X32 FILLER_64_1720 ();
 FILLCELL_X32 FILLER_64_1752 ();
 FILLCELL_X32 FILLER_64_1784 ();
 FILLCELL_X32 FILLER_64_1816 ();
 FILLCELL_X32 FILLER_64_1848 ();
 FILLCELL_X8 FILLER_64_1880 ();
 FILLCELL_X4 FILLER_64_1888 ();
 FILLCELL_X2 FILLER_64_1892 ();
 FILLCELL_X1 FILLER_64_1895 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X32 FILLER_65_1584 ();
 FILLCELL_X32 FILLER_65_1616 ();
 FILLCELL_X32 FILLER_65_1648 ();
 FILLCELL_X32 FILLER_65_1680 ();
 FILLCELL_X32 FILLER_65_1712 ();
 FILLCELL_X32 FILLER_65_1744 ();
 FILLCELL_X32 FILLER_65_1776 ();
 FILLCELL_X32 FILLER_65_1808 ();
 FILLCELL_X32 FILLER_65_1840 ();
 FILLCELL_X16 FILLER_65_1872 ();
 FILLCELL_X8 FILLER_65_1888 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X32 FILLER_66_1592 ();
 FILLCELL_X32 FILLER_66_1624 ();
 FILLCELL_X32 FILLER_66_1656 ();
 FILLCELL_X32 FILLER_66_1688 ();
 FILLCELL_X32 FILLER_66_1720 ();
 FILLCELL_X32 FILLER_66_1752 ();
 FILLCELL_X32 FILLER_66_1784 ();
 FILLCELL_X32 FILLER_66_1816 ();
 FILLCELL_X32 FILLER_66_1848 ();
 FILLCELL_X8 FILLER_66_1880 ();
 FILLCELL_X4 FILLER_66_1888 ();
 FILLCELL_X2 FILLER_66_1892 ();
 FILLCELL_X1 FILLER_66_1895 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X32 FILLER_67_801 ();
 FILLCELL_X32 FILLER_67_833 ();
 FILLCELL_X32 FILLER_67_865 ();
 FILLCELL_X32 FILLER_67_897 ();
 FILLCELL_X32 FILLER_67_929 ();
 FILLCELL_X32 FILLER_67_961 ();
 FILLCELL_X32 FILLER_67_993 ();
 FILLCELL_X32 FILLER_67_1025 ();
 FILLCELL_X32 FILLER_67_1057 ();
 FILLCELL_X32 FILLER_67_1089 ();
 FILLCELL_X32 FILLER_67_1121 ();
 FILLCELL_X32 FILLER_67_1153 ();
 FILLCELL_X32 FILLER_67_1185 ();
 FILLCELL_X32 FILLER_67_1217 ();
 FILLCELL_X8 FILLER_67_1249 ();
 FILLCELL_X4 FILLER_67_1257 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X32 FILLER_67_1584 ();
 FILLCELL_X32 FILLER_67_1616 ();
 FILLCELL_X32 FILLER_67_1648 ();
 FILLCELL_X32 FILLER_67_1680 ();
 FILLCELL_X32 FILLER_67_1712 ();
 FILLCELL_X32 FILLER_67_1744 ();
 FILLCELL_X32 FILLER_67_1776 ();
 FILLCELL_X32 FILLER_67_1808 ();
 FILLCELL_X32 FILLER_67_1840 ();
 FILLCELL_X16 FILLER_67_1872 ();
 FILLCELL_X8 FILLER_67_1888 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X32 FILLER_68_952 ();
 FILLCELL_X32 FILLER_68_984 ();
 FILLCELL_X32 FILLER_68_1016 ();
 FILLCELL_X32 FILLER_68_1048 ();
 FILLCELL_X32 FILLER_68_1080 ();
 FILLCELL_X32 FILLER_68_1112 ();
 FILLCELL_X32 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_68_1176 ();
 FILLCELL_X32 FILLER_68_1208 ();
 FILLCELL_X32 FILLER_68_1240 ();
 FILLCELL_X32 FILLER_68_1272 ();
 FILLCELL_X32 FILLER_68_1304 ();
 FILLCELL_X32 FILLER_68_1336 ();
 FILLCELL_X32 FILLER_68_1368 ();
 FILLCELL_X32 FILLER_68_1400 ();
 FILLCELL_X32 FILLER_68_1432 ();
 FILLCELL_X32 FILLER_68_1464 ();
 FILLCELL_X32 FILLER_68_1496 ();
 FILLCELL_X32 FILLER_68_1528 ();
 FILLCELL_X32 FILLER_68_1560 ();
 FILLCELL_X32 FILLER_68_1592 ();
 FILLCELL_X32 FILLER_68_1624 ();
 FILLCELL_X32 FILLER_68_1656 ();
 FILLCELL_X32 FILLER_68_1688 ();
 FILLCELL_X32 FILLER_68_1720 ();
 FILLCELL_X32 FILLER_68_1752 ();
 FILLCELL_X32 FILLER_68_1784 ();
 FILLCELL_X32 FILLER_68_1816 ();
 FILLCELL_X32 FILLER_68_1848 ();
 FILLCELL_X8 FILLER_68_1880 ();
 FILLCELL_X4 FILLER_68_1888 ();
 FILLCELL_X2 FILLER_68_1892 ();
 FILLCELL_X1 FILLER_68_1895 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X32 FILLER_69_833 ();
 FILLCELL_X32 FILLER_69_865 ();
 FILLCELL_X32 FILLER_69_897 ();
 FILLCELL_X32 FILLER_69_929 ();
 FILLCELL_X32 FILLER_69_961 ();
 FILLCELL_X32 FILLER_69_993 ();
 FILLCELL_X32 FILLER_69_1025 ();
 FILLCELL_X32 FILLER_69_1057 ();
 FILLCELL_X32 FILLER_69_1089 ();
 FILLCELL_X32 FILLER_69_1121 ();
 FILLCELL_X32 FILLER_69_1153 ();
 FILLCELL_X32 FILLER_69_1185 ();
 FILLCELL_X32 FILLER_69_1217 ();
 FILLCELL_X8 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1257 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X32 FILLER_69_1584 ();
 FILLCELL_X32 FILLER_69_1616 ();
 FILLCELL_X32 FILLER_69_1648 ();
 FILLCELL_X32 FILLER_69_1680 ();
 FILLCELL_X32 FILLER_69_1712 ();
 FILLCELL_X32 FILLER_69_1744 ();
 FILLCELL_X32 FILLER_69_1776 ();
 FILLCELL_X32 FILLER_69_1808 ();
 FILLCELL_X32 FILLER_69_1840 ();
 FILLCELL_X16 FILLER_69_1872 ();
 FILLCELL_X8 FILLER_69_1888 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X32 FILLER_70_1592 ();
 FILLCELL_X32 FILLER_70_1624 ();
 FILLCELL_X32 FILLER_70_1656 ();
 FILLCELL_X32 FILLER_70_1688 ();
 FILLCELL_X32 FILLER_70_1720 ();
 FILLCELL_X32 FILLER_70_1752 ();
 FILLCELL_X32 FILLER_70_1784 ();
 FILLCELL_X32 FILLER_70_1816 ();
 FILLCELL_X32 FILLER_70_1848 ();
 FILLCELL_X8 FILLER_70_1880 ();
 FILLCELL_X4 FILLER_70_1888 ();
 FILLCELL_X2 FILLER_70_1892 ();
 FILLCELL_X1 FILLER_70_1895 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1584 ();
 FILLCELL_X32 FILLER_71_1616 ();
 FILLCELL_X32 FILLER_71_1648 ();
 FILLCELL_X32 FILLER_71_1680 ();
 FILLCELL_X32 FILLER_71_1712 ();
 FILLCELL_X32 FILLER_71_1744 ();
 FILLCELL_X32 FILLER_71_1776 ();
 FILLCELL_X32 FILLER_71_1808 ();
 FILLCELL_X32 FILLER_71_1840 ();
 FILLCELL_X16 FILLER_71_1872 ();
 FILLCELL_X8 FILLER_71_1888 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X32 FILLER_72_1592 ();
 FILLCELL_X32 FILLER_72_1624 ();
 FILLCELL_X32 FILLER_72_1656 ();
 FILLCELL_X32 FILLER_72_1688 ();
 FILLCELL_X32 FILLER_72_1720 ();
 FILLCELL_X32 FILLER_72_1752 ();
 FILLCELL_X32 FILLER_72_1784 ();
 FILLCELL_X32 FILLER_72_1816 ();
 FILLCELL_X32 FILLER_72_1848 ();
 FILLCELL_X8 FILLER_72_1880 ();
 FILLCELL_X4 FILLER_72_1888 ();
 FILLCELL_X2 FILLER_72_1892 ();
 FILLCELL_X1 FILLER_72_1895 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X32 FILLER_73_1584 ();
 FILLCELL_X32 FILLER_73_1616 ();
 FILLCELL_X32 FILLER_73_1648 ();
 FILLCELL_X32 FILLER_73_1680 ();
 FILLCELL_X32 FILLER_73_1712 ();
 FILLCELL_X32 FILLER_73_1744 ();
 FILLCELL_X32 FILLER_73_1776 ();
 FILLCELL_X32 FILLER_73_1808 ();
 FILLCELL_X32 FILLER_73_1840 ();
 FILLCELL_X16 FILLER_73_1872 ();
 FILLCELL_X8 FILLER_73_1888 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X32 FILLER_74_1592 ();
 FILLCELL_X32 FILLER_74_1624 ();
 FILLCELL_X32 FILLER_74_1656 ();
 FILLCELL_X32 FILLER_74_1688 ();
 FILLCELL_X32 FILLER_74_1720 ();
 FILLCELL_X32 FILLER_74_1752 ();
 FILLCELL_X32 FILLER_74_1784 ();
 FILLCELL_X32 FILLER_74_1816 ();
 FILLCELL_X32 FILLER_74_1848 ();
 FILLCELL_X8 FILLER_74_1880 ();
 FILLCELL_X4 FILLER_74_1888 ();
 FILLCELL_X2 FILLER_74_1892 ();
 FILLCELL_X1 FILLER_74_1895 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X32 FILLER_75_865 ();
 FILLCELL_X32 FILLER_75_897 ();
 FILLCELL_X32 FILLER_75_929 ();
 FILLCELL_X32 FILLER_75_961 ();
 FILLCELL_X32 FILLER_75_993 ();
 FILLCELL_X32 FILLER_75_1025 ();
 FILLCELL_X32 FILLER_75_1057 ();
 FILLCELL_X32 FILLER_75_1089 ();
 FILLCELL_X32 FILLER_75_1121 ();
 FILLCELL_X32 FILLER_75_1153 ();
 FILLCELL_X32 FILLER_75_1185 ();
 FILLCELL_X32 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1249 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X32 FILLER_75_1584 ();
 FILLCELL_X32 FILLER_75_1616 ();
 FILLCELL_X32 FILLER_75_1648 ();
 FILLCELL_X32 FILLER_75_1680 ();
 FILLCELL_X32 FILLER_75_1712 ();
 FILLCELL_X32 FILLER_75_1744 ();
 FILLCELL_X32 FILLER_75_1776 ();
 FILLCELL_X32 FILLER_75_1808 ();
 FILLCELL_X32 FILLER_75_1840 ();
 FILLCELL_X16 FILLER_75_1872 ();
 FILLCELL_X8 FILLER_75_1888 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X32 FILLER_76_952 ();
 FILLCELL_X32 FILLER_76_984 ();
 FILLCELL_X32 FILLER_76_1016 ();
 FILLCELL_X32 FILLER_76_1048 ();
 FILLCELL_X32 FILLER_76_1080 ();
 FILLCELL_X32 FILLER_76_1112 ();
 FILLCELL_X32 FILLER_76_1144 ();
 FILLCELL_X32 FILLER_76_1176 ();
 FILLCELL_X32 FILLER_76_1208 ();
 FILLCELL_X32 FILLER_76_1240 ();
 FILLCELL_X32 FILLER_76_1272 ();
 FILLCELL_X32 FILLER_76_1304 ();
 FILLCELL_X32 FILLER_76_1336 ();
 FILLCELL_X32 FILLER_76_1368 ();
 FILLCELL_X32 FILLER_76_1400 ();
 FILLCELL_X32 FILLER_76_1432 ();
 FILLCELL_X32 FILLER_76_1464 ();
 FILLCELL_X32 FILLER_76_1496 ();
 FILLCELL_X32 FILLER_76_1528 ();
 FILLCELL_X32 FILLER_76_1560 ();
 FILLCELL_X32 FILLER_76_1592 ();
 FILLCELL_X32 FILLER_76_1624 ();
 FILLCELL_X32 FILLER_76_1656 ();
 FILLCELL_X32 FILLER_76_1688 ();
 FILLCELL_X32 FILLER_76_1720 ();
 FILLCELL_X32 FILLER_76_1752 ();
 FILLCELL_X32 FILLER_76_1784 ();
 FILLCELL_X32 FILLER_76_1816 ();
 FILLCELL_X32 FILLER_76_1848 ();
 FILLCELL_X8 FILLER_76_1880 ();
 FILLCELL_X4 FILLER_76_1888 ();
 FILLCELL_X2 FILLER_76_1892 ();
 FILLCELL_X1 FILLER_76_1895 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_961 ();
 FILLCELL_X32 FILLER_77_993 ();
 FILLCELL_X32 FILLER_77_1025 ();
 FILLCELL_X32 FILLER_77_1057 ();
 FILLCELL_X32 FILLER_77_1089 ();
 FILLCELL_X32 FILLER_77_1121 ();
 FILLCELL_X32 FILLER_77_1153 ();
 FILLCELL_X32 FILLER_77_1185 ();
 FILLCELL_X32 FILLER_77_1217 ();
 FILLCELL_X8 FILLER_77_1249 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X32 FILLER_77_1584 ();
 FILLCELL_X32 FILLER_77_1616 ();
 FILLCELL_X32 FILLER_77_1648 ();
 FILLCELL_X32 FILLER_77_1680 ();
 FILLCELL_X32 FILLER_77_1712 ();
 FILLCELL_X32 FILLER_77_1744 ();
 FILLCELL_X32 FILLER_77_1776 ();
 FILLCELL_X32 FILLER_77_1808 ();
 FILLCELL_X32 FILLER_77_1840 ();
 FILLCELL_X16 FILLER_77_1872 ();
 FILLCELL_X8 FILLER_77_1888 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X32 FILLER_78_952 ();
 FILLCELL_X32 FILLER_78_984 ();
 FILLCELL_X32 FILLER_78_1016 ();
 FILLCELL_X32 FILLER_78_1048 ();
 FILLCELL_X32 FILLER_78_1080 ();
 FILLCELL_X32 FILLER_78_1112 ();
 FILLCELL_X32 FILLER_78_1144 ();
 FILLCELL_X32 FILLER_78_1176 ();
 FILLCELL_X32 FILLER_78_1208 ();
 FILLCELL_X32 FILLER_78_1240 ();
 FILLCELL_X32 FILLER_78_1272 ();
 FILLCELL_X32 FILLER_78_1304 ();
 FILLCELL_X32 FILLER_78_1336 ();
 FILLCELL_X32 FILLER_78_1368 ();
 FILLCELL_X32 FILLER_78_1400 ();
 FILLCELL_X32 FILLER_78_1432 ();
 FILLCELL_X32 FILLER_78_1464 ();
 FILLCELL_X32 FILLER_78_1496 ();
 FILLCELL_X32 FILLER_78_1528 ();
 FILLCELL_X32 FILLER_78_1560 ();
 FILLCELL_X32 FILLER_78_1592 ();
 FILLCELL_X32 FILLER_78_1624 ();
 FILLCELL_X32 FILLER_78_1656 ();
 FILLCELL_X32 FILLER_78_1688 ();
 FILLCELL_X32 FILLER_78_1720 ();
 FILLCELL_X32 FILLER_78_1752 ();
 FILLCELL_X32 FILLER_78_1784 ();
 FILLCELL_X32 FILLER_78_1816 ();
 FILLCELL_X32 FILLER_78_1848 ();
 FILLCELL_X8 FILLER_78_1880 ();
 FILLCELL_X4 FILLER_78_1888 ();
 FILLCELL_X2 FILLER_78_1892 ();
 FILLCELL_X1 FILLER_78_1895 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X32 FILLER_79_961 ();
 FILLCELL_X32 FILLER_79_993 ();
 FILLCELL_X32 FILLER_79_1025 ();
 FILLCELL_X32 FILLER_79_1057 ();
 FILLCELL_X32 FILLER_79_1089 ();
 FILLCELL_X32 FILLER_79_1121 ();
 FILLCELL_X32 FILLER_79_1153 ();
 FILLCELL_X32 FILLER_79_1185 ();
 FILLCELL_X32 FILLER_79_1217 ();
 FILLCELL_X8 FILLER_79_1249 ();
 FILLCELL_X4 FILLER_79_1257 ();
 FILLCELL_X2 FILLER_79_1261 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X32 FILLER_79_1584 ();
 FILLCELL_X32 FILLER_79_1616 ();
 FILLCELL_X32 FILLER_79_1648 ();
 FILLCELL_X32 FILLER_79_1680 ();
 FILLCELL_X32 FILLER_79_1712 ();
 FILLCELL_X32 FILLER_79_1744 ();
 FILLCELL_X32 FILLER_79_1776 ();
 FILLCELL_X32 FILLER_79_1808 ();
 FILLCELL_X32 FILLER_79_1840 ();
 FILLCELL_X16 FILLER_79_1872 ();
 FILLCELL_X8 FILLER_79_1888 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X32 FILLER_80_952 ();
 FILLCELL_X32 FILLER_80_984 ();
 FILLCELL_X32 FILLER_80_1016 ();
 FILLCELL_X32 FILLER_80_1048 ();
 FILLCELL_X32 FILLER_80_1080 ();
 FILLCELL_X32 FILLER_80_1112 ();
 FILLCELL_X32 FILLER_80_1144 ();
 FILLCELL_X32 FILLER_80_1176 ();
 FILLCELL_X32 FILLER_80_1208 ();
 FILLCELL_X32 FILLER_80_1240 ();
 FILLCELL_X32 FILLER_80_1272 ();
 FILLCELL_X32 FILLER_80_1304 ();
 FILLCELL_X32 FILLER_80_1336 ();
 FILLCELL_X32 FILLER_80_1368 ();
 FILLCELL_X32 FILLER_80_1400 ();
 FILLCELL_X32 FILLER_80_1432 ();
 FILLCELL_X32 FILLER_80_1464 ();
 FILLCELL_X32 FILLER_80_1496 ();
 FILLCELL_X32 FILLER_80_1528 ();
 FILLCELL_X32 FILLER_80_1560 ();
 FILLCELL_X32 FILLER_80_1592 ();
 FILLCELL_X32 FILLER_80_1624 ();
 FILLCELL_X32 FILLER_80_1656 ();
 FILLCELL_X32 FILLER_80_1688 ();
 FILLCELL_X32 FILLER_80_1720 ();
 FILLCELL_X32 FILLER_80_1752 ();
 FILLCELL_X32 FILLER_80_1784 ();
 FILLCELL_X32 FILLER_80_1816 ();
 FILLCELL_X32 FILLER_80_1848 ();
 FILLCELL_X8 FILLER_80_1880 ();
 FILLCELL_X4 FILLER_80_1888 ();
 FILLCELL_X2 FILLER_80_1892 ();
 FILLCELL_X1 FILLER_80_1895 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X32 FILLER_81_1584 ();
 FILLCELL_X32 FILLER_81_1616 ();
 FILLCELL_X32 FILLER_81_1648 ();
 FILLCELL_X32 FILLER_81_1680 ();
 FILLCELL_X32 FILLER_81_1712 ();
 FILLCELL_X32 FILLER_81_1744 ();
 FILLCELL_X32 FILLER_81_1776 ();
 FILLCELL_X32 FILLER_81_1808 ();
 FILLCELL_X32 FILLER_81_1840 ();
 FILLCELL_X16 FILLER_81_1872 ();
 FILLCELL_X8 FILLER_81_1888 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X32 FILLER_82_1592 ();
 FILLCELL_X32 FILLER_82_1624 ();
 FILLCELL_X32 FILLER_82_1656 ();
 FILLCELL_X32 FILLER_82_1688 ();
 FILLCELL_X32 FILLER_82_1720 ();
 FILLCELL_X32 FILLER_82_1752 ();
 FILLCELL_X32 FILLER_82_1784 ();
 FILLCELL_X32 FILLER_82_1816 ();
 FILLCELL_X32 FILLER_82_1848 ();
 FILLCELL_X8 FILLER_82_1880 ();
 FILLCELL_X4 FILLER_82_1888 ();
 FILLCELL_X2 FILLER_82_1892 ();
 FILLCELL_X1 FILLER_82_1895 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X32 FILLER_83_1584 ();
 FILLCELL_X32 FILLER_83_1616 ();
 FILLCELL_X32 FILLER_83_1648 ();
 FILLCELL_X32 FILLER_83_1680 ();
 FILLCELL_X32 FILLER_83_1712 ();
 FILLCELL_X32 FILLER_83_1744 ();
 FILLCELL_X32 FILLER_83_1776 ();
 FILLCELL_X32 FILLER_83_1808 ();
 FILLCELL_X32 FILLER_83_1840 ();
 FILLCELL_X16 FILLER_83_1872 ();
 FILLCELL_X8 FILLER_83_1888 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X32 FILLER_84_1592 ();
 FILLCELL_X32 FILLER_84_1624 ();
 FILLCELL_X32 FILLER_84_1656 ();
 FILLCELL_X32 FILLER_84_1688 ();
 FILLCELL_X32 FILLER_84_1720 ();
 FILLCELL_X32 FILLER_84_1752 ();
 FILLCELL_X32 FILLER_84_1784 ();
 FILLCELL_X32 FILLER_84_1816 ();
 FILLCELL_X32 FILLER_84_1848 ();
 FILLCELL_X8 FILLER_84_1880 ();
 FILLCELL_X4 FILLER_84_1888 ();
 FILLCELL_X2 FILLER_84_1892 ();
 FILLCELL_X1 FILLER_84_1895 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X32 FILLER_85_1584 ();
 FILLCELL_X32 FILLER_85_1616 ();
 FILLCELL_X32 FILLER_85_1648 ();
 FILLCELL_X32 FILLER_85_1680 ();
 FILLCELL_X32 FILLER_85_1712 ();
 FILLCELL_X32 FILLER_85_1744 ();
 FILLCELL_X32 FILLER_85_1776 ();
 FILLCELL_X32 FILLER_85_1808 ();
 FILLCELL_X32 FILLER_85_1840 ();
 FILLCELL_X16 FILLER_85_1872 ();
 FILLCELL_X8 FILLER_85_1888 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X32 FILLER_86_1592 ();
 FILLCELL_X32 FILLER_86_1624 ();
 FILLCELL_X32 FILLER_86_1656 ();
 FILLCELL_X32 FILLER_86_1688 ();
 FILLCELL_X32 FILLER_86_1720 ();
 FILLCELL_X32 FILLER_86_1752 ();
 FILLCELL_X32 FILLER_86_1784 ();
 FILLCELL_X32 FILLER_86_1816 ();
 FILLCELL_X32 FILLER_86_1848 ();
 FILLCELL_X8 FILLER_86_1880 ();
 FILLCELL_X4 FILLER_86_1888 ();
 FILLCELL_X2 FILLER_86_1892 ();
 FILLCELL_X1 FILLER_86_1895 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X32 FILLER_87_1584 ();
 FILLCELL_X32 FILLER_87_1616 ();
 FILLCELL_X32 FILLER_87_1648 ();
 FILLCELL_X32 FILLER_87_1680 ();
 FILLCELL_X32 FILLER_87_1712 ();
 FILLCELL_X32 FILLER_87_1744 ();
 FILLCELL_X32 FILLER_87_1776 ();
 FILLCELL_X32 FILLER_87_1808 ();
 FILLCELL_X32 FILLER_87_1840 ();
 FILLCELL_X16 FILLER_87_1872 ();
 FILLCELL_X8 FILLER_87_1888 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X32 FILLER_88_1592 ();
 FILLCELL_X32 FILLER_88_1624 ();
 FILLCELL_X32 FILLER_88_1656 ();
 FILLCELL_X32 FILLER_88_1688 ();
 FILLCELL_X32 FILLER_88_1720 ();
 FILLCELL_X32 FILLER_88_1752 ();
 FILLCELL_X32 FILLER_88_1784 ();
 FILLCELL_X32 FILLER_88_1816 ();
 FILLCELL_X32 FILLER_88_1848 ();
 FILLCELL_X8 FILLER_88_1880 ();
 FILLCELL_X4 FILLER_88_1888 ();
 FILLCELL_X2 FILLER_88_1892 ();
 FILLCELL_X1 FILLER_88_1895 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X32 FILLER_89_1584 ();
 FILLCELL_X32 FILLER_89_1616 ();
 FILLCELL_X32 FILLER_89_1648 ();
 FILLCELL_X32 FILLER_89_1680 ();
 FILLCELL_X32 FILLER_89_1712 ();
 FILLCELL_X32 FILLER_89_1744 ();
 FILLCELL_X32 FILLER_89_1776 ();
 FILLCELL_X32 FILLER_89_1808 ();
 FILLCELL_X32 FILLER_89_1840 ();
 FILLCELL_X16 FILLER_89_1872 ();
 FILLCELL_X8 FILLER_89_1888 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X32 FILLER_90_1592 ();
 FILLCELL_X32 FILLER_90_1624 ();
 FILLCELL_X32 FILLER_90_1656 ();
 FILLCELL_X32 FILLER_90_1688 ();
 FILLCELL_X32 FILLER_90_1720 ();
 FILLCELL_X32 FILLER_90_1752 ();
 FILLCELL_X32 FILLER_90_1784 ();
 FILLCELL_X32 FILLER_90_1816 ();
 FILLCELL_X32 FILLER_90_1848 ();
 FILLCELL_X8 FILLER_90_1880 ();
 FILLCELL_X4 FILLER_90_1888 ();
 FILLCELL_X2 FILLER_90_1892 ();
 FILLCELL_X1 FILLER_90_1895 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X32 FILLER_91_1584 ();
 FILLCELL_X32 FILLER_91_1616 ();
 FILLCELL_X32 FILLER_91_1648 ();
 FILLCELL_X32 FILLER_91_1680 ();
 FILLCELL_X32 FILLER_91_1712 ();
 FILLCELL_X32 FILLER_91_1744 ();
 FILLCELL_X32 FILLER_91_1776 ();
 FILLCELL_X32 FILLER_91_1808 ();
 FILLCELL_X32 FILLER_91_1840 ();
 FILLCELL_X16 FILLER_91_1872 ();
 FILLCELL_X8 FILLER_91_1888 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X32 FILLER_92_1592 ();
 FILLCELL_X32 FILLER_92_1624 ();
 FILLCELL_X32 FILLER_92_1656 ();
 FILLCELL_X32 FILLER_92_1688 ();
 FILLCELL_X32 FILLER_92_1720 ();
 FILLCELL_X32 FILLER_92_1752 ();
 FILLCELL_X32 FILLER_92_1784 ();
 FILLCELL_X32 FILLER_92_1816 ();
 FILLCELL_X32 FILLER_92_1848 ();
 FILLCELL_X8 FILLER_92_1880 ();
 FILLCELL_X4 FILLER_92_1888 ();
 FILLCELL_X2 FILLER_92_1892 ();
 FILLCELL_X1 FILLER_92_1895 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X32 FILLER_93_1584 ();
 FILLCELL_X32 FILLER_93_1616 ();
 FILLCELL_X32 FILLER_93_1648 ();
 FILLCELL_X32 FILLER_93_1680 ();
 FILLCELL_X32 FILLER_93_1712 ();
 FILLCELL_X32 FILLER_93_1744 ();
 FILLCELL_X32 FILLER_93_1776 ();
 FILLCELL_X32 FILLER_93_1808 ();
 FILLCELL_X32 FILLER_93_1840 ();
 FILLCELL_X16 FILLER_93_1872 ();
 FILLCELL_X8 FILLER_93_1888 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X32 FILLER_94_1592 ();
 FILLCELL_X32 FILLER_94_1624 ();
 FILLCELL_X32 FILLER_94_1656 ();
 FILLCELL_X32 FILLER_94_1688 ();
 FILLCELL_X32 FILLER_94_1720 ();
 FILLCELL_X32 FILLER_94_1752 ();
 FILLCELL_X32 FILLER_94_1784 ();
 FILLCELL_X32 FILLER_94_1816 ();
 FILLCELL_X32 FILLER_94_1848 ();
 FILLCELL_X8 FILLER_94_1880 ();
 FILLCELL_X4 FILLER_94_1888 ();
 FILLCELL_X2 FILLER_94_1892 ();
 FILLCELL_X1 FILLER_94_1895 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X32 FILLER_95_961 ();
 FILLCELL_X32 FILLER_95_993 ();
 FILLCELL_X32 FILLER_95_1025 ();
 FILLCELL_X32 FILLER_95_1057 ();
 FILLCELL_X32 FILLER_95_1089 ();
 FILLCELL_X32 FILLER_95_1121 ();
 FILLCELL_X32 FILLER_95_1153 ();
 FILLCELL_X32 FILLER_95_1185 ();
 FILLCELL_X32 FILLER_95_1217 ();
 FILLCELL_X8 FILLER_95_1249 ();
 FILLCELL_X4 FILLER_95_1257 ();
 FILLCELL_X2 FILLER_95_1261 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X32 FILLER_95_1584 ();
 FILLCELL_X32 FILLER_95_1616 ();
 FILLCELL_X32 FILLER_95_1648 ();
 FILLCELL_X32 FILLER_95_1680 ();
 FILLCELL_X32 FILLER_95_1712 ();
 FILLCELL_X32 FILLER_95_1744 ();
 FILLCELL_X32 FILLER_95_1776 ();
 FILLCELL_X32 FILLER_95_1808 ();
 FILLCELL_X32 FILLER_95_1840 ();
 FILLCELL_X16 FILLER_95_1872 ();
 FILLCELL_X8 FILLER_95_1888 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X32 FILLER_96_1592 ();
 FILLCELL_X32 FILLER_96_1624 ();
 FILLCELL_X32 FILLER_96_1656 ();
 FILLCELL_X32 FILLER_96_1688 ();
 FILLCELL_X32 FILLER_96_1720 ();
 FILLCELL_X32 FILLER_96_1752 ();
 FILLCELL_X32 FILLER_96_1784 ();
 FILLCELL_X32 FILLER_96_1816 ();
 FILLCELL_X32 FILLER_96_1848 ();
 FILLCELL_X8 FILLER_96_1880 ();
 FILLCELL_X4 FILLER_96_1888 ();
 FILLCELL_X2 FILLER_96_1892 ();
 FILLCELL_X1 FILLER_96_1895 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X32 FILLER_97_961 ();
 FILLCELL_X32 FILLER_97_993 ();
 FILLCELL_X32 FILLER_97_1025 ();
 FILLCELL_X32 FILLER_97_1057 ();
 FILLCELL_X32 FILLER_97_1089 ();
 FILLCELL_X32 FILLER_97_1121 ();
 FILLCELL_X32 FILLER_97_1153 ();
 FILLCELL_X32 FILLER_97_1185 ();
 FILLCELL_X32 FILLER_97_1217 ();
 FILLCELL_X8 FILLER_97_1249 ();
 FILLCELL_X4 FILLER_97_1257 ();
 FILLCELL_X2 FILLER_97_1261 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X32 FILLER_97_1584 ();
 FILLCELL_X32 FILLER_97_1616 ();
 FILLCELL_X32 FILLER_97_1648 ();
 FILLCELL_X32 FILLER_97_1680 ();
 FILLCELL_X32 FILLER_97_1712 ();
 FILLCELL_X32 FILLER_97_1744 ();
 FILLCELL_X32 FILLER_97_1776 ();
 FILLCELL_X32 FILLER_97_1808 ();
 FILLCELL_X32 FILLER_97_1840 ();
 FILLCELL_X16 FILLER_97_1872 ();
 FILLCELL_X8 FILLER_97_1888 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X32 FILLER_98_1304 ();
 FILLCELL_X32 FILLER_98_1336 ();
 FILLCELL_X32 FILLER_98_1368 ();
 FILLCELL_X32 FILLER_98_1400 ();
 FILLCELL_X32 FILLER_98_1432 ();
 FILLCELL_X32 FILLER_98_1464 ();
 FILLCELL_X32 FILLER_98_1496 ();
 FILLCELL_X32 FILLER_98_1528 ();
 FILLCELL_X32 FILLER_98_1560 ();
 FILLCELL_X32 FILLER_98_1592 ();
 FILLCELL_X32 FILLER_98_1624 ();
 FILLCELL_X32 FILLER_98_1656 ();
 FILLCELL_X32 FILLER_98_1688 ();
 FILLCELL_X32 FILLER_98_1720 ();
 FILLCELL_X32 FILLER_98_1752 ();
 FILLCELL_X32 FILLER_98_1784 ();
 FILLCELL_X32 FILLER_98_1816 ();
 FILLCELL_X32 FILLER_98_1848 ();
 FILLCELL_X8 FILLER_98_1880 ();
 FILLCELL_X4 FILLER_98_1888 ();
 FILLCELL_X2 FILLER_98_1892 ();
 FILLCELL_X1 FILLER_98_1895 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X32 FILLER_99_1584 ();
 FILLCELL_X32 FILLER_99_1616 ();
 FILLCELL_X32 FILLER_99_1648 ();
 FILLCELL_X32 FILLER_99_1680 ();
 FILLCELL_X32 FILLER_99_1712 ();
 FILLCELL_X32 FILLER_99_1744 ();
 FILLCELL_X32 FILLER_99_1776 ();
 FILLCELL_X32 FILLER_99_1808 ();
 FILLCELL_X32 FILLER_99_1840 ();
 FILLCELL_X16 FILLER_99_1872 ();
 FILLCELL_X8 FILLER_99_1888 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X32 FILLER_100_952 ();
 FILLCELL_X32 FILLER_100_984 ();
 FILLCELL_X32 FILLER_100_1016 ();
 FILLCELL_X32 FILLER_100_1048 ();
 FILLCELL_X32 FILLER_100_1080 ();
 FILLCELL_X32 FILLER_100_1112 ();
 FILLCELL_X32 FILLER_100_1144 ();
 FILLCELL_X32 FILLER_100_1176 ();
 FILLCELL_X32 FILLER_100_1208 ();
 FILLCELL_X32 FILLER_100_1240 ();
 FILLCELL_X32 FILLER_100_1272 ();
 FILLCELL_X32 FILLER_100_1304 ();
 FILLCELL_X32 FILLER_100_1336 ();
 FILLCELL_X32 FILLER_100_1368 ();
 FILLCELL_X32 FILLER_100_1400 ();
 FILLCELL_X32 FILLER_100_1432 ();
 FILLCELL_X32 FILLER_100_1464 ();
 FILLCELL_X32 FILLER_100_1496 ();
 FILLCELL_X32 FILLER_100_1528 ();
 FILLCELL_X32 FILLER_100_1560 ();
 FILLCELL_X32 FILLER_100_1592 ();
 FILLCELL_X32 FILLER_100_1624 ();
 FILLCELL_X32 FILLER_100_1656 ();
 FILLCELL_X32 FILLER_100_1688 ();
 FILLCELL_X32 FILLER_100_1720 ();
 FILLCELL_X32 FILLER_100_1752 ();
 FILLCELL_X32 FILLER_100_1784 ();
 FILLCELL_X32 FILLER_100_1816 ();
 FILLCELL_X32 FILLER_100_1848 ();
 FILLCELL_X8 FILLER_100_1880 ();
 FILLCELL_X4 FILLER_100_1888 ();
 FILLCELL_X2 FILLER_100_1892 ();
 FILLCELL_X1 FILLER_100_1895 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X32 FILLER_101_1584 ();
 FILLCELL_X32 FILLER_101_1616 ();
 FILLCELL_X32 FILLER_101_1648 ();
 FILLCELL_X32 FILLER_101_1680 ();
 FILLCELL_X32 FILLER_101_1712 ();
 FILLCELL_X32 FILLER_101_1744 ();
 FILLCELL_X32 FILLER_101_1776 ();
 FILLCELL_X32 FILLER_101_1808 ();
 FILLCELL_X32 FILLER_101_1840 ();
 FILLCELL_X16 FILLER_101_1872 ();
 FILLCELL_X8 FILLER_101_1888 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X32 FILLER_102_1304 ();
 FILLCELL_X32 FILLER_102_1336 ();
 FILLCELL_X32 FILLER_102_1368 ();
 FILLCELL_X32 FILLER_102_1400 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X32 FILLER_102_1496 ();
 FILLCELL_X32 FILLER_102_1528 ();
 FILLCELL_X32 FILLER_102_1560 ();
 FILLCELL_X32 FILLER_102_1592 ();
 FILLCELL_X32 FILLER_102_1624 ();
 FILLCELL_X32 FILLER_102_1656 ();
 FILLCELL_X32 FILLER_102_1688 ();
 FILLCELL_X32 FILLER_102_1720 ();
 FILLCELL_X32 FILLER_102_1752 ();
 FILLCELL_X32 FILLER_102_1784 ();
 FILLCELL_X32 FILLER_102_1816 ();
 FILLCELL_X32 FILLER_102_1848 ();
 FILLCELL_X8 FILLER_102_1880 ();
 FILLCELL_X4 FILLER_102_1888 ();
 FILLCELL_X2 FILLER_102_1892 ();
 FILLCELL_X1 FILLER_102_1895 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X32 FILLER_103_1584 ();
 FILLCELL_X32 FILLER_103_1616 ();
 FILLCELL_X32 FILLER_103_1648 ();
 FILLCELL_X32 FILLER_103_1680 ();
 FILLCELL_X32 FILLER_103_1712 ();
 FILLCELL_X32 FILLER_103_1744 ();
 FILLCELL_X32 FILLER_103_1776 ();
 FILLCELL_X32 FILLER_103_1808 ();
 FILLCELL_X32 FILLER_103_1840 ();
 FILLCELL_X16 FILLER_103_1872 ();
 FILLCELL_X8 FILLER_103_1888 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X32 FILLER_104_1304 ();
 FILLCELL_X32 FILLER_104_1336 ();
 FILLCELL_X32 FILLER_104_1368 ();
 FILLCELL_X32 FILLER_104_1400 ();
 FILLCELL_X32 FILLER_104_1432 ();
 FILLCELL_X32 FILLER_104_1464 ();
 FILLCELL_X32 FILLER_104_1496 ();
 FILLCELL_X32 FILLER_104_1528 ();
 FILLCELL_X32 FILLER_104_1560 ();
 FILLCELL_X32 FILLER_104_1592 ();
 FILLCELL_X32 FILLER_104_1624 ();
 FILLCELL_X32 FILLER_104_1656 ();
 FILLCELL_X32 FILLER_104_1688 ();
 FILLCELL_X32 FILLER_104_1720 ();
 FILLCELL_X32 FILLER_104_1752 ();
 FILLCELL_X32 FILLER_104_1784 ();
 FILLCELL_X32 FILLER_104_1816 ();
 FILLCELL_X32 FILLER_104_1848 ();
 FILLCELL_X8 FILLER_104_1880 ();
 FILLCELL_X4 FILLER_104_1888 ();
 FILLCELL_X2 FILLER_104_1892 ();
 FILLCELL_X1 FILLER_104_1895 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X16 FILLER_105_929 ();
 FILLCELL_X4 FILLER_105_945 ();
 FILLCELL_X2 FILLER_105_949 ();
 FILLCELL_X32 FILLER_105_976 ();
 FILLCELL_X32 FILLER_105_1008 ();
 FILLCELL_X32 FILLER_105_1040 ();
 FILLCELL_X32 FILLER_105_1072 ();
 FILLCELL_X32 FILLER_105_1104 ();
 FILLCELL_X32 FILLER_105_1136 ();
 FILLCELL_X32 FILLER_105_1168 ();
 FILLCELL_X32 FILLER_105_1200 ();
 FILLCELL_X16 FILLER_105_1232 ();
 FILLCELL_X8 FILLER_105_1248 ();
 FILLCELL_X4 FILLER_105_1256 ();
 FILLCELL_X2 FILLER_105_1260 ();
 FILLCELL_X1 FILLER_105_1262 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X32 FILLER_105_1584 ();
 FILLCELL_X32 FILLER_105_1616 ();
 FILLCELL_X32 FILLER_105_1648 ();
 FILLCELL_X32 FILLER_105_1680 ();
 FILLCELL_X32 FILLER_105_1712 ();
 FILLCELL_X32 FILLER_105_1744 ();
 FILLCELL_X32 FILLER_105_1776 ();
 FILLCELL_X32 FILLER_105_1808 ();
 FILLCELL_X32 FILLER_105_1840 ();
 FILLCELL_X16 FILLER_105_1872 ();
 FILLCELL_X8 FILLER_105_1888 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X32 FILLER_106_1304 ();
 FILLCELL_X32 FILLER_106_1336 ();
 FILLCELL_X32 FILLER_106_1368 ();
 FILLCELL_X32 FILLER_106_1400 ();
 FILLCELL_X32 FILLER_106_1432 ();
 FILLCELL_X32 FILLER_106_1464 ();
 FILLCELL_X32 FILLER_106_1496 ();
 FILLCELL_X32 FILLER_106_1528 ();
 FILLCELL_X32 FILLER_106_1560 ();
 FILLCELL_X32 FILLER_106_1592 ();
 FILLCELL_X32 FILLER_106_1624 ();
 FILLCELL_X32 FILLER_106_1656 ();
 FILLCELL_X32 FILLER_106_1688 ();
 FILLCELL_X32 FILLER_106_1720 ();
 FILLCELL_X32 FILLER_106_1752 ();
 FILLCELL_X32 FILLER_106_1784 ();
 FILLCELL_X32 FILLER_106_1816 ();
 FILLCELL_X32 FILLER_106_1848 ();
 FILLCELL_X8 FILLER_106_1880 ();
 FILLCELL_X4 FILLER_106_1888 ();
 FILLCELL_X2 FILLER_106_1892 ();
 FILLCELL_X1 FILLER_106_1895 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X16 FILLER_107_961 ();
 FILLCELL_X8 FILLER_107_977 ();
 FILLCELL_X4 FILLER_107_985 ();
 FILLCELL_X1 FILLER_107_989 ();
 FILLCELL_X32 FILLER_107_1003 ();
 FILLCELL_X32 FILLER_107_1035 ();
 FILLCELL_X32 FILLER_107_1067 ();
 FILLCELL_X32 FILLER_107_1099 ();
 FILLCELL_X32 FILLER_107_1131 ();
 FILLCELL_X32 FILLER_107_1163 ();
 FILLCELL_X32 FILLER_107_1195 ();
 FILLCELL_X32 FILLER_107_1227 ();
 FILLCELL_X4 FILLER_107_1259 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X32 FILLER_107_1584 ();
 FILLCELL_X32 FILLER_107_1616 ();
 FILLCELL_X32 FILLER_107_1648 ();
 FILLCELL_X32 FILLER_107_1680 ();
 FILLCELL_X32 FILLER_107_1712 ();
 FILLCELL_X32 FILLER_107_1744 ();
 FILLCELL_X32 FILLER_107_1776 ();
 FILLCELL_X32 FILLER_107_1808 ();
 FILLCELL_X32 FILLER_107_1840 ();
 FILLCELL_X16 FILLER_107_1872 ();
 FILLCELL_X8 FILLER_107_1888 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X16 FILLER_108_792 ();
 FILLCELL_X2 FILLER_108_808 ();
 FILLCELL_X1 FILLER_108_810 ();
 FILLCELL_X16 FILLER_108_836 ();
 FILLCELL_X8 FILLER_108_852 ();
 FILLCELL_X8 FILLER_108_873 ();
 FILLCELL_X2 FILLER_108_881 ();
 FILLCELL_X1 FILLER_108_883 ();
 FILLCELL_X32 FILLER_108_909 ();
 FILLCELL_X32 FILLER_108_941 ();
 FILLCELL_X32 FILLER_108_973 ();
 FILLCELL_X32 FILLER_108_1005 ();
 FILLCELL_X32 FILLER_108_1037 ();
 FILLCELL_X32 FILLER_108_1069 ();
 FILLCELL_X32 FILLER_108_1101 ();
 FILLCELL_X32 FILLER_108_1133 ();
 FILLCELL_X32 FILLER_108_1165 ();
 FILLCELL_X32 FILLER_108_1197 ();
 FILLCELL_X32 FILLER_108_1229 ();
 FILLCELL_X32 FILLER_108_1261 ();
 FILLCELL_X32 FILLER_108_1293 ();
 FILLCELL_X32 FILLER_108_1325 ();
 FILLCELL_X32 FILLER_108_1357 ();
 FILLCELL_X32 FILLER_108_1389 ();
 FILLCELL_X32 FILLER_108_1421 ();
 FILLCELL_X32 FILLER_108_1453 ();
 FILLCELL_X32 FILLER_108_1485 ();
 FILLCELL_X32 FILLER_108_1517 ();
 FILLCELL_X32 FILLER_108_1549 ();
 FILLCELL_X32 FILLER_108_1581 ();
 FILLCELL_X32 FILLER_108_1613 ();
 FILLCELL_X32 FILLER_108_1645 ();
 FILLCELL_X32 FILLER_108_1677 ();
 FILLCELL_X32 FILLER_108_1709 ();
 FILLCELL_X32 FILLER_108_1741 ();
 FILLCELL_X32 FILLER_108_1773 ();
 FILLCELL_X32 FILLER_108_1805 ();
 FILLCELL_X32 FILLER_108_1837 ();
 FILLCELL_X16 FILLER_108_1869 ();
 FILLCELL_X8 FILLER_108_1885 ();
 FILLCELL_X1 FILLER_108_1893 ();
 FILLCELL_X1 FILLER_108_1895 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X2 FILLER_109_833 ();
 FILLCELL_X1 FILLER_109_835 ();
 FILLCELL_X32 FILLER_109_849 ();
 FILLCELL_X4 FILLER_109_881 ();
 FILLCELL_X1 FILLER_109_885 ();
 FILLCELL_X32 FILLER_109_899 ();
 FILLCELL_X8 FILLER_109_931 ();
 FILLCELL_X4 FILLER_109_939 ();
 FILLCELL_X2 FILLER_109_943 ();
 FILLCELL_X1 FILLER_109_945 ();
 FILLCELL_X1 FILLER_109_951 ();
 FILLCELL_X8 FILLER_109_961 ();
 FILLCELL_X4 FILLER_109_969 ();
 FILLCELL_X2 FILLER_109_973 ();
 FILLCELL_X1 FILLER_109_975 ();
 FILLCELL_X32 FILLER_109_1001 ();
 FILLCELL_X32 FILLER_109_1033 ();
 FILLCELL_X32 FILLER_109_1065 ();
 FILLCELL_X32 FILLER_109_1097 ();
 FILLCELL_X32 FILLER_109_1129 ();
 FILLCELL_X32 FILLER_109_1161 ();
 FILLCELL_X32 FILLER_109_1193 ();
 FILLCELL_X32 FILLER_109_1225 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X32 FILLER_109_1584 ();
 FILLCELL_X32 FILLER_109_1616 ();
 FILLCELL_X32 FILLER_109_1648 ();
 FILLCELL_X32 FILLER_109_1680 ();
 FILLCELL_X32 FILLER_109_1712 ();
 FILLCELL_X32 FILLER_109_1744 ();
 FILLCELL_X32 FILLER_109_1776 ();
 FILLCELL_X32 FILLER_109_1808 ();
 FILLCELL_X32 FILLER_109_1840 ();
 FILLCELL_X16 FILLER_109_1872 ();
 FILLCELL_X8 FILLER_109_1888 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X16 FILLER_110_792 ();
 FILLCELL_X2 FILLER_110_808 ();
 FILLCELL_X32 FILLER_110_823 ();
 FILLCELL_X32 FILLER_110_855 ();
 FILLCELL_X32 FILLER_110_887 ();
 FILLCELL_X16 FILLER_110_919 ();
 FILLCELL_X8 FILLER_110_935 ();
 FILLCELL_X2 FILLER_110_943 ();
 FILLCELL_X1 FILLER_110_945 ();
 FILLCELL_X8 FILLER_110_962 ();
 FILLCELL_X4 FILLER_110_970 ();
 FILLCELL_X16 FILLER_110_979 ();
 FILLCELL_X1 FILLER_110_995 ();
 FILLCELL_X32 FILLER_110_1009 ();
 FILLCELL_X32 FILLER_110_1041 ();
 FILLCELL_X32 FILLER_110_1073 ();
 FILLCELL_X32 FILLER_110_1105 ();
 FILLCELL_X32 FILLER_110_1137 ();
 FILLCELL_X32 FILLER_110_1169 ();
 FILLCELL_X32 FILLER_110_1201 ();
 FILLCELL_X32 FILLER_110_1233 ();
 FILLCELL_X32 FILLER_110_1265 ();
 FILLCELL_X32 FILLER_110_1297 ();
 FILLCELL_X32 FILLER_110_1329 ();
 FILLCELL_X32 FILLER_110_1361 ();
 FILLCELL_X32 FILLER_110_1393 ();
 FILLCELL_X32 FILLER_110_1425 ();
 FILLCELL_X32 FILLER_110_1457 ();
 FILLCELL_X32 FILLER_110_1489 ();
 FILLCELL_X32 FILLER_110_1521 ();
 FILLCELL_X32 FILLER_110_1553 ();
 FILLCELL_X32 FILLER_110_1585 ();
 FILLCELL_X32 FILLER_110_1617 ();
 FILLCELL_X32 FILLER_110_1649 ();
 FILLCELL_X32 FILLER_110_1681 ();
 FILLCELL_X32 FILLER_110_1713 ();
 FILLCELL_X32 FILLER_110_1745 ();
 FILLCELL_X32 FILLER_110_1777 ();
 FILLCELL_X32 FILLER_110_1809 ();
 FILLCELL_X32 FILLER_110_1841 ();
 FILLCELL_X16 FILLER_110_1873 ();
 FILLCELL_X4 FILLER_110_1889 ();
 FILLCELL_X1 FILLER_110_1893 ();
 FILLCELL_X1 FILLER_110_1895 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X4 FILLER_111_801 ();
 FILLCELL_X2 FILLER_111_805 ();
 FILLCELL_X1 FILLER_111_807 ();
 FILLCELL_X32 FILLER_111_815 ();
 FILLCELL_X32 FILLER_111_847 ();
 FILLCELL_X32 FILLER_111_879 ();
 FILLCELL_X32 FILLER_111_911 ();
 FILLCELL_X8 FILLER_111_943 ();
 FILLCELL_X8 FILLER_111_956 ();
 FILLCELL_X4 FILLER_111_964 ();
 FILLCELL_X2 FILLER_111_968 ();
 FILLCELL_X1 FILLER_111_970 ();
 FILLCELL_X32 FILLER_111_980 ();
 FILLCELL_X32 FILLER_111_1012 ();
 FILLCELL_X32 FILLER_111_1044 ();
 FILLCELL_X32 FILLER_111_1076 ();
 FILLCELL_X32 FILLER_111_1108 ();
 FILLCELL_X32 FILLER_111_1140 ();
 FILLCELL_X32 FILLER_111_1172 ();
 FILLCELL_X32 FILLER_111_1204 ();
 FILLCELL_X16 FILLER_111_1236 ();
 FILLCELL_X8 FILLER_111_1252 ();
 FILLCELL_X2 FILLER_111_1260 ();
 FILLCELL_X1 FILLER_111_1262 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X32 FILLER_111_1584 ();
 FILLCELL_X32 FILLER_111_1616 ();
 FILLCELL_X32 FILLER_111_1648 ();
 FILLCELL_X32 FILLER_111_1680 ();
 FILLCELL_X32 FILLER_111_1712 ();
 FILLCELL_X32 FILLER_111_1744 ();
 FILLCELL_X32 FILLER_111_1776 ();
 FILLCELL_X32 FILLER_111_1808 ();
 FILLCELL_X32 FILLER_111_1840 ();
 FILLCELL_X16 FILLER_111_1872 ();
 FILLCELL_X8 FILLER_111_1888 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X16 FILLER_112_856 ();
 FILLCELL_X8 FILLER_112_872 ();
 FILLCELL_X4 FILLER_112_880 ();
 FILLCELL_X2 FILLER_112_884 ();
 FILLCELL_X1 FILLER_112_886 ();
 FILLCELL_X16 FILLER_112_893 ();
 FILLCELL_X2 FILLER_112_909 ();
 FILLCELL_X4 FILLER_112_915 ();
 FILLCELL_X32 FILLER_112_929 ();
 FILLCELL_X4 FILLER_112_961 ();
 FILLCELL_X2 FILLER_112_965 ();
 FILLCELL_X1 FILLER_112_971 ();
 FILLCELL_X32 FILLER_112_981 ();
 FILLCELL_X32 FILLER_112_1013 ();
 FILLCELL_X32 FILLER_112_1045 ();
 FILLCELL_X32 FILLER_112_1077 ();
 FILLCELL_X32 FILLER_112_1109 ();
 FILLCELL_X32 FILLER_112_1141 ();
 FILLCELL_X32 FILLER_112_1173 ();
 FILLCELL_X32 FILLER_112_1205 ();
 FILLCELL_X32 FILLER_112_1237 ();
 FILLCELL_X32 FILLER_112_1269 ();
 FILLCELL_X32 FILLER_112_1301 ();
 FILLCELL_X32 FILLER_112_1333 ();
 FILLCELL_X32 FILLER_112_1365 ();
 FILLCELL_X32 FILLER_112_1397 ();
 FILLCELL_X32 FILLER_112_1429 ();
 FILLCELL_X32 FILLER_112_1461 ();
 FILLCELL_X32 FILLER_112_1493 ();
 FILLCELL_X32 FILLER_112_1525 ();
 FILLCELL_X32 FILLER_112_1557 ();
 FILLCELL_X32 FILLER_112_1589 ();
 FILLCELL_X32 FILLER_112_1621 ();
 FILLCELL_X32 FILLER_112_1653 ();
 FILLCELL_X32 FILLER_112_1685 ();
 FILLCELL_X32 FILLER_112_1717 ();
 FILLCELL_X32 FILLER_112_1749 ();
 FILLCELL_X32 FILLER_112_1781 ();
 FILLCELL_X32 FILLER_112_1813 ();
 FILLCELL_X16 FILLER_112_1845 ();
 FILLCELL_X4 FILLER_112_1861 ();
 FILLCELL_X2 FILLER_112_1865 ();
 FILLCELL_X16 FILLER_112_1870 ();
 FILLCELL_X8 FILLER_112_1886 ();
 FILLCELL_X1 FILLER_112_1895 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X32 FILLER_113_833 ();
 FILLCELL_X16 FILLER_113_865 ();
 FILLCELL_X8 FILLER_113_897 ();
 FILLCELL_X4 FILLER_113_905 ();
 FILLCELL_X1 FILLER_113_909 ();
 FILLCELL_X8 FILLER_113_926 ();
 FILLCELL_X4 FILLER_113_934 ();
 FILLCELL_X32 FILLER_113_940 ();
 FILLCELL_X8 FILLER_113_972 ();
 FILLCELL_X4 FILLER_113_980 ();
 FILLCELL_X2 FILLER_113_984 ();
 FILLCELL_X8 FILLER_113_1018 ();
 FILLCELL_X4 FILLER_113_1026 ();
 FILLCELL_X2 FILLER_113_1036 ();
 FILLCELL_X8 FILLER_113_1044 ();
 FILLCELL_X1 FILLER_113_1052 ();
 FILLCELL_X8 FILLER_113_1056 ();
 FILLCELL_X4 FILLER_113_1064 ();
 FILLCELL_X1 FILLER_113_1068 ();
 FILLCELL_X32 FILLER_113_1072 ();
 FILLCELL_X1 FILLER_113_1104 ();
 FILLCELL_X16 FILLER_113_1108 ();
 FILLCELL_X8 FILLER_113_1124 ();
 FILLCELL_X2 FILLER_113_1132 ();
 FILLCELL_X2 FILLER_113_1140 ();
 FILLCELL_X2 FILLER_113_1146 ();
 FILLCELL_X32 FILLER_113_1162 ();
 FILLCELL_X1 FILLER_113_1194 ();
 FILLCELL_X2 FILLER_113_1199 ();
 FILLCELL_X2 FILLER_113_1206 ();
 FILLCELL_X32 FILLER_113_1221 ();
 FILLCELL_X8 FILLER_113_1253 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X32 FILLER_113_1552 ();
 FILLCELL_X32 FILLER_113_1584 ();
 FILLCELL_X32 FILLER_113_1616 ();
 FILLCELL_X32 FILLER_113_1648 ();
 FILLCELL_X32 FILLER_113_1680 ();
 FILLCELL_X32 FILLER_113_1712 ();
 FILLCELL_X32 FILLER_113_1744 ();
 FILLCELL_X32 FILLER_113_1776 ();
 FILLCELL_X32 FILLER_113_1808 ();
 FILLCELL_X32 FILLER_113_1840 ();
 FILLCELL_X16 FILLER_113_1872 ();
 FILLCELL_X4 FILLER_113_1888 ();
 FILLCELL_X1 FILLER_113_1892 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X8 FILLER_114_856 ();
 FILLCELL_X4 FILLER_114_864 ();
 FILLCELL_X8 FILLER_114_871 ();
 FILLCELL_X2 FILLER_114_879 ();
 FILLCELL_X4 FILLER_114_883 ();
 FILLCELL_X2 FILLER_114_887 ();
 FILLCELL_X32 FILLER_114_898 ();
 FILLCELL_X2 FILLER_114_930 ();
 FILLCELL_X2 FILLER_114_950 ();
 FILLCELL_X1 FILLER_114_952 ();
 FILLCELL_X4 FILLER_114_956 ();
 FILLCELL_X2 FILLER_114_960 ();
 FILLCELL_X16 FILLER_114_976 ();
 FILLCELL_X8 FILLER_114_992 ();
 FILLCELL_X4 FILLER_114_1000 ();
 FILLCELL_X2 FILLER_114_1004 ();
 FILLCELL_X1 FILLER_114_1010 ();
 FILLCELL_X8 FILLER_114_1014 ();
 FILLCELL_X2 FILLER_114_1022 ();
 FILLCELL_X1 FILLER_114_1024 ();
 FILLCELL_X4 FILLER_114_1027 ();
 FILLCELL_X8 FILLER_114_1047 ();
 FILLCELL_X2 FILLER_114_1055 ();
 FILLCELL_X8 FILLER_114_1073 ();
 FILLCELL_X1 FILLER_114_1081 ();
 FILLCELL_X4 FILLER_114_1088 ();
 FILLCELL_X16 FILLER_114_1095 ();
 FILLCELL_X4 FILLER_114_1111 ();
 FILLCELL_X4 FILLER_114_1118 ();
 FILLCELL_X2 FILLER_114_1122 ();
 FILLCELL_X1 FILLER_114_1124 ();
 FILLCELL_X2 FILLER_114_1144 ();
 FILLCELL_X1 FILLER_114_1146 ();
 FILLCELL_X4 FILLER_114_1149 ();
 FILLCELL_X2 FILLER_114_1153 ();
 FILLCELL_X1 FILLER_114_1155 ();
 FILLCELL_X4 FILLER_114_1166 ();
 FILLCELL_X2 FILLER_114_1170 ();
 FILLCELL_X1 FILLER_114_1172 ();
 FILLCELL_X32 FILLER_114_1177 ();
 FILLCELL_X32 FILLER_114_1209 ();
 FILLCELL_X32 FILLER_114_1241 ();
 FILLCELL_X32 FILLER_114_1273 ();
 FILLCELL_X32 FILLER_114_1305 ();
 FILLCELL_X32 FILLER_114_1337 ();
 FILLCELL_X32 FILLER_114_1369 ();
 FILLCELL_X32 FILLER_114_1401 ();
 FILLCELL_X32 FILLER_114_1433 ();
 FILLCELL_X32 FILLER_114_1465 ();
 FILLCELL_X32 FILLER_114_1497 ();
 FILLCELL_X32 FILLER_114_1529 ();
 FILLCELL_X32 FILLER_114_1561 ();
 FILLCELL_X32 FILLER_114_1593 ();
 FILLCELL_X32 FILLER_114_1625 ();
 FILLCELL_X32 FILLER_114_1657 ();
 FILLCELL_X32 FILLER_114_1689 ();
 FILLCELL_X32 FILLER_114_1721 ();
 FILLCELL_X32 FILLER_114_1753 ();
 FILLCELL_X32 FILLER_114_1785 ();
 FILLCELL_X32 FILLER_114_1817 ();
 FILLCELL_X4 FILLER_114_1849 ();
 FILLCELL_X4 FILLER_114_1878 ();
 FILLCELL_X2 FILLER_114_1882 ();
 FILLCELL_X4 FILLER_114_1887 ();
 FILLCELL_X2 FILLER_114_1891 ();
 FILLCELL_X1 FILLER_114_1893 ();
 FILLCELL_X1 FILLER_114_1895 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X16 FILLER_115_801 ();
 FILLCELL_X4 FILLER_115_817 ();
 FILLCELL_X2 FILLER_115_821 ();
 FILLCELL_X16 FILLER_115_828 ();
 FILLCELL_X2 FILLER_115_844 ();
 FILLCELL_X1 FILLER_115_846 ();
 FILLCELL_X2 FILLER_115_849 ();
 FILLCELL_X1 FILLER_115_851 ();
 FILLCELL_X16 FILLER_115_870 ();
 FILLCELL_X2 FILLER_115_886 ();
 FILLCELL_X16 FILLER_115_891 ();
 FILLCELL_X8 FILLER_115_907 ();
 FILLCELL_X4 FILLER_115_915 ();
 FILLCELL_X2 FILLER_115_919 ();
 FILLCELL_X1 FILLER_115_921 ();
 FILLCELL_X16 FILLER_115_924 ();
 FILLCELL_X2 FILLER_115_940 ();
 FILLCELL_X16 FILLER_115_944 ();
 FILLCELL_X8 FILLER_115_960 ();
 FILLCELL_X4 FILLER_115_968 ();
 FILLCELL_X2 FILLER_115_972 ();
 FILLCELL_X16 FILLER_115_976 ();
 FILLCELL_X8 FILLER_115_992 ();
 FILLCELL_X2 FILLER_115_1000 ();
 FILLCELL_X1 FILLER_115_1002 ();
 FILLCELL_X32 FILLER_115_1010 ();
 FILLCELL_X4 FILLER_115_1042 ();
 FILLCELL_X2 FILLER_115_1046 ();
 FILLCELL_X1 FILLER_115_1048 ();
 FILLCELL_X8 FILLER_115_1065 ();
 FILLCELL_X4 FILLER_115_1073 ();
 FILLCELL_X8 FILLER_115_1093 ();
 FILLCELL_X1 FILLER_115_1101 ();
 FILLCELL_X32 FILLER_115_1118 ();
 FILLCELL_X32 FILLER_115_1150 ();
 FILLCELL_X32 FILLER_115_1182 ();
 FILLCELL_X32 FILLER_115_1214 ();
 FILLCELL_X16 FILLER_115_1246 ();
 FILLCELL_X1 FILLER_115_1262 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X32 FILLER_115_1552 ();
 FILLCELL_X32 FILLER_115_1584 ();
 FILLCELL_X32 FILLER_115_1616 ();
 FILLCELL_X32 FILLER_115_1648 ();
 FILLCELL_X32 FILLER_115_1680 ();
 FILLCELL_X32 FILLER_115_1712 ();
 FILLCELL_X32 FILLER_115_1744 ();
 FILLCELL_X32 FILLER_115_1776 ();
 FILLCELL_X32 FILLER_115_1808 ();
 FILLCELL_X32 FILLER_115_1840 ();
 FILLCELL_X8 FILLER_115_1872 ();
 FILLCELL_X8 FILLER_115_1883 ();
 FILLCELL_X4 FILLER_115_1891 ();
 FILLCELL_X1 FILLER_115_1895 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X16 FILLER_116_792 ();
 FILLCELL_X4 FILLER_116_808 ();
 FILLCELL_X16 FILLER_116_816 ();
 FILLCELL_X2 FILLER_116_832 ();
 FILLCELL_X1 FILLER_116_834 ();
 FILLCELL_X4 FILLER_116_851 ();
 FILLCELL_X2 FILLER_116_855 ();
 FILLCELL_X1 FILLER_116_857 ();
 FILLCELL_X16 FILLER_116_868 ();
 FILLCELL_X8 FILLER_116_884 ();
 FILLCELL_X4 FILLER_116_894 ();
 FILLCELL_X2 FILLER_116_898 ();
 FILLCELL_X4 FILLER_116_903 ();
 FILLCELL_X2 FILLER_116_907 ();
 FILLCELL_X8 FILLER_116_925 ();
 FILLCELL_X4 FILLER_116_933 ();
 FILLCELL_X2 FILLER_116_937 ();
 FILLCELL_X8 FILLER_116_949 ();
 FILLCELL_X2 FILLER_116_957 ();
 FILLCELL_X1 FILLER_116_959 ();
 FILLCELL_X1 FILLER_116_970 ();
 FILLCELL_X8 FILLER_116_987 ();
 FILLCELL_X4 FILLER_116_995 ();
 FILLCELL_X2 FILLER_116_999 ();
 FILLCELL_X32 FILLER_116_1017 ();
 FILLCELL_X2 FILLER_116_1049 ();
 FILLCELL_X2 FILLER_116_1054 ();
 FILLCELL_X32 FILLER_116_1059 ();
 FILLCELL_X8 FILLER_116_1091 ();
 FILLCELL_X2 FILLER_116_1099 ();
 FILLCELL_X4 FILLER_116_1104 ();
 FILLCELL_X2 FILLER_116_1108 ();
 FILLCELL_X1 FILLER_116_1110 ();
 FILLCELL_X2 FILLER_116_1127 ();
 FILLCELL_X1 FILLER_116_1129 ();
 FILLCELL_X16 FILLER_116_1132 ();
 FILLCELL_X4 FILLER_116_1148 ();
 FILLCELL_X2 FILLER_116_1152 ();
 FILLCELL_X1 FILLER_116_1154 ();
 FILLCELL_X2 FILLER_116_1165 ();
 FILLCELL_X4 FILLER_116_1171 ();
 FILLCELL_X2 FILLER_116_1175 ();
 FILLCELL_X32 FILLER_116_1215 ();
 FILLCELL_X32 FILLER_116_1247 ();
 FILLCELL_X32 FILLER_116_1279 ();
 FILLCELL_X32 FILLER_116_1311 ();
 FILLCELL_X32 FILLER_116_1343 ();
 FILLCELL_X32 FILLER_116_1375 ();
 FILLCELL_X32 FILLER_116_1407 ();
 FILLCELL_X32 FILLER_116_1439 ();
 FILLCELL_X32 FILLER_116_1471 ();
 FILLCELL_X32 FILLER_116_1503 ();
 FILLCELL_X32 FILLER_116_1535 ();
 FILLCELL_X32 FILLER_116_1567 ();
 FILLCELL_X32 FILLER_116_1599 ();
 FILLCELL_X32 FILLER_116_1631 ();
 FILLCELL_X32 FILLER_116_1663 ();
 FILLCELL_X32 FILLER_116_1695 ();
 FILLCELL_X32 FILLER_116_1727 ();
 FILLCELL_X32 FILLER_116_1759 ();
 FILLCELL_X32 FILLER_116_1791 ();
 FILLCELL_X32 FILLER_116_1823 ();
 FILLCELL_X32 FILLER_116_1855 ();
 FILLCELL_X4 FILLER_116_1887 ();
 FILLCELL_X2 FILLER_116_1891 ();
 FILLCELL_X1 FILLER_116_1893 ();
 FILLCELL_X1 FILLER_116_1895 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X8 FILLER_117_801 ();
 FILLCELL_X2 FILLER_117_809 ();
 FILLCELL_X4 FILLER_117_837 ();
 FILLCELL_X2 FILLER_117_841 ();
 FILLCELL_X1 FILLER_117_843 ();
 FILLCELL_X4 FILLER_117_863 ();
 FILLCELL_X1 FILLER_117_867 ();
 FILLCELL_X16 FILLER_117_870 ();
 FILLCELL_X1 FILLER_117_893 ();
 FILLCELL_X16 FILLER_117_914 ();
 FILLCELL_X4 FILLER_117_930 ();
 FILLCELL_X1 FILLER_117_934 ();
 FILLCELL_X8 FILLER_117_939 ();
 FILLCELL_X8 FILLER_117_951 ();
 FILLCELL_X4 FILLER_117_959 ();
 FILLCELL_X2 FILLER_117_963 ();
 FILLCELL_X8 FILLER_117_970 ();
 FILLCELL_X2 FILLER_117_978 ();
 FILLCELL_X16 FILLER_117_987 ();
 FILLCELL_X4 FILLER_117_1003 ();
 FILLCELL_X1 FILLER_117_1007 ();
 FILLCELL_X32 FILLER_117_1011 ();
 FILLCELL_X1 FILLER_117_1043 ();
 FILLCELL_X16 FILLER_117_1060 ();
 FILLCELL_X4 FILLER_117_1076 ();
 FILLCELL_X2 FILLER_117_1080 ();
 FILLCELL_X1 FILLER_117_1082 ();
 FILLCELL_X16 FILLER_117_1087 ();
 FILLCELL_X8 FILLER_117_1103 ();
 FILLCELL_X2 FILLER_117_1111 ();
 FILLCELL_X1 FILLER_117_1113 ();
 FILLCELL_X32 FILLER_117_1116 ();
 FILLCELL_X32 FILLER_117_1148 ();
 FILLCELL_X32 FILLER_117_1180 ();
 FILLCELL_X32 FILLER_117_1212 ();
 FILLCELL_X16 FILLER_117_1244 ();
 FILLCELL_X2 FILLER_117_1260 ();
 FILLCELL_X1 FILLER_117_1262 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X32 FILLER_117_1552 ();
 FILLCELL_X32 FILLER_117_1584 ();
 FILLCELL_X32 FILLER_117_1616 ();
 FILLCELL_X32 FILLER_117_1648 ();
 FILLCELL_X32 FILLER_117_1680 ();
 FILLCELL_X32 FILLER_117_1712 ();
 FILLCELL_X32 FILLER_117_1744 ();
 FILLCELL_X32 FILLER_117_1776 ();
 FILLCELL_X32 FILLER_117_1808 ();
 FILLCELL_X32 FILLER_117_1840 ();
 FILLCELL_X16 FILLER_117_1872 ();
 FILLCELL_X8 FILLER_117_1888 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_741 ();
 FILLCELL_X32 FILLER_118_773 ();
 FILLCELL_X16 FILLER_118_805 ();
 FILLCELL_X4 FILLER_118_821 ();
 FILLCELL_X2 FILLER_118_825 ();
 FILLCELL_X16 FILLER_118_836 ();
 FILLCELL_X16 FILLER_118_856 ();
 FILLCELL_X8 FILLER_118_872 ();
 FILLCELL_X2 FILLER_118_880 ();
 FILLCELL_X16 FILLER_118_898 ();
 FILLCELL_X8 FILLER_118_914 ();
 FILLCELL_X4 FILLER_118_922 ();
 FILLCELL_X2 FILLER_118_926 ();
 FILLCELL_X1 FILLER_118_928 ();
 FILLCELL_X16 FILLER_118_945 ();
 FILLCELL_X8 FILLER_118_961 ();
 FILLCELL_X2 FILLER_118_969 ();
 FILLCELL_X8 FILLER_118_987 ();
 FILLCELL_X4 FILLER_118_995 ();
 FILLCELL_X1 FILLER_118_999 ();
 FILLCELL_X32 FILLER_118_1016 ();
 FILLCELL_X4 FILLER_118_1048 ();
 FILLCELL_X1 FILLER_118_1052 ();
 FILLCELL_X16 FILLER_118_1056 ();
 FILLCELL_X4 FILLER_118_1072 ();
 FILLCELL_X1 FILLER_118_1076 ();
 FILLCELL_X2 FILLER_118_1081 ();
 FILLCELL_X32 FILLER_118_1095 ();
 FILLCELL_X32 FILLER_118_1127 ();
 FILLCELL_X32 FILLER_118_1159 ();
 FILLCELL_X32 FILLER_118_1191 ();
 FILLCELL_X32 FILLER_118_1223 ();
 FILLCELL_X32 FILLER_118_1255 ();
 FILLCELL_X32 FILLER_118_1287 ();
 FILLCELL_X32 FILLER_118_1319 ();
 FILLCELL_X32 FILLER_118_1351 ();
 FILLCELL_X32 FILLER_118_1383 ();
 FILLCELL_X32 FILLER_118_1415 ();
 FILLCELL_X32 FILLER_118_1447 ();
 FILLCELL_X32 FILLER_118_1479 ();
 FILLCELL_X32 FILLER_118_1511 ();
 FILLCELL_X32 FILLER_118_1543 ();
 FILLCELL_X32 FILLER_118_1575 ();
 FILLCELL_X32 FILLER_118_1607 ();
 FILLCELL_X32 FILLER_118_1639 ();
 FILLCELL_X32 FILLER_118_1671 ();
 FILLCELL_X32 FILLER_118_1703 ();
 FILLCELL_X32 FILLER_118_1735 ();
 FILLCELL_X32 FILLER_118_1767 ();
 FILLCELL_X32 FILLER_118_1799 ();
 FILLCELL_X32 FILLER_118_1831 ();
 FILLCELL_X8 FILLER_118_1863 ();
 FILLCELL_X4 FILLER_118_1871 ();
 FILLCELL_X1 FILLER_118_1875 ();
 FILLCELL_X8 FILLER_118_1879 ();
 FILLCELL_X4 FILLER_118_1887 ();
 FILLCELL_X2 FILLER_118_1891 ();
 FILLCELL_X1 FILLER_118_1893 ();
 FILLCELL_X1 FILLER_118_1895 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X8 FILLER_119_801 ();
 FILLCELL_X2 FILLER_119_809 ();
 FILLCELL_X4 FILLER_119_827 ();
 FILLCELL_X2 FILLER_119_831 ();
 FILLCELL_X16 FILLER_119_836 ();
 FILLCELL_X8 FILLER_119_852 ();
 FILLCELL_X4 FILLER_119_860 ();
 FILLCELL_X1 FILLER_119_867 ();
 FILLCELL_X16 FILLER_119_873 ();
 FILLCELL_X8 FILLER_119_889 ();
 FILLCELL_X2 FILLER_119_897 ();
 FILLCELL_X1 FILLER_119_899 ();
 FILLCELL_X32 FILLER_119_905 ();
 FILLCELL_X32 FILLER_119_937 ();
 FILLCELL_X32 FILLER_119_969 ();
 FILLCELL_X2 FILLER_119_1001 ();
 FILLCELL_X1 FILLER_119_1003 ();
 FILLCELL_X2 FILLER_119_1007 ();
 FILLCELL_X4 FILLER_119_1014 ();
 FILLCELL_X2 FILLER_119_1018 ();
 FILLCELL_X16 FILLER_119_1036 ();
 FILLCELL_X8 FILLER_119_1052 ();
 FILLCELL_X4 FILLER_119_1060 ();
 FILLCELL_X8 FILLER_119_1078 ();
 FILLCELL_X2 FILLER_119_1086 ();
 FILLCELL_X1 FILLER_119_1088 ();
 FILLCELL_X4 FILLER_119_1105 ();
 FILLCELL_X4 FILLER_119_1111 ();
 FILLCELL_X2 FILLER_119_1115 ();
 FILLCELL_X32 FILLER_119_1141 ();
 FILLCELL_X32 FILLER_119_1173 ();
 FILLCELL_X32 FILLER_119_1205 ();
 FILLCELL_X16 FILLER_119_1237 ();
 FILLCELL_X8 FILLER_119_1253 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X32 FILLER_119_1552 ();
 FILLCELL_X32 FILLER_119_1584 ();
 FILLCELL_X32 FILLER_119_1616 ();
 FILLCELL_X32 FILLER_119_1648 ();
 FILLCELL_X32 FILLER_119_1680 ();
 FILLCELL_X32 FILLER_119_1712 ();
 FILLCELL_X32 FILLER_119_1744 ();
 FILLCELL_X32 FILLER_119_1776 ();
 FILLCELL_X32 FILLER_119_1808 ();
 FILLCELL_X32 FILLER_119_1840 ();
 FILLCELL_X16 FILLER_119_1872 ();
 FILLCELL_X8 FILLER_119_1888 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X8 FILLER_120_760 ();
 FILLCELL_X4 FILLER_120_768 ();
 FILLCELL_X2 FILLER_120_772 ();
 FILLCELL_X16 FILLER_120_778 ();
 FILLCELL_X8 FILLER_120_794 ();
 FILLCELL_X4 FILLER_120_802 ();
 FILLCELL_X8 FILLER_120_810 ();
 FILLCELL_X1 FILLER_120_818 ();
 FILLCELL_X2 FILLER_120_826 ();
 FILLCELL_X1 FILLER_120_828 ();
 FILLCELL_X4 FILLER_120_845 ();
 FILLCELL_X4 FILLER_120_865 ();
 FILLCELL_X16 FILLER_120_879 ();
 FILLCELL_X1 FILLER_120_895 ();
 FILLCELL_X16 FILLER_120_909 ();
 FILLCELL_X8 FILLER_120_927 ();
 FILLCELL_X1 FILLER_120_935 ();
 FILLCELL_X1 FILLER_120_942 ();
 FILLCELL_X4 FILLER_120_945 ();
 FILLCELL_X16 FILLER_120_965 ();
 FILLCELL_X16 FILLER_120_984 ();
 FILLCELL_X1 FILLER_120_1000 ();
 FILLCELL_X32 FILLER_120_1017 ();
 FILLCELL_X1 FILLER_120_1049 ();
 FILLCELL_X32 FILLER_120_1093 ();
 FILLCELL_X32 FILLER_120_1125 ();
 FILLCELL_X32 FILLER_120_1157 ();
 FILLCELL_X32 FILLER_120_1189 ();
 FILLCELL_X32 FILLER_120_1221 ();
 FILLCELL_X32 FILLER_120_1253 ();
 FILLCELL_X32 FILLER_120_1285 ();
 FILLCELL_X32 FILLER_120_1317 ();
 FILLCELL_X32 FILLER_120_1349 ();
 FILLCELL_X32 FILLER_120_1381 ();
 FILLCELL_X32 FILLER_120_1413 ();
 FILLCELL_X32 FILLER_120_1445 ();
 FILLCELL_X32 FILLER_120_1477 ();
 FILLCELL_X32 FILLER_120_1509 ();
 FILLCELL_X32 FILLER_120_1541 ();
 FILLCELL_X32 FILLER_120_1573 ();
 FILLCELL_X32 FILLER_120_1605 ();
 FILLCELL_X32 FILLER_120_1637 ();
 FILLCELL_X32 FILLER_120_1669 ();
 FILLCELL_X32 FILLER_120_1701 ();
 FILLCELL_X32 FILLER_120_1733 ();
 FILLCELL_X32 FILLER_120_1765 ();
 FILLCELL_X32 FILLER_120_1797 ();
 FILLCELL_X32 FILLER_120_1829 ();
 FILLCELL_X32 FILLER_120_1861 ();
 FILLCELL_X1 FILLER_120_1893 ();
 FILLCELL_X1 FILLER_120_1895 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X16 FILLER_121_769 ();
 FILLCELL_X8 FILLER_121_785 ();
 FILLCELL_X4 FILLER_121_793 ();
 FILLCELL_X1 FILLER_121_801 ();
 FILLCELL_X8 FILLER_121_812 ();
 FILLCELL_X1 FILLER_121_820 ();
 FILLCELL_X8 FILLER_121_831 ();
 FILLCELL_X4 FILLER_121_839 ();
 FILLCELL_X1 FILLER_121_843 ();
 FILLCELL_X8 FILLER_121_860 ();
 FILLCELL_X4 FILLER_121_868 ();
 FILLCELL_X2 FILLER_121_872 ();
 FILLCELL_X1 FILLER_121_874 ();
 FILLCELL_X16 FILLER_121_891 ();
 FILLCELL_X8 FILLER_121_907 ();
 FILLCELL_X2 FILLER_121_915 ();
 FILLCELL_X16 FILLER_121_949 ();
 FILLCELL_X8 FILLER_121_965 ();
 FILLCELL_X1 FILLER_121_973 ();
 FILLCELL_X16 FILLER_121_990 ();
 FILLCELL_X2 FILLER_121_1006 ();
 FILLCELL_X1 FILLER_121_1008 ();
 FILLCELL_X32 FILLER_121_1025 ();
 FILLCELL_X2 FILLER_121_1057 ();
 FILLCELL_X1 FILLER_121_1059 ();
 FILLCELL_X32 FILLER_121_1062 ();
 FILLCELL_X32 FILLER_121_1097 ();
 FILLCELL_X32 FILLER_121_1129 ();
 FILLCELL_X32 FILLER_121_1161 ();
 FILLCELL_X32 FILLER_121_1193 ();
 FILLCELL_X32 FILLER_121_1225 ();
 FILLCELL_X4 FILLER_121_1257 ();
 FILLCELL_X2 FILLER_121_1261 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X32 FILLER_121_1552 ();
 FILLCELL_X32 FILLER_121_1584 ();
 FILLCELL_X32 FILLER_121_1616 ();
 FILLCELL_X32 FILLER_121_1648 ();
 FILLCELL_X32 FILLER_121_1680 ();
 FILLCELL_X32 FILLER_121_1712 ();
 FILLCELL_X32 FILLER_121_1744 ();
 FILLCELL_X32 FILLER_121_1776 ();
 FILLCELL_X32 FILLER_121_1808 ();
 FILLCELL_X32 FILLER_121_1840 ();
 FILLCELL_X16 FILLER_121_1872 ();
 FILLCELL_X8 FILLER_121_1888 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X8 FILLER_122_792 ();
 FILLCELL_X2 FILLER_122_800 ();
 FILLCELL_X1 FILLER_122_802 ();
 FILLCELL_X32 FILLER_122_809 ();
 FILLCELL_X16 FILLER_122_841 ();
 FILLCELL_X8 FILLER_122_857 ();
 FILLCELL_X16 FILLER_122_867 ();
 FILLCELL_X4 FILLER_122_883 ();
 FILLCELL_X2 FILLER_122_887 ();
 FILLCELL_X4 FILLER_122_895 ();
 FILLCELL_X16 FILLER_122_915 ();
 FILLCELL_X4 FILLER_122_931 ();
 FILLCELL_X1 FILLER_122_935 ();
 FILLCELL_X16 FILLER_122_941 ();
 FILLCELL_X2 FILLER_122_957 ();
 FILLCELL_X1 FILLER_122_959 ();
 FILLCELL_X2 FILLER_122_976 ();
 FILLCELL_X4 FILLER_122_981 ();
 FILLCELL_X2 FILLER_122_985 ();
 FILLCELL_X1 FILLER_122_987 ();
 FILLCELL_X32 FILLER_122_1004 ();
 FILLCELL_X32 FILLER_122_1036 ();
 FILLCELL_X16 FILLER_122_1068 ();
 FILLCELL_X8 FILLER_122_1084 ();
 FILLCELL_X32 FILLER_122_1108 ();
 FILLCELL_X32 FILLER_122_1140 ();
 FILLCELL_X32 FILLER_122_1172 ();
 FILLCELL_X32 FILLER_122_1204 ();
 FILLCELL_X32 FILLER_122_1236 ();
 FILLCELL_X32 FILLER_122_1268 ();
 FILLCELL_X32 FILLER_122_1300 ();
 FILLCELL_X32 FILLER_122_1332 ();
 FILLCELL_X32 FILLER_122_1364 ();
 FILLCELL_X32 FILLER_122_1396 ();
 FILLCELL_X32 FILLER_122_1428 ();
 FILLCELL_X32 FILLER_122_1460 ();
 FILLCELL_X32 FILLER_122_1492 ();
 FILLCELL_X32 FILLER_122_1524 ();
 FILLCELL_X32 FILLER_122_1556 ();
 FILLCELL_X32 FILLER_122_1588 ();
 FILLCELL_X32 FILLER_122_1620 ();
 FILLCELL_X32 FILLER_122_1652 ();
 FILLCELL_X32 FILLER_122_1684 ();
 FILLCELL_X32 FILLER_122_1716 ();
 FILLCELL_X32 FILLER_122_1748 ();
 FILLCELL_X32 FILLER_122_1780 ();
 FILLCELL_X32 FILLER_122_1812 ();
 FILLCELL_X32 FILLER_122_1844 ();
 FILLCELL_X16 FILLER_122_1876 ();
 FILLCELL_X2 FILLER_122_1892 ();
 FILLCELL_X1 FILLER_122_1895 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X4 FILLER_123_769 ();
 FILLCELL_X2 FILLER_123_773 ();
 FILLCELL_X4 FILLER_123_809 ();
 FILLCELL_X2 FILLER_123_813 ();
 FILLCELL_X8 FILLER_123_831 ();
 FILLCELL_X4 FILLER_123_839 ();
 FILLCELL_X32 FILLER_123_846 ();
 FILLCELL_X8 FILLER_123_878 ();
 FILLCELL_X2 FILLER_123_886 ();
 FILLCELL_X1 FILLER_123_888 ();
 FILLCELL_X4 FILLER_123_893 ();
 FILLCELL_X2 FILLER_123_897 ();
 FILLCELL_X16 FILLER_123_917 ();
 FILLCELL_X4 FILLER_123_933 ();
 FILLCELL_X2 FILLER_123_937 ();
 FILLCELL_X1 FILLER_123_939 ();
 FILLCELL_X16 FILLER_123_950 ();
 FILLCELL_X8 FILLER_123_966 ();
 FILLCELL_X4 FILLER_123_974 ();
 FILLCELL_X1 FILLER_123_978 ();
 FILLCELL_X1 FILLER_123_981 ();
 FILLCELL_X16 FILLER_123_985 ();
 FILLCELL_X4 FILLER_123_1001 ();
 FILLCELL_X2 FILLER_123_1005 ();
 FILLCELL_X16 FILLER_123_1011 ();
 FILLCELL_X4 FILLER_123_1027 ();
 FILLCELL_X1 FILLER_123_1031 ();
 FILLCELL_X16 FILLER_123_1038 ();
 FILLCELL_X1 FILLER_123_1058 ();
 FILLCELL_X32 FILLER_123_1069 ();
 FILLCELL_X8 FILLER_123_1101 ();
 FILLCELL_X4 FILLER_123_1109 ();
 FILLCELL_X2 FILLER_123_1113 ();
 FILLCELL_X32 FILLER_123_1135 ();
 FILLCELL_X32 FILLER_123_1167 ();
 FILLCELL_X32 FILLER_123_1199 ();
 FILLCELL_X32 FILLER_123_1231 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X32 FILLER_123_1552 ();
 FILLCELL_X32 FILLER_123_1584 ();
 FILLCELL_X32 FILLER_123_1616 ();
 FILLCELL_X32 FILLER_123_1648 ();
 FILLCELL_X32 FILLER_123_1680 ();
 FILLCELL_X32 FILLER_123_1712 ();
 FILLCELL_X32 FILLER_123_1744 ();
 FILLCELL_X32 FILLER_123_1776 ();
 FILLCELL_X32 FILLER_123_1808 ();
 FILLCELL_X32 FILLER_123_1840 ();
 FILLCELL_X16 FILLER_123_1872 ();
 FILLCELL_X8 FILLER_123_1888 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X4 FILLER_124_760 ();
 FILLCELL_X2 FILLER_124_764 ();
 FILLCELL_X1 FILLER_124_766 ();
 FILLCELL_X4 FILLER_124_773 ();
 FILLCELL_X4 FILLER_124_793 ();
 FILLCELL_X16 FILLER_124_799 ();
 FILLCELL_X16 FILLER_124_817 ();
 FILLCELL_X4 FILLER_124_833 ();
 FILLCELL_X4 FILLER_124_853 ();
 FILLCELL_X1 FILLER_124_857 ();
 FILLCELL_X4 FILLER_124_874 ();
 FILLCELL_X1 FILLER_124_878 ();
 FILLCELL_X16 FILLER_124_895 ();
 FILLCELL_X2 FILLER_124_911 ();
 FILLCELL_X1 FILLER_124_913 ();
 FILLCELL_X4 FILLER_124_916 ();
 FILLCELL_X1 FILLER_124_920 ();
 FILLCELL_X8 FILLER_124_923 ();
 FILLCELL_X4 FILLER_124_931 ();
 FILLCELL_X1 FILLER_124_935 ();
 FILLCELL_X16 FILLER_124_952 ();
 FILLCELL_X8 FILLER_124_968 ();
 FILLCELL_X2 FILLER_124_976 ();
 FILLCELL_X8 FILLER_124_988 ();
 FILLCELL_X4 FILLER_124_996 ();
 FILLCELL_X2 FILLER_124_1000 ();
 FILLCELL_X8 FILLER_124_1018 ();
 FILLCELL_X1 FILLER_124_1026 ();
 FILLCELL_X2 FILLER_124_1059 ();
 FILLCELL_X1 FILLER_124_1061 ();
 FILLCELL_X32 FILLER_124_1064 ();
 FILLCELL_X32 FILLER_124_1096 ();
 FILLCELL_X1 FILLER_124_1128 ();
 FILLCELL_X32 FILLER_124_1133 ();
 FILLCELL_X32 FILLER_124_1165 ();
 FILLCELL_X32 FILLER_124_1197 ();
 FILLCELL_X32 FILLER_124_1229 ();
 FILLCELL_X32 FILLER_124_1261 ();
 FILLCELL_X32 FILLER_124_1293 ();
 FILLCELL_X32 FILLER_124_1325 ();
 FILLCELL_X32 FILLER_124_1357 ();
 FILLCELL_X32 FILLER_124_1389 ();
 FILLCELL_X32 FILLER_124_1421 ();
 FILLCELL_X32 FILLER_124_1453 ();
 FILLCELL_X32 FILLER_124_1485 ();
 FILLCELL_X32 FILLER_124_1517 ();
 FILLCELL_X32 FILLER_124_1549 ();
 FILLCELL_X32 FILLER_124_1581 ();
 FILLCELL_X32 FILLER_124_1613 ();
 FILLCELL_X32 FILLER_124_1645 ();
 FILLCELL_X32 FILLER_124_1677 ();
 FILLCELL_X32 FILLER_124_1709 ();
 FILLCELL_X32 FILLER_124_1741 ();
 FILLCELL_X32 FILLER_124_1773 ();
 FILLCELL_X32 FILLER_124_1805 ();
 FILLCELL_X32 FILLER_124_1837 ();
 FILLCELL_X16 FILLER_124_1869 ();
 FILLCELL_X8 FILLER_124_1885 ();
 FILLCELL_X1 FILLER_124_1893 ();
 FILLCELL_X1 FILLER_124_1895 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X16 FILLER_125_769 ();
 FILLCELL_X4 FILLER_125_785 ();
 FILLCELL_X2 FILLER_125_789 ();
 FILLCELL_X1 FILLER_125_791 ();
 FILLCELL_X16 FILLER_125_808 ();
 FILLCELL_X4 FILLER_125_824 ();
 FILLCELL_X2 FILLER_125_828 ();
 FILLCELL_X1 FILLER_125_830 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X16 FILLER_125_865 ();
 FILLCELL_X8 FILLER_125_881 ();
 FILLCELL_X4 FILLER_125_889 ();
 FILLCELL_X2 FILLER_125_893 ();
 FILLCELL_X1 FILLER_125_895 ();
 FILLCELL_X8 FILLER_125_898 ();
 FILLCELL_X2 FILLER_125_906 ();
 FILLCELL_X1 FILLER_125_908 ();
 FILLCELL_X32 FILLER_125_925 ();
 FILLCELL_X4 FILLER_125_957 ();
 FILLCELL_X32 FILLER_125_965 ();
 FILLCELL_X16 FILLER_125_997 ();
 FILLCELL_X2 FILLER_125_1013 ();
 FILLCELL_X1 FILLER_125_1015 ();
 FILLCELL_X32 FILLER_125_1032 ();
 FILLCELL_X32 FILLER_125_1080 ();
 FILLCELL_X32 FILLER_125_1112 ();
 FILLCELL_X32 FILLER_125_1144 ();
 FILLCELL_X32 FILLER_125_1176 ();
 FILLCELL_X32 FILLER_125_1208 ();
 FILLCELL_X16 FILLER_125_1240 ();
 FILLCELL_X4 FILLER_125_1256 ();
 FILLCELL_X2 FILLER_125_1260 ();
 FILLCELL_X1 FILLER_125_1262 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X32 FILLER_125_1648 ();
 FILLCELL_X32 FILLER_125_1680 ();
 FILLCELL_X32 FILLER_125_1712 ();
 FILLCELL_X32 FILLER_125_1744 ();
 FILLCELL_X32 FILLER_125_1776 ();
 FILLCELL_X32 FILLER_125_1808 ();
 FILLCELL_X16 FILLER_125_1840 ();
 FILLCELL_X1 FILLER_125_1856 ();
 FILLCELL_X32 FILLER_125_1860 ();
 FILLCELL_X4 FILLER_125_1892 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X16 FILLER_126_760 ();
 FILLCELL_X8 FILLER_126_776 ();
 FILLCELL_X2 FILLER_126_796 ();
 FILLCELL_X8 FILLER_126_801 ();
 FILLCELL_X1 FILLER_126_809 ();
 FILLCELL_X2 FILLER_126_826 ();
 FILLCELL_X1 FILLER_126_828 ();
 FILLCELL_X4 FILLER_126_845 ();
 FILLCELL_X2 FILLER_126_849 ();
 FILLCELL_X1 FILLER_126_851 ();
 FILLCELL_X1 FILLER_126_856 ();
 FILLCELL_X16 FILLER_126_859 ();
 FILLCELL_X8 FILLER_126_875 ();
 FILLCELL_X4 FILLER_126_883 ();
 FILLCELL_X1 FILLER_126_887 ();
 FILLCELL_X16 FILLER_126_904 ();
 FILLCELL_X8 FILLER_126_920 ();
 FILLCELL_X2 FILLER_126_928 ();
 FILLCELL_X1 FILLER_126_930 ();
 FILLCELL_X16 FILLER_126_933 ();
 FILLCELL_X2 FILLER_126_949 ();
 FILLCELL_X1 FILLER_126_951 ();
 FILLCELL_X2 FILLER_126_954 ();
 FILLCELL_X8 FILLER_126_972 ();
 FILLCELL_X4 FILLER_126_980 ();
 FILLCELL_X1 FILLER_126_984 ();
 FILLCELL_X2 FILLER_126_987 ();
 FILLCELL_X1 FILLER_126_989 ();
 FILLCELL_X32 FILLER_126_993 ();
 FILLCELL_X32 FILLER_126_1025 ();
 FILLCELL_X4 FILLER_126_1057 ();
 FILLCELL_X2 FILLER_126_1061 ();
 FILLCELL_X8 FILLER_126_1065 ();
 FILLCELL_X4 FILLER_126_1073 ();
 FILLCELL_X2 FILLER_126_1077 ();
 FILLCELL_X32 FILLER_126_1081 ();
 FILLCELL_X32 FILLER_126_1113 ();
 FILLCELL_X32 FILLER_126_1145 ();
 FILLCELL_X32 FILLER_126_1177 ();
 FILLCELL_X32 FILLER_126_1209 ();
 FILLCELL_X32 FILLER_126_1241 ();
 FILLCELL_X32 FILLER_126_1273 ();
 FILLCELL_X32 FILLER_126_1305 ();
 FILLCELL_X32 FILLER_126_1337 ();
 FILLCELL_X32 FILLER_126_1369 ();
 FILLCELL_X32 FILLER_126_1401 ();
 FILLCELL_X32 FILLER_126_1433 ();
 FILLCELL_X32 FILLER_126_1465 ();
 FILLCELL_X32 FILLER_126_1497 ();
 FILLCELL_X32 FILLER_126_1529 ();
 FILLCELL_X32 FILLER_126_1561 ();
 FILLCELL_X32 FILLER_126_1593 ();
 FILLCELL_X32 FILLER_126_1625 ();
 FILLCELL_X32 FILLER_126_1657 ();
 FILLCELL_X32 FILLER_126_1689 ();
 FILLCELL_X32 FILLER_126_1721 ();
 FILLCELL_X32 FILLER_126_1753 ();
 FILLCELL_X32 FILLER_126_1785 ();
 FILLCELL_X32 FILLER_126_1817 ();
 FILLCELL_X32 FILLER_126_1849 ();
 FILLCELL_X8 FILLER_126_1881 ();
 FILLCELL_X4 FILLER_126_1889 ();
 FILLCELL_X1 FILLER_126_1893 ();
 FILLCELL_X1 FILLER_126_1895 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_803 ();
 FILLCELL_X8 FILLER_127_835 ();
 FILLCELL_X4 FILLER_127_843 ();
 FILLCELL_X8 FILLER_127_865 ();
 FILLCELL_X1 FILLER_127_873 ();
 FILLCELL_X16 FILLER_127_876 ();
 FILLCELL_X8 FILLER_127_892 ();
 FILLCELL_X4 FILLER_127_900 ();
 FILLCELL_X2 FILLER_127_904 ();
 FILLCELL_X4 FILLER_127_908 ();
 FILLCELL_X2 FILLER_127_912 ();
 FILLCELL_X1 FILLER_127_914 ();
 FILLCELL_X4 FILLER_127_917 ();
 FILLCELL_X2 FILLER_127_921 ();
 FILLCELL_X1 FILLER_127_923 ();
 FILLCELL_X32 FILLER_127_940 ();
 FILLCELL_X4 FILLER_127_972 ();
 FILLCELL_X2 FILLER_127_976 ();
 FILLCELL_X1 FILLER_127_978 ();
 FILLCELL_X16 FILLER_127_995 ();
 FILLCELL_X4 FILLER_127_1011 ();
 FILLCELL_X2 FILLER_127_1015 ();
 FILLCELL_X1 FILLER_127_1017 ();
 FILLCELL_X8 FILLER_127_1021 ();
 FILLCELL_X2 FILLER_127_1029 ();
 FILLCELL_X1 FILLER_127_1031 ();
 FILLCELL_X16 FILLER_127_1034 ();
 FILLCELL_X4 FILLER_127_1050 ();
 FILLCELL_X2 FILLER_127_1057 ();
 FILLCELL_X1 FILLER_127_1059 ();
 FILLCELL_X32 FILLER_127_1062 ();
 FILLCELL_X32 FILLER_127_1094 ();
 FILLCELL_X32 FILLER_127_1126 ();
 FILLCELL_X32 FILLER_127_1158 ();
 FILLCELL_X32 FILLER_127_1190 ();
 FILLCELL_X32 FILLER_127_1222 ();
 FILLCELL_X8 FILLER_127_1254 ();
 FILLCELL_X1 FILLER_127_1262 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X32 FILLER_127_1584 ();
 FILLCELL_X32 FILLER_127_1616 ();
 FILLCELL_X32 FILLER_127_1648 ();
 FILLCELL_X32 FILLER_127_1680 ();
 FILLCELL_X32 FILLER_127_1712 ();
 FILLCELL_X32 FILLER_127_1744 ();
 FILLCELL_X32 FILLER_127_1776 ();
 FILLCELL_X32 FILLER_127_1808 ();
 FILLCELL_X32 FILLER_127_1840 ();
 FILLCELL_X16 FILLER_127_1872 ();
 FILLCELL_X8 FILLER_127_1888 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X4 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_798 ();
 FILLCELL_X8 FILLER_128_830 ();
 FILLCELL_X1 FILLER_128_838 ();
 FILLCELL_X8 FILLER_128_855 ();
 FILLCELL_X2 FILLER_128_863 ();
 FILLCELL_X1 FILLER_128_865 ();
 FILLCELL_X1 FILLER_128_882 ();
 FILLCELL_X16 FILLER_128_885 ();
 FILLCELL_X2 FILLER_128_901 ();
 FILLCELL_X16 FILLER_128_905 ();
 FILLCELL_X8 FILLER_128_921 ();
 FILLCELL_X2 FILLER_128_929 ();
 FILLCELL_X8 FILLER_128_933 ();
 FILLCELL_X2 FILLER_128_941 ();
 FILLCELL_X1 FILLER_128_943 ();
 FILLCELL_X4 FILLER_128_946 ();
 FILLCELL_X2 FILLER_128_950 ();
 FILLCELL_X1 FILLER_128_952 ();
 FILLCELL_X16 FILLER_128_955 ();
 FILLCELL_X1 FILLER_128_971 ();
 FILLCELL_X8 FILLER_128_1004 ();
 FILLCELL_X4 FILLER_128_1012 ();
 FILLCELL_X16 FILLER_128_1045 ();
 FILLCELL_X1 FILLER_128_1061 ();
 FILLCELL_X8 FILLER_128_1078 ();
 FILLCELL_X32 FILLER_128_1096 ();
 FILLCELL_X32 FILLER_128_1128 ();
 FILLCELL_X32 FILLER_128_1160 ();
 FILLCELL_X32 FILLER_128_1192 ();
 FILLCELL_X32 FILLER_128_1224 ();
 FILLCELL_X32 FILLER_128_1256 ();
 FILLCELL_X32 FILLER_128_1288 ();
 FILLCELL_X32 FILLER_128_1320 ();
 FILLCELL_X32 FILLER_128_1352 ();
 FILLCELL_X32 FILLER_128_1384 ();
 FILLCELL_X32 FILLER_128_1416 ();
 FILLCELL_X32 FILLER_128_1448 ();
 FILLCELL_X32 FILLER_128_1480 ();
 FILLCELL_X32 FILLER_128_1512 ();
 FILLCELL_X32 FILLER_128_1544 ();
 FILLCELL_X32 FILLER_128_1576 ();
 FILLCELL_X32 FILLER_128_1608 ();
 FILLCELL_X32 FILLER_128_1640 ();
 FILLCELL_X32 FILLER_128_1672 ();
 FILLCELL_X32 FILLER_128_1704 ();
 FILLCELL_X32 FILLER_128_1736 ();
 FILLCELL_X32 FILLER_128_1768 ();
 FILLCELL_X32 FILLER_128_1800 ();
 FILLCELL_X32 FILLER_128_1832 ();
 FILLCELL_X16 FILLER_128_1864 ();
 FILLCELL_X8 FILLER_128_1880 ();
 FILLCELL_X4 FILLER_128_1888 ();
 FILLCELL_X2 FILLER_128_1892 ();
 FILLCELL_X1 FILLER_128_1895 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X16 FILLER_129_769 ();
 FILLCELL_X4 FILLER_129_785 ();
 FILLCELL_X8 FILLER_129_805 ();
 FILLCELL_X4 FILLER_129_813 ();
 FILLCELL_X2 FILLER_129_817 ();
 FILLCELL_X1 FILLER_129_819 ();
 FILLCELL_X32 FILLER_129_830 ();
 FILLCELL_X16 FILLER_129_862 ();
 FILLCELL_X4 FILLER_129_878 ();
 FILLCELL_X1 FILLER_129_882 ();
 FILLCELL_X8 FILLER_129_893 ();
 FILLCELL_X4 FILLER_129_901 ();
 FILLCELL_X2 FILLER_129_905 ();
 FILLCELL_X8 FILLER_129_919 ();
 FILLCELL_X4 FILLER_129_927 ();
 FILLCELL_X2 FILLER_129_931 ();
 FILLCELL_X4 FILLER_129_943 ();
 FILLCELL_X32 FILLER_129_949 ();
 FILLCELL_X16 FILLER_129_981 ();
 FILLCELL_X8 FILLER_129_997 ();
 FILLCELL_X2 FILLER_129_1023 ();
 FILLCELL_X1 FILLER_129_1025 ();
 FILLCELL_X8 FILLER_129_1028 ();
 FILLCELL_X4 FILLER_129_1036 ();
 FILLCELL_X2 FILLER_129_1040 ();
 FILLCELL_X32 FILLER_129_1058 ();
 FILLCELL_X8 FILLER_129_1090 ();
 FILLCELL_X32 FILLER_129_1108 ();
 FILLCELL_X32 FILLER_129_1140 ();
 FILLCELL_X32 FILLER_129_1172 ();
 FILLCELL_X32 FILLER_129_1204 ();
 FILLCELL_X16 FILLER_129_1236 ();
 FILLCELL_X8 FILLER_129_1252 ();
 FILLCELL_X2 FILLER_129_1260 ();
 FILLCELL_X1 FILLER_129_1262 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X32 FILLER_129_1584 ();
 FILLCELL_X32 FILLER_129_1616 ();
 FILLCELL_X32 FILLER_129_1648 ();
 FILLCELL_X32 FILLER_129_1680 ();
 FILLCELL_X32 FILLER_129_1712 ();
 FILLCELL_X32 FILLER_129_1744 ();
 FILLCELL_X32 FILLER_129_1776 ();
 FILLCELL_X32 FILLER_129_1808 ();
 FILLCELL_X32 FILLER_129_1840 ();
 FILLCELL_X16 FILLER_129_1872 ();
 FILLCELL_X8 FILLER_129_1888 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X16 FILLER_130_760 ();
 FILLCELL_X8 FILLER_130_776 ();
 FILLCELL_X4 FILLER_130_784 ();
 FILLCELL_X1 FILLER_130_788 ();
 FILLCELL_X8 FILLER_130_795 ();
 FILLCELL_X16 FILLER_130_813 ();
 FILLCELL_X4 FILLER_130_829 ();
 FILLCELL_X2 FILLER_130_833 ();
 FILLCELL_X1 FILLER_130_835 ();
 FILLCELL_X4 FILLER_130_838 ();
 FILLCELL_X1 FILLER_130_842 ();
 FILLCELL_X8 FILLER_130_845 ();
 FILLCELL_X1 FILLER_130_853 ();
 FILLCELL_X16 FILLER_130_856 ();
 FILLCELL_X8 FILLER_130_872 ();
 FILLCELL_X16 FILLER_130_883 ();
 FILLCELL_X8 FILLER_130_899 ();
 FILLCELL_X2 FILLER_130_907 ();
 FILLCELL_X1 FILLER_130_909 ();
 FILLCELL_X16 FILLER_130_913 ();
 FILLCELL_X8 FILLER_130_929 ();
 FILLCELL_X4 FILLER_130_937 ();
 FILLCELL_X2 FILLER_130_941 ();
 FILLCELL_X1 FILLER_130_943 ();
 FILLCELL_X32 FILLER_130_954 ();
 FILLCELL_X8 FILLER_130_986 ();
 FILLCELL_X4 FILLER_130_994 ();
 FILLCELL_X2 FILLER_130_998 ();
 FILLCELL_X16 FILLER_130_1005 ();
 FILLCELL_X4 FILLER_130_1021 ();
 FILLCELL_X1 FILLER_130_1025 ();
 FILLCELL_X16 FILLER_130_1029 ();
 FILLCELL_X8 FILLER_130_1045 ();
 FILLCELL_X4 FILLER_130_1053 ();
 FILLCELL_X1 FILLER_130_1057 ();
 FILLCELL_X16 FILLER_130_1068 ();
 FILLCELL_X8 FILLER_130_1084 ();
 FILLCELL_X2 FILLER_130_1092 ();
 FILLCELL_X4 FILLER_130_1107 ();
 FILLCELL_X2 FILLER_130_1113 ();
 FILLCELL_X1 FILLER_130_1115 ();
 FILLCELL_X32 FILLER_130_1124 ();
 FILLCELL_X32 FILLER_130_1156 ();
 FILLCELL_X32 FILLER_130_1188 ();
 FILLCELL_X32 FILLER_130_1220 ();
 FILLCELL_X32 FILLER_130_1252 ();
 FILLCELL_X32 FILLER_130_1284 ();
 FILLCELL_X32 FILLER_130_1316 ();
 FILLCELL_X32 FILLER_130_1348 ();
 FILLCELL_X32 FILLER_130_1380 ();
 FILLCELL_X32 FILLER_130_1412 ();
 FILLCELL_X32 FILLER_130_1444 ();
 FILLCELL_X32 FILLER_130_1476 ();
 FILLCELL_X32 FILLER_130_1508 ();
 FILLCELL_X32 FILLER_130_1540 ();
 FILLCELL_X32 FILLER_130_1572 ();
 FILLCELL_X32 FILLER_130_1604 ();
 FILLCELL_X32 FILLER_130_1636 ();
 FILLCELL_X32 FILLER_130_1668 ();
 FILLCELL_X32 FILLER_130_1700 ();
 FILLCELL_X32 FILLER_130_1732 ();
 FILLCELL_X32 FILLER_130_1764 ();
 FILLCELL_X32 FILLER_130_1796 ();
 FILLCELL_X32 FILLER_130_1828 ();
 FILLCELL_X32 FILLER_130_1860 ();
 FILLCELL_X2 FILLER_130_1892 ();
 FILLCELL_X1 FILLER_130_1895 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X8 FILLER_131_801 ();
 FILLCELL_X2 FILLER_131_809 ();
 FILLCELL_X16 FILLER_131_824 ();
 FILLCELL_X2 FILLER_131_840 ();
 FILLCELL_X1 FILLER_131_842 ();
 FILLCELL_X8 FILLER_131_853 ();
 FILLCELL_X2 FILLER_131_861 ();
 FILLCELL_X1 FILLER_131_863 ();
 FILLCELL_X8 FILLER_131_866 ();
 FILLCELL_X4 FILLER_131_874 ();
 FILLCELL_X1 FILLER_131_878 ();
 FILLCELL_X4 FILLER_131_881 ();
 FILLCELL_X2 FILLER_131_885 ();
 FILLCELL_X1 FILLER_131_887 ();
 FILLCELL_X16 FILLER_131_891 ();
 FILLCELL_X8 FILLER_131_907 ();
 FILLCELL_X2 FILLER_131_915 ();
 FILLCELL_X1 FILLER_131_923 ();
 FILLCELL_X32 FILLER_131_928 ();
 FILLCELL_X16 FILLER_131_960 ();
 FILLCELL_X8 FILLER_131_976 ();
 FILLCELL_X2 FILLER_131_984 ();
 FILLCELL_X4 FILLER_131_989 ();
 FILLCELL_X2 FILLER_131_993 ();
 FILLCELL_X32 FILLER_131_998 ();
 FILLCELL_X16 FILLER_131_1030 ();
 FILLCELL_X8 FILLER_131_1046 ();
 FILLCELL_X4 FILLER_131_1054 ();
 FILLCELL_X8 FILLER_131_1064 ();
 FILLCELL_X2 FILLER_131_1072 ();
 FILLCELL_X1 FILLER_131_1074 ();
 FILLCELL_X16 FILLER_131_1085 ();
 FILLCELL_X8 FILLER_131_1101 ();
 FILLCELL_X32 FILLER_131_1125 ();
 FILLCELL_X32 FILLER_131_1157 ();
 FILLCELL_X32 FILLER_131_1189 ();
 FILLCELL_X32 FILLER_131_1221 ();
 FILLCELL_X8 FILLER_131_1253 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X32 FILLER_131_1584 ();
 FILLCELL_X32 FILLER_131_1616 ();
 FILLCELL_X32 FILLER_131_1648 ();
 FILLCELL_X32 FILLER_131_1680 ();
 FILLCELL_X32 FILLER_131_1712 ();
 FILLCELL_X32 FILLER_131_1744 ();
 FILLCELL_X32 FILLER_131_1776 ();
 FILLCELL_X32 FILLER_131_1808 ();
 FILLCELL_X32 FILLER_131_1840 ();
 FILLCELL_X16 FILLER_131_1872 ();
 FILLCELL_X8 FILLER_131_1888 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X16 FILLER_132_792 ();
 FILLCELL_X8 FILLER_132_808 ();
 FILLCELL_X4 FILLER_132_816 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X8 FILLER_132_866 ();
 FILLCELL_X4 FILLER_132_874 ();
 FILLCELL_X2 FILLER_132_878 ();
 FILLCELL_X8 FILLER_132_903 ();
 FILLCELL_X2 FILLER_132_911 ();
 FILLCELL_X1 FILLER_132_913 ();
 FILLCELL_X1 FILLER_132_921 ();
 FILLCELL_X4 FILLER_132_926 ();
 FILLCELL_X1 FILLER_132_930 ();
 FILLCELL_X2 FILLER_132_934 ();
 FILLCELL_X1 FILLER_132_936 ();
 FILLCELL_X32 FILLER_132_939 ();
 FILLCELL_X8 FILLER_132_971 ();
 FILLCELL_X4 FILLER_132_979 ();
 FILLCELL_X2 FILLER_132_983 ();
 FILLCELL_X2 FILLER_132_995 ();
 FILLCELL_X1 FILLER_132_997 ();
 FILLCELL_X16 FILLER_132_1008 ();
 FILLCELL_X1 FILLER_132_1024 ();
 FILLCELL_X8 FILLER_132_1035 ();
 FILLCELL_X4 FILLER_132_1043 ();
 FILLCELL_X1 FILLER_132_1047 ();
 FILLCELL_X32 FILLER_132_1078 ();
 FILLCELL_X32 FILLER_132_1110 ();
 FILLCELL_X32 FILLER_132_1142 ();
 FILLCELL_X32 FILLER_132_1174 ();
 FILLCELL_X32 FILLER_132_1206 ();
 FILLCELL_X32 FILLER_132_1238 ();
 FILLCELL_X32 FILLER_132_1270 ();
 FILLCELL_X32 FILLER_132_1302 ();
 FILLCELL_X32 FILLER_132_1334 ();
 FILLCELL_X32 FILLER_132_1366 ();
 FILLCELL_X32 FILLER_132_1398 ();
 FILLCELL_X32 FILLER_132_1430 ();
 FILLCELL_X32 FILLER_132_1462 ();
 FILLCELL_X32 FILLER_132_1494 ();
 FILLCELL_X32 FILLER_132_1526 ();
 FILLCELL_X32 FILLER_132_1558 ();
 FILLCELL_X32 FILLER_132_1590 ();
 FILLCELL_X32 FILLER_132_1622 ();
 FILLCELL_X32 FILLER_132_1654 ();
 FILLCELL_X32 FILLER_132_1686 ();
 FILLCELL_X32 FILLER_132_1718 ();
 FILLCELL_X32 FILLER_132_1750 ();
 FILLCELL_X32 FILLER_132_1782 ();
 FILLCELL_X32 FILLER_132_1814 ();
 FILLCELL_X8 FILLER_132_1846 ();
 FILLCELL_X4 FILLER_132_1854 ();
 FILLCELL_X32 FILLER_132_1862 ();
 FILLCELL_X1 FILLER_132_1895 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X16 FILLER_133_801 ();
 FILLCELL_X2 FILLER_133_817 ();
 FILLCELL_X16 FILLER_133_837 ();
 FILLCELL_X4 FILLER_133_855 ();
 FILLCELL_X32 FILLER_133_861 ();
 FILLCELL_X8 FILLER_133_893 ();
 FILLCELL_X4 FILLER_133_911 ();
 FILLCELL_X2 FILLER_133_915 ();
 FILLCELL_X1 FILLER_133_917 ();
 FILLCELL_X1 FILLER_133_922 ();
 FILLCELL_X1 FILLER_133_926 ();
 FILLCELL_X1 FILLER_133_931 ();
 FILLCELL_X4 FILLER_133_945 ();
 FILLCELL_X32 FILLER_133_968 ();
 FILLCELL_X32 FILLER_133_1000 ();
 FILLCELL_X16 FILLER_133_1032 ();
 FILLCELL_X8 FILLER_133_1048 ();
 FILLCELL_X32 FILLER_133_1096 ();
 FILLCELL_X32 FILLER_133_1128 ();
 FILLCELL_X32 FILLER_133_1160 ();
 FILLCELL_X32 FILLER_133_1192 ();
 FILLCELL_X32 FILLER_133_1224 ();
 FILLCELL_X4 FILLER_133_1256 ();
 FILLCELL_X2 FILLER_133_1260 ();
 FILLCELL_X1 FILLER_133_1262 ();
 FILLCELL_X32 FILLER_133_1264 ();
 FILLCELL_X32 FILLER_133_1296 ();
 FILLCELL_X32 FILLER_133_1328 ();
 FILLCELL_X32 FILLER_133_1360 ();
 FILLCELL_X32 FILLER_133_1392 ();
 FILLCELL_X32 FILLER_133_1424 ();
 FILLCELL_X32 FILLER_133_1456 ();
 FILLCELL_X32 FILLER_133_1488 ();
 FILLCELL_X32 FILLER_133_1520 ();
 FILLCELL_X32 FILLER_133_1552 ();
 FILLCELL_X32 FILLER_133_1584 ();
 FILLCELL_X32 FILLER_133_1616 ();
 FILLCELL_X32 FILLER_133_1648 ();
 FILLCELL_X32 FILLER_133_1680 ();
 FILLCELL_X32 FILLER_133_1712 ();
 FILLCELL_X32 FILLER_133_1744 ();
 FILLCELL_X32 FILLER_133_1776 ();
 FILLCELL_X32 FILLER_133_1808 ();
 FILLCELL_X32 FILLER_133_1840 ();
 FILLCELL_X16 FILLER_133_1872 ();
 FILLCELL_X8 FILLER_133_1888 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X16 FILLER_134_792 ();
 FILLCELL_X1 FILLER_134_808 ();
 FILLCELL_X4 FILLER_134_819 ();
 FILLCELL_X2 FILLER_134_823 ();
 FILLCELL_X8 FILLER_134_833 ();
 FILLCELL_X16 FILLER_134_881 ();
 FILLCELL_X4 FILLER_134_897 ();
 FILLCELL_X16 FILLER_134_905 ();
 FILLCELL_X8 FILLER_134_921 ();
 FILLCELL_X1 FILLER_134_929 ();
 FILLCELL_X2 FILLER_134_950 ();
 FILLCELL_X1 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_966 ();
 FILLCELL_X1 FILLER_134_998 ();
 FILLCELL_X4 FILLER_134_1006 ();
 FILLCELL_X2 FILLER_134_1010 ();
 FILLCELL_X1 FILLER_134_1012 ();
 FILLCELL_X8 FILLER_134_1016 ();
 FILLCELL_X2 FILLER_134_1024 ();
 FILLCELL_X1 FILLER_134_1030 ();
 FILLCELL_X2 FILLER_134_1038 ();
 FILLCELL_X1 FILLER_134_1040 ();
 FILLCELL_X2 FILLER_134_1043 ();
 FILLCELL_X1 FILLER_134_1045 ();
 FILLCELL_X8 FILLER_134_1050 ();
 FILLCELL_X4 FILLER_134_1058 ();
 FILLCELL_X2 FILLER_134_1062 ();
 FILLCELL_X32 FILLER_134_1080 ();
 FILLCELL_X32 FILLER_134_1112 ();
 FILLCELL_X32 FILLER_134_1144 ();
 FILLCELL_X32 FILLER_134_1176 ();
 FILLCELL_X32 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_134_1240 ();
 FILLCELL_X32 FILLER_134_1272 ();
 FILLCELL_X32 FILLER_134_1304 ();
 FILLCELL_X32 FILLER_134_1336 ();
 FILLCELL_X32 FILLER_134_1368 ();
 FILLCELL_X32 FILLER_134_1400 ();
 FILLCELL_X32 FILLER_134_1432 ();
 FILLCELL_X32 FILLER_134_1464 ();
 FILLCELL_X32 FILLER_134_1496 ();
 FILLCELL_X32 FILLER_134_1528 ();
 FILLCELL_X32 FILLER_134_1560 ();
 FILLCELL_X32 FILLER_134_1592 ();
 FILLCELL_X32 FILLER_134_1624 ();
 FILLCELL_X32 FILLER_134_1656 ();
 FILLCELL_X32 FILLER_134_1688 ();
 FILLCELL_X32 FILLER_134_1720 ();
 FILLCELL_X32 FILLER_134_1752 ();
 FILLCELL_X32 FILLER_134_1784 ();
 FILLCELL_X32 FILLER_134_1816 ();
 FILLCELL_X32 FILLER_134_1848 ();
 FILLCELL_X8 FILLER_134_1880 ();
 FILLCELL_X4 FILLER_134_1888 ();
 FILLCELL_X2 FILLER_134_1892 ();
 FILLCELL_X1 FILLER_134_1895 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X1 FILLER_135_801 ();
 FILLCELL_X8 FILLER_135_813 ();
 FILLCELL_X4 FILLER_135_821 ();
 FILLCELL_X2 FILLER_135_825 ();
 FILLCELL_X1 FILLER_135_827 ();
 FILLCELL_X2 FILLER_135_837 ();
 FILLCELL_X1 FILLER_135_839 ();
 FILLCELL_X2 FILLER_135_850 ();
 FILLCELL_X1 FILLER_135_852 ();
 FILLCELL_X2 FILLER_135_862 ();
 FILLCELL_X1 FILLER_135_864 ();
 FILLCELL_X32 FILLER_135_874 ();
 FILLCELL_X16 FILLER_135_906 ();
 FILLCELL_X2 FILLER_135_922 ();
 FILLCELL_X1 FILLER_135_924 ();
 FILLCELL_X4 FILLER_135_931 ();
 FILLCELL_X2 FILLER_135_935 ();
 FILLCELL_X16 FILLER_135_940 ();
 FILLCELL_X8 FILLER_135_963 ();
 FILLCELL_X16 FILLER_135_975 ();
 FILLCELL_X8 FILLER_135_991 ();
 FILLCELL_X4 FILLER_135_999 ();
 FILLCELL_X2 FILLER_135_1003 ();
 FILLCELL_X1 FILLER_135_1005 ();
 FILLCELL_X1 FILLER_135_1015 ();
 FILLCELL_X1 FILLER_135_1034 ();
 FILLCELL_X4 FILLER_135_1051 ();
 FILLCELL_X1 FILLER_135_1055 ();
 FILLCELL_X1 FILLER_135_1070 ();
 FILLCELL_X32 FILLER_135_1081 ();
 FILLCELL_X32 FILLER_135_1113 ();
 FILLCELL_X32 FILLER_135_1145 ();
 FILLCELL_X32 FILLER_135_1177 ();
 FILLCELL_X32 FILLER_135_1209 ();
 FILLCELL_X16 FILLER_135_1241 ();
 FILLCELL_X4 FILLER_135_1257 ();
 FILLCELL_X2 FILLER_135_1261 ();
 FILLCELL_X32 FILLER_135_1264 ();
 FILLCELL_X32 FILLER_135_1296 ();
 FILLCELL_X32 FILLER_135_1328 ();
 FILLCELL_X32 FILLER_135_1360 ();
 FILLCELL_X32 FILLER_135_1392 ();
 FILLCELL_X32 FILLER_135_1424 ();
 FILLCELL_X32 FILLER_135_1456 ();
 FILLCELL_X32 FILLER_135_1488 ();
 FILLCELL_X32 FILLER_135_1520 ();
 FILLCELL_X32 FILLER_135_1552 ();
 FILLCELL_X32 FILLER_135_1584 ();
 FILLCELL_X32 FILLER_135_1616 ();
 FILLCELL_X32 FILLER_135_1648 ();
 FILLCELL_X32 FILLER_135_1680 ();
 FILLCELL_X32 FILLER_135_1712 ();
 FILLCELL_X32 FILLER_135_1744 ();
 FILLCELL_X32 FILLER_135_1776 ();
 FILLCELL_X32 FILLER_135_1808 ();
 FILLCELL_X32 FILLER_135_1840 ();
 FILLCELL_X16 FILLER_135_1872 ();
 FILLCELL_X8 FILLER_135_1888 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X4 FILLER_136_792 ();
 FILLCELL_X4 FILLER_136_822 ();
 FILLCELL_X2 FILLER_136_826 ();
 FILLCELL_X1 FILLER_136_828 ();
 FILLCELL_X4 FILLER_136_840 ();
 FILLCELL_X2 FILLER_136_844 ();
 FILLCELL_X1 FILLER_136_846 ();
 FILLCELL_X2 FILLER_136_858 ();
 FILLCELL_X4 FILLER_136_867 ();
 FILLCELL_X2 FILLER_136_871 ();
 FILLCELL_X16 FILLER_136_880 ();
 FILLCELL_X4 FILLER_136_896 ();
 FILLCELL_X1 FILLER_136_900 ();
 FILLCELL_X8 FILLER_136_914 ();
 FILLCELL_X2 FILLER_136_922 ();
 FILLCELL_X16 FILLER_136_930 ();
 FILLCELL_X2 FILLER_136_946 ();
 FILLCELL_X1 FILLER_136_965 ();
 FILLCELL_X1 FILLER_136_980 ();
 FILLCELL_X8 FILLER_136_1001 ();
 FILLCELL_X2 FILLER_136_1009 ();
 FILLCELL_X8 FILLER_136_1016 ();
 FILLCELL_X2 FILLER_136_1028 ();
 FILLCELL_X1 FILLER_136_1030 ();
 FILLCELL_X2 FILLER_136_1048 ();
 FILLCELL_X4 FILLER_136_1056 ();
 FILLCELL_X2 FILLER_136_1060 ();
 FILLCELL_X4 FILLER_136_1068 ();
 FILLCELL_X1 FILLER_136_1072 ();
 FILLCELL_X32 FILLER_136_1077 ();
 FILLCELL_X32 FILLER_136_1109 ();
 FILLCELL_X32 FILLER_136_1141 ();
 FILLCELL_X32 FILLER_136_1173 ();
 FILLCELL_X32 FILLER_136_1205 ();
 FILLCELL_X32 FILLER_136_1237 ();
 FILLCELL_X32 FILLER_136_1269 ();
 FILLCELL_X32 FILLER_136_1301 ();
 FILLCELL_X32 FILLER_136_1333 ();
 FILLCELL_X32 FILLER_136_1365 ();
 FILLCELL_X32 FILLER_136_1397 ();
 FILLCELL_X32 FILLER_136_1429 ();
 FILLCELL_X32 FILLER_136_1461 ();
 FILLCELL_X32 FILLER_136_1493 ();
 FILLCELL_X32 FILLER_136_1525 ();
 FILLCELL_X32 FILLER_136_1557 ();
 FILLCELL_X32 FILLER_136_1589 ();
 FILLCELL_X32 FILLER_136_1621 ();
 FILLCELL_X32 FILLER_136_1653 ();
 FILLCELL_X32 FILLER_136_1685 ();
 FILLCELL_X32 FILLER_136_1717 ();
 FILLCELL_X32 FILLER_136_1749 ();
 FILLCELL_X32 FILLER_136_1781 ();
 FILLCELL_X32 FILLER_136_1813 ();
 FILLCELL_X32 FILLER_136_1845 ();
 FILLCELL_X16 FILLER_136_1877 ();
 FILLCELL_X1 FILLER_136_1893 ();
 FILLCELL_X1 FILLER_136_1895 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X4 FILLER_137_801 ();
 FILLCELL_X1 FILLER_137_805 ();
 FILLCELL_X2 FILLER_137_826 ();
 FILLCELL_X1 FILLER_137_839 ();
 FILLCELL_X4 FILLER_137_845 ();
 FILLCELL_X2 FILLER_137_849 ();
 FILLCELL_X1 FILLER_137_851 ();
 FILLCELL_X4 FILLER_137_863 ();
 FILLCELL_X2 FILLER_137_874 ();
 FILLCELL_X1 FILLER_137_886 ();
 FILLCELL_X2 FILLER_137_904 ();
 FILLCELL_X1 FILLER_137_906 ();
 FILLCELL_X8 FILLER_137_916 ();
 FILLCELL_X2 FILLER_137_924 ();
 FILLCELL_X1 FILLER_137_926 ();
 FILLCELL_X16 FILLER_137_936 ();
 FILLCELL_X1 FILLER_137_952 ();
 FILLCELL_X16 FILLER_137_963 ();
 FILLCELL_X2 FILLER_137_979 ();
 FILLCELL_X16 FILLER_137_994 ();
 FILLCELL_X2 FILLER_137_1010 ();
 FILLCELL_X1 FILLER_137_1012 ();
 FILLCELL_X4 FILLER_137_1018 ();
 FILLCELL_X1 FILLER_137_1022 ();
 FILLCELL_X4 FILLER_137_1029 ();
 FILLCELL_X1 FILLER_137_1033 ();
 FILLCELL_X4 FILLER_137_1040 ();
 FILLCELL_X2 FILLER_137_1044 ();
 FILLCELL_X1 FILLER_137_1046 ();
 FILLCELL_X32 FILLER_137_1056 ();
 FILLCELL_X32 FILLER_137_1088 ();
 FILLCELL_X32 FILLER_137_1120 ();
 FILLCELL_X32 FILLER_137_1152 ();
 FILLCELL_X32 FILLER_137_1184 ();
 FILLCELL_X32 FILLER_137_1216 ();
 FILLCELL_X8 FILLER_137_1248 ();
 FILLCELL_X4 FILLER_137_1256 ();
 FILLCELL_X2 FILLER_137_1260 ();
 FILLCELL_X1 FILLER_137_1262 ();
 FILLCELL_X32 FILLER_137_1264 ();
 FILLCELL_X32 FILLER_137_1296 ();
 FILLCELL_X32 FILLER_137_1328 ();
 FILLCELL_X32 FILLER_137_1360 ();
 FILLCELL_X32 FILLER_137_1392 ();
 FILLCELL_X32 FILLER_137_1424 ();
 FILLCELL_X32 FILLER_137_1456 ();
 FILLCELL_X32 FILLER_137_1488 ();
 FILLCELL_X32 FILLER_137_1520 ();
 FILLCELL_X32 FILLER_137_1552 ();
 FILLCELL_X32 FILLER_137_1584 ();
 FILLCELL_X32 FILLER_137_1616 ();
 FILLCELL_X32 FILLER_137_1648 ();
 FILLCELL_X32 FILLER_137_1680 ();
 FILLCELL_X32 FILLER_137_1712 ();
 FILLCELL_X32 FILLER_137_1744 ();
 FILLCELL_X32 FILLER_137_1776 ();
 FILLCELL_X32 FILLER_137_1808 ();
 FILLCELL_X32 FILLER_137_1840 ();
 FILLCELL_X16 FILLER_137_1872 ();
 FILLCELL_X8 FILLER_137_1888 ();
 FILLCELL_X16 FILLER_138_1 ();
 FILLCELL_X8 FILLER_138_17 ();
 FILLCELL_X4 FILLER_138_25 ();
 FILLCELL_X32 FILLER_138_39 ();
 FILLCELL_X32 FILLER_138_71 ();
 FILLCELL_X32 FILLER_138_103 ();
 FILLCELL_X32 FILLER_138_135 ();
 FILLCELL_X32 FILLER_138_167 ();
 FILLCELL_X32 FILLER_138_199 ();
 FILLCELL_X32 FILLER_138_231 ();
 FILLCELL_X32 FILLER_138_263 ();
 FILLCELL_X32 FILLER_138_295 ();
 FILLCELL_X32 FILLER_138_327 ();
 FILLCELL_X32 FILLER_138_359 ();
 FILLCELL_X32 FILLER_138_391 ();
 FILLCELL_X32 FILLER_138_423 ();
 FILLCELL_X32 FILLER_138_455 ();
 FILLCELL_X32 FILLER_138_487 ();
 FILLCELL_X32 FILLER_138_519 ();
 FILLCELL_X32 FILLER_138_551 ();
 FILLCELL_X32 FILLER_138_583 ();
 FILLCELL_X16 FILLER_138_615 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X8 FILLER_138_824 ();
 FILLCELL_X2 FILLER_138_832 ();
 FILLCELL_X1 FILLER_138_834 ();
 FILLCELL_X8 FILLER_138_848 ();
 FILLCELL_X2 FILLER_138_856 ();
 FILLCELL_X16 FILLER_138_870 ();
 FILLCELL_X2 FILLER_138_886 ();
 FILLCELL_X1 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_901 ();
 FILLCELL_X16 FILLER_138_933 ();
 FILLCELL_X8 FILLER_138_949 ();
 FILLCELL_X32 FILLER_138_970 ();
 FILLCELL_X32 FILLER_138_1002 ();
 FILLCELL_X8 FILLER_138_1034 ();
 FILLCELL_X4 FILLER_138_1042 ();
 FILLCELL_X32 FILLER_138_1055 ();
 FILLCELL_X32 FILLER_138_1087 ();
 FILLCELL_X32 FILLER_138_1119 ();
 FILLCELL_X32 FILLER_138_1151 ();
 FILLCELL_X32 FILLER_138_1183 ();
 FILLCELL_X32 FILLER_138_1215 ();
 FILLCELL_X32 FILLER_138_1247 ();
 FILLCELL_X32 FILLER_138_1279 ();
 FILLCELL_X32 FILLER_138_1311 ();
 FILLCELL_X32 FILLER_138_1343 ();
 FILLCELL_X32 FILLER_138_1375 ();
 FILLCELL_X32 FILLER_138_1407 ();
 FILLCELL_X32 FILLER_138_1439 ();
 FILLCELL_X32 FILLER_138_1471 ();
 FILLCELL_X32 FILLER_138_1503 ();
 FILLCELL_X32 FILLER_138_1535 ();
 FILLCELL_X32 FILLER_138_1567 ();
 FILLCELL_X32 FILLER_138_1599 ();
 FILLCELL_X32 FILLER_138_1631 ();
 FILLCELL_X32 FILLER_138_1663 ();
 FILLCELL_X32 FILLER_138_1695 ();
 FILLCELL_X32 FILLER_138_1727 ();
 FILLCELL_X32 FILLER_138_1759 ();
 FILLCELL_X32 FILLER_138_1791 ();
 FILLCELL_X32 FILLER_138_1823 ();
 FILLCELL_X32 FILLER_138_1855 ();
 FILLCELL_X4 FILLER_138_1887 ();
 FILLCELL_X2 FILLER_138_1891 ();
 FILLCELL_X1 FILLER_138_1893 ();
 FILLCELL_X1 FILLER_138_1895 ();
 FILLCELL_X8 FILLER_139_1 ();
 FILLCELL_X2 FILLER_139_9 ();
 FILLCELL_X32 FILLER_139_15 ();
 FILLCELL_X32 FILLER_139_47 ();
 FILLCELL_X32 FILLER_139_79 ();
 FILLCELL_X32 FILLER_139_111 ();
 FILLCELL_X32 FILLER_139_143 ();
 FILLCELL_X32 FILLER_139_175 ();
 FILLCELL_X32 FILLER_139_207 ();
 FILLCELL_X32 FILLER_139_239 ();
 FILLCELL_X32 FILLER_139_271 ();
 FILLCELL_X32 FILLER_139_303 ();
 FILLCELL_X32 FILLER_139_335 ();
 FILLCELL_X32 FILLER_139_367 ();
 FILLCELL_X32 FILLER_139_399 ();
 FILLCELL_X32 FILLER_139_431 ();
 FILLCELL_X32 FILLER_139_463 ();
 FILLCELL_X32 FILLER_139_495 ();
 FILLCELL_X32 FILLER_139_527 ();
 FILLCELL_X32 FILLER_139_559 ();
 FILLCELL_X32 FILLER_139_591 ();
 FILLCELL_X32 FILLER_139_623 ();
 FILLCELL_X32 FILLER_139_655 ();
 FILLCELL_X32 FILLER_139_687 ();
 FILLCELL_X32 FILLER_139_719 ();
 FILLCELL_X32 FILLER_139_751 ();
 FILLCELL_X32 FILLER_139_783 ();
 FILLCELL_X32 FILLER_139_815 ();
 FILLCELL_X32 FILLER_139_847 ();
 FILLCELL_X32 FILLER_139_879 ();
 FILLCELL_X32 FILLER_139_911 ();
 FILLCELL_X32 FILLER_139_943 ();
 FILLCELL_X32 FILLER_139_975 ();
 FILLCELL_X32 FILLER_139_1007 ();
 FILLCELL_X32 FILLER_139_1039 ();
 FILLCELL_X32 FILLER_139_1071 ();
 FILLCELL_X32 FILLER_139_1103 ();
 FILLCELL_X32 FILLER_139_1135 ();
 FILLCELL_X32 FILLER_139_1167 ();
 FILLCELL_X32 FILLER_139_1199 ();
 FILLCELL_X32 FILLER_139_1231 ();
 FILLCELL_X32 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1296 ();
 FILLCELL_X32 FILLER_139_1328 ();
 FILLCELL_X32 FILLER_139_1360 ();
 FILLCELL_X32 FILLER_139_1392 ();
 FILLCELL_X32 FILLER_139_1424 ();
 FILLCELL_X32 FILLER_139_1456 ();
 FILLCELL_X32 FILLER_139_1488 ();
 FILLCELL_X32 FILLER_139_1520 ();
 FILLCELL_X32 FILLER_139_1552 ();
 FILLCELL_X32 FILLER_139_1584 ();
 FILLCELL_X32 FILLER_139_1616 ();
 FILLCELL_X32 FILLER_139_1648 ();
 FILLCELL_X32 FILLER_139_1680 ();
 FILLCELL_X32 FILLER_139_1712 ();
 FILLCELL_X32 FILLER_139_1744 ();
 FILLCELL_X32 FILLER_139_1776 ();
 FILLCELL_X32 FILLER_139_1808 ();
 FILLCELL_X32 FILLER_139_1840 ();
 FILLCELL_X16 FILLER_139_1872 ();
 FILLCELL_X8 FILLER_139_1888 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X32 FILLER_140_1048 ();
 FILLCELL_X32 FILLER_140_1080 ();
 FILLCELL_X32 FILLER_140_1112 ();
 FILLCELL_X32 FILLER_140_1144 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X32 FILLER_140_1240 ();
 FILLCELL_X32 FILLER_140_1272 ();
 FILLCELL_X32 FILLER_140_1304 ();
 FILLCELL_X32 FILLER_140_1336 ();
 FILLCELL_X32 FILLER_140_1368 ();
 FILLCELL_X32 FILLER_140_1400 ();
 FILLCELL_X32 FILLER_140_1432 ();
 FILLCELL_X32 FILLER_140_1464 ();
 FILLCELL_X32 FILLER_140_1496 ();
 FILLCELL_X32 FILLER_140_1528 ();
 FILLCELL_X32 FILLER_140_1560 ();
 FILLCELL_X32 FILLER_140_1592 ();
 FILLCELL_X32 FILLER_140_1624 ();
 FILLCELL_X32 FILLER_140_1656 ();
 FILLCELL_X32 FILLER_140_1688 ();
 FILLCELL_X32 FILLER_140_1720 ();
 FILLCELL_X32 FILLER_140_1752 ();
 FILLCELL_X32 FILLER_140_1784 ();
 FILLCELL_X32 FILLER_140_1816 ();
 FILLCELL_X32 FILLER_140_1848 ();
 FILLCELL_X8 FILLER_140_1880 ();
 FILLCELL_X4 FILLER_140_1888 ();
 FILLCELL_X2 FILLER_140_1892 ();
 FILLCELL_X1 FILLER_140_1895 ();
 FILLCELL_X32 FILLER_141_6 ();
 FILLCELL_X32 FILLER_141_38 ();
 FILLCELL_X32 FILLER_141_70 ();
 FILLCELL_X32 FILLER_141_102 ();
 FILLCELL_X32 FILLER_141_134 ();
 FILLCELL_X32 FILLER_141_166 ();
 FILLCELL_X32 FILLER_141_198 ();
 FILLCELL_X32 FILLER_141_230 ();
 FILLCELL_X32 FILLER_141_262 ();
 FILLCELL_X32 FILLER_141_294 ();
 FILLCELL_X32 FILLER_141_326 ();
 FILLCELL_X32 FILLER_141_358 ();
 FILLCELL_X32 FILLER_141_390 ();
 FILLCELL_X32 FILLER_141_422 ();
 FILLCELL_X32 FILLER_141_454 ();
 FILLCELL_X32 FILLER_141_486 ();
 FILLCELL_X32 FILLER_141_518 ();
 FILLCELL_X32 FILLER_141_550 ();
 FILLCELL_X32 FILLER_141_582 ();
 FILLCELL_X32 FILLER_141_614 ();
 FILLCELL_X32 FILLER_141_646 ();
 FILLCELL_X32 FILLER_141_678 ();
 FILLCELL_X32 FILLER_141_710 ();
 FILLCELL_X32 FILLER_141_742 ();
 FILLCELL_X32 FILLER_141_774 ();
 FILLCELL_X32 FILLER_141_806 ();
 FILLCELL_X32 FILLER_141_838 ();
 FILLCELL_X32 FILLER_141_870 ();
 FILLCELL_X32 FILLER_141_902 ();
 FILLCELL_X32 FILLER_141_934 ();
 FILLCELL_X32 FILLER_141_966 ();
 FILLCELL_X32 FILLER_141_998 ();
 FILLCELL_X32 FILLER_141_1030 ();
 FILLCELL_X32 FILLER_141_1062 ();
 FILLCELL_X32 FILLER_141_1094 ();
 FILLCELL_X32 FILLER_141_1126 ();
 FILLCELL_X32 FILLER_141_1158 ();
 FILLCELL_X32 FILLER_141_1190 ();
 FILLCELL_X32 FILLER_141_1222 ();
 FILLCELL_X8 FILLER_141_1254 ();
 FILLCELL_X1 FILLER_141_1262 ();
 FILLCELL_X32 FILLER_141_1264 ();
 FILLCELL_X32 FILLER_141_1296 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X32 FILLER_141_1360 ();
 FILLCELL_X32 FILLER_141_1392 ();
 FILLCELL_X32 FILLER_141_1424 ();
 FILLCELL_X32 FILLER_141_1456 ();
 FILLCELL_X32 FILLER_141_1488 ();
 FILLCELL_X32 FILLER_141_1520 ();
 FILLCELL_X32 FILLER_141_1552 ();
 FILLCELL_X32 FILLER_141_1584 ();
 FILLCELL_X32 FILLER_141_1616 ();
 FILLCELL_X32 FILLER_141_1648 ();
 FILLCELL_X32 FILLER_141_1680 ();
 FILLCELL_X32 FILLER_141_1712 ();
 FILLCELL_X32 FILLER_141_1744 ();
 FILLCELL_X32 FILLER_141_1776 ();
 FILLCELL_X32 FILLER_141_1808 ();
 FILLCELL_X32 FILLER_141_1840 ();
 FILLCELL_X16 FILLER_141_1872 ();
 FILLCELL_X8 FILLER_141_1888 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X32 FILLER_142_1112 ();
 FILLCELL_X32 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_142_1176 ();
 FILLCELL_X32 FILLER_142_1208 ();
 FILLCELL_X32 FILLER_142_1240 ();
 FILLCELL_X32 FILLER_142_1272 ();
 FILLCELL_X32 FILLER_142_1304 ();
 FILLCELL_X32 FILLER_142_1336 ();
 FILLCELL_X32 FILLER_142_1368 ();
 FILLCELL_X32 FILLER_142_1400 ();
 FILLCELL_X32 FILLER_142_1432 ();
 FILLCELL_X32 FILLER_142_1464 ();
 FILLCELL_X32 FILLER_142_1496 ();
 FILLCELL_X32 FILLER_142_1528 ();
 FILLCELL_X32 FILLER_142_1560 ();
 FILLCELL_X32 FILLER_142_1592 ();
 FILLCELL_X32 FILLER_142_1624 ();
 FILLCELL_X32 FILLER_142_1656 ();
 FILLCELL_X32 FILLER_142_1688 ();
 FILLCELL_X32 FILLER_142_1720 ();
 FILLCELL_X32 FILLER_142_1752 ();
 FILLCELL_X32 FILLER_142_1784 ();
 FILLCELL_X32 FILLER_142_1816 ();
 FILLCELL_X32 FILLER_142_1848 ();
 FILLCELL_X8 FILLER_142_1880 ();
 FILLCELL_X4 FILLER_142_1888 ();
 FILLCELL_X2 FILLER_142_1892 ();
 FILLCELL_X1 FILLER_142_1895 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X32 FILLER_143_1089 ();
 FILLCELL_X32 FILLER_143_1121 ();
 FILLCELL_X32 FILLER_143_1153 ();
 FILLCELL_X32 FILLER_143_1185 ();
 FILLCELL_X32 FILLER_143_1217 ();
 FILLCELL_X8 FILLER_143_1249 ();
 FILLCELL_X4 FILLER_143_1257 ();
 FILLCELL_X2 FILLER_143_1261 ();
 FILLCELL_X32 FILLER_143_1264 ();
 FILLCELL_X32 FILLER_143_1296 ();
 FILLCELL_X32 FILLER_143_1328 ();
 FILLCELL_X32 FILLER_143_1360 ();
 FILLCELL_X32 FILLER_143_1392 ();
 FILLCELL_X32 FILLER_143_1424 ();
 FILLCELL_X32 FILLER_143_1456 ();
 FILLCELL_X32 FILLER_143_1488 ();
 FILLCELL_X32 FILLER_143_1520 ();
 FILLCELL_X32 FILLER_143_1552 ();
 FILLCELL_X32 FILLER_143_1584 ();
 FILLCELL_X32 FILLER_143_1616 ();
 FILLCELL_X32 FILLER_143_1648 ();
 FILLCELL_X32 FILLER_143_1680 ();
 FILLCELL_X32 FILLER_143_1712 ();
 FILLCELL_X32 FILLER_143_1744 ();
 FILLCELL_X32 FILLER_143_1776 ();
 FILLCELL_X32 FILLER_143_1808 ();
 FILLCELL_X32 FILLER_143_1840 ();
 FILLCELL_X16 FILLER_143_1872 ();
 FILLCELL_X8 FILLER_143_1888 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X32 FILLER_144_1144 ();
 FILLCELL_X32 FILLER_144_1176 ();
 FILLCELL_X32 FILLER_144_1208 ();
 FILLCELL_X32 FILLER_144_1240 ();
 FILLCELL_X32 FILLER_144_1272 ();
 FILLCELL_X32 FILLER_144_1304 ();
 FILLCELL_X32 FILLER_144_1336 ();
 FILLCELL_X32 FILLER_144_1368 ();
 FILLCELL_X32 FILLER_144_1400 ();
 FILLCELL_X32 FILLER_144_1432 ();
 FILLCELL_X32 FILLER_144_1464 ();
 FILLCELL_X32 FILLER_144_1496 ();
 FILLCELL_X32 FILLER_144_1528 ();
 FILLCELL_X32 FILLER_144_1560 ();
 FILLCELL_X32 FILLER_144_1592 ();
 FILLCELL_X32 FILLER_144_1624 ();
 FILLCELL_X32 FILLER_144_1656 ();
 FILLCELL_X32 FILLER_144_1688 ();
 FILLCELL_X32 FILLER_144_1720 ();
 FILLCELL_X32 FILLER_144_1752 ();
 FILLCELL_X32 FILLER_144_1784 ();
 FILLCELL_X32 FILLER_144_1816 ();
 FILLCELL_X32 FILLER_144_1848 ();
 FILLCELL_X8 FILLER_144_1880 ();
 FILLCELL_X4 FILLER_144_1888 ();
 FILLCELL_X2 FILLER_144_1892 ();
 FILLCELL_X1 FILLER_144_1895 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X32 FILLER_145_1153 ();
 FILLCELL_X32 FILLER_145_1185 ();
 FILLCELL_X32 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1249 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X32 FILLER_145_1584 ();
 FILLCELL_X32 FILLER_145_1616 ();
 FILLCELL_X32 FILLER_145_1648 ();
 FILLCELL_X32 FILLER_145_1680 ();
 FILLCELL_X32 FILLER_145_1712 ();
 FILLCELL_X32 FILLER_145_1744 ();
 FILLCELL_X32 FILLER_145_1776 ();
 FILLCELL_X32 FILLER_145_1808 ();
 FILLCELL_X32 FILLER_145_1840 ();
 FILLCELL_X16 FILLER_145_1872 ();
 FILLCELL_X8 FILLER_145_1888 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X32 FILLER_146_1144 ();
 FILLCELL_X32 FILLER_146_1176 ();
 FILLCELL_X32 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_146_1240 ();
 FILLCELL_X32 FILLER_146_1272 ();
 FILLCELL_X32 FILLER_146_1304 ();
 FILLCELL_X32 FILLER_146_1336 ();
 FILLCELL_X32 FILLER_146_1368 ();
 FILLCELL_X32 FILLER_146_1400 ();
 FILLCELL_X32 FILLER_146_1432 ();
 FILLCELL_X32 FILLER_146_1464 ();
 FILLCELL_X32 FILLER_146_1496 ();
 FILLCELL_X32 FILLER_146_1528 ();
 FILLCELL_X32 FILLER_146_1560 ();
 FILLCELL_X32 FILLER_146_1592 ();
 FILLCELL_X32 FILLER_146_1624 ();
 FILLCELL_X32 FILLER_146_1656 ();
 FILLCELL_X32 FILLER_146_1688 ();
 FILLCELL_X32 FILLER_146_1720 ();
 FILLCELL_X32 FILLER_146_1752 ();
 FILLCELL_X32 FILLER_146_1784 ();
 FILLCELL_X32 FILLER_146_1816 ();
 FILLCELL_X32 FILLER_146_1848 ();
 FILLCELL_X8 FILLER_146_1880 ();
 FILLCELL_X4 FILLER_146_1888 ();
 FILLCELL_X2 FILLER_146_1892 ();
 FILLCELL_X1 FILLER_146_1895 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X32 FILLER_147_1185 ();
 FILLCELL_X32 FILLER_147_1217 ();
 FILLCELL_X8 FILLER_147_1249 ();
 FILLCELL_X4 FILLER_147_1257 ();
 FILLCELL_X2 FILLER_147_1261 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X32 FILLER_147_1584 ();
 FILLCELL_X32 FILLER_147_1616 ();
 FILLCELL_X32 FILLER_147_1648 ();
 FILLCELL_X32 FILLER_147_1680 ();
 FILLCELL_X32 FILLER_147_1712 ();
 FILLCELL_X32 FILLER_147_1744 ();
 FILLCELL_X32 FILLER_147_1776 ();
 FILLCELL_X32 FILLER_147_1808 ();
 FILLCELL_X32 FILLER_147_1840 ();
 FILLCELL_X16 FILLER_147_1872 ();
 FILLCELL_X8 FILLER_147_1888 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X32 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_148_1240 ();
 FILLCELL_X32 FILLER_148_1272 ();
 FILLCELL_X32 FILLER_148_1304 ();
 FILLCELL_X32 FILLER_148_1336 ();
 FILLCELL_X32 FILLER_148_1368 ();
 FILLCELL_X32 FILLER_148_1400 ();
 FILLCELL_X32 FILLER_148_1432 ();
 FILLCELL_X32 FILLER_148_1464 ();
 FILLCELL_X32 FILLER_148_1496 ();
 FILLCELL_X32 FILLER_148_1528 ();
 FILLCELL_X32 FILLER_148_1560 ();
 FILLCELL_X32 FILLER_148_1592 ();
 FILLCELL_X32 FILLER_148_1624 ();
 FILLCELL_X32 FILLER_148_1656 ();
 FILLCELL_X32 FILLER_148_1688 ();
 FILLCELL_X32 FILLER_148_1720 ();
 FILLCELL_X32 FILLER_148_1752 ();
 FILLCELL_X32 FILLER_148_1784 ();
 FILLCELL_X32 FILLER_148_1816 ();
 FILLCELL_X32 FILLER_148_1848 ();
 FILLCELL_X8 FILLER_148_1880 ();
 FILLCELL_X4 FILLER_148_1888 ();
 FILLCELL_X2 FILLER_148_1892 ();
 FILLCELL_X1 FILLER_148_1895 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X32 FILLER_149_1584 ();
 FILLCELL_X32 FILLER_149_1616 ();
 FILLCELL_X32 FILLER_149_1648 ();
 FILLCELL_X32 FILLER_149_1680 ();
 FILLCELL_X32 FILLER_149_1712 ();
 FILLCELL_X32 FILLER_149_1744 ();
 FILLCELL_X32 FILLER_149_1776 ();
 FILLCELL_X32 FILLER_149_1808 ();
 FILLCELL_X32 FILLER_149_1840 ();
 FILLCELL_X16 FILLER_149_1872 ();
 FILLCELL_X8 FILLER_149_1888 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X32 FILLER_150_1304 ();
 FILLCELL_X32 FILLER_150_1336 ();
 FILLCELL_X32 FILLER_150_1368 ();
 FILLCELL_X32 FILLER_150_1400 ();
 FILLCELL_X32 FILLER_150_1432 ();
 FILLCELL_X32 FILLER_150_1464 ();
 FILLCELL_X32 FILLER_150_1496 ();
 FILLCELL_X32 FILLER_150_1528 ();
 FILLCELL_X32 FILLER_150_1560 ();
 FILLCELL_X32 FILLER_150_1592 ();
 FILLCELL_X32 FILLER_150_1624 ();
 FILLCELL_X32 FILLER_150_1656 ();
 FILLCELL_X32 FILLER_150_1688 ();
 FILLCELL_X32 FILLER_150_1720 ();
 FILLCELL_X32 FILLER_150_1752 ();
 FILLCELL_X32 FILLER_150_1784 ();
 FILLCELL_X32 FILLER_150_1816 ();
 FILLCELL_X32 FILLER_150_1848 ();
 FILLCELL_X8 FILLER_150_1880 ();
 FILLCELL_X4 FILLER_150_1888 ();
 FILLCELL_X2 FILLER_150_1892 ();
 FILLCELL_X1 FILLER_150_1895 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X32 FILLER_151_1025 ();
 FILLCELL_X32 FILLER_151_1057 ();
 FILLCELL_X32 FILLER_151_1089 ();
 FILLCELL_X32 FILLER_151_1121 ();
 FILLCELL_X32 FILLER_151_1153 ();
 FILLCELL_X32 FILLER_151_1185 ();
 FILLCELL_X32 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1249 ();
 FILLCELL_X4 FILLER_151_1257 ();
 FILLCELL_X2 FILLER_151_1261 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X32 FILLER_151_1648 ();
 FILLCELL_X32 FILLER_151_1680 ();
 FILLCELL_X32 FILLER_151_1712 ();
 FILLCELL_X32 FILLER_151_1744 ();
 FILLCELL_X32 FILLER_151_1776 ();
 FILLCELL_X32 FILLER_151_1808 ();
 FILLCELL_X32 FILLER_151_1840 ();
 FILLCELL_X16 FILLER_151_1872 ();
 FILLCELL_X8 FILLER_151_1888 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X32 FILLER_152_1304 ();
 FILLCELL_X32 FILLER_152_1336 ();
 FILLCELL_X32 FILLER_152_1368 ();
 FILLCELL_X32 FILLER_152_1400 ();
 FILLCELL_X32 FILLER_152_1432 ();
 FILLCELL_X32 FILLER_152_1464 ();
 FILLCELL_X32 FILLER_152_1496 ();
 FILLCELL_X32 FILLER_152_1528 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X32 FILLER_152_1592 ();
 FILLCELL_X32 FILLER_152_1624 ();
 FILLCELL_X32 FILLER_152_1656 ();
 FILLCELL_X32 FILLER_152_1688 ();
 FILLCELL_X32 FILLER_152_1720 ();
 FILLCELL_X32 FILLER_152_1752 ();
 FILLCELL_X32 FILLER_152_1784 ();
 FILLCELL_X32 FILLER_152_1816 ();
 FILLCELL_X32 FILLER_152_1848 ();
 FILLCELL_X8 FILLER_152_1880 ();
 FILLCELL_X4 FILLER_152_1888 ();
 FILLCELL_X2 FILLER_152_1892 ();
 FILLCELL_X1 FILLER_152_1895 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X32 FILLER_153_961 ();
 FILLCELL_X32 FILLER_153_993 ();
 FILLCELL_X32 FILLER_153_1025 ();
 FILLCELL_X32 FILLER_153_1057 ();
 FILLCELL_X32 FILLER_153_1089 ();
 FILLCELL_X32 FILLER_153_1121 ();
 FILLCELL_X32 FILLER_153_1153 ();
 FILLCELL_X32 FILLER_153_1185 ();
 FILLCELL_X32 FILLER_153_1217 ();
 FILLCELL_X8 FILLER_153_1249 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X32 FILLER_153_1584 ();
 FILLCELL_X32 FILLER_153_1616 ();
 FILLCELL_X32 FILLER_153_1648 ();
 FILLCELL_X32 FILLER_153_1680 ();
 FILLCELL_X32 FILLER_153_1712 ();
 FILLCELL_X32 FILLER_153_1744 ();
 FILLCELL_X32 FILLER_153_1776 ();
 FILLCELL_X32 FILLER_153_1808 ();
 FILLCELL_X32 FILLER_153_1840 ();
 FILLCELL_X16 FILLER_153_1872 ();
 FILLCELL_X8 FILLER_153_1888 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X32 FILLER_154_1304 ();
 FILLCELL_X32 FILLER_154_1336 ();
 FILLCELL_X32 FILLER_154_1368 ();
 FILLCELL_X32 FILLER_154_1400 ();
 FILLCELL_X32 FILLER_154_1432 ();
 FILLCELL_X32 FILLER_154_1464 ();
 FILLCELL_X32 FILLER_154_1496 ();
 FILLCELL_X32 FILLER_154_1528 ();
 FILLCELL_X32 FILLER_154_1560 ();
 FILLCELL_X32 FILLER_154_1592 ();
 FILLCELL_X32 FILLER_154_1624 ();
 FILLCELL_X32 FILLER_154_1656 ();
 FILLCELL_X32 FILLER_154_1688 ();
 FILLCELL_X32 FILLER_154_1720 ();
 FILLCELL_X32 FILLER_154_1752 ();
 FILLCELL_X32 FILLER_154_1784 ();
 FILLCELL_X32 FILLER_154_1816 ();
 FILLCELL_X32 FILLER_154_1848 ();
 FILLCELL_X8 FILLER_154_1880 ();
 FILLCELL_X4 FILLER_154_1888 ();
 FILLCELL_X2 FILLER_154_1892 ();
 FILLCELL_X1 FILLER_154_1895 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X32 FILLER_155_929 ();
 FILLCELL_X32 FILLER_155_961 ();
 FILLCELL_X32 FILLER_155_993 ();
 FILLCELL_X32 FILLER_155_1025 ();
 FILLCELL_X32 FILLER_155_1057 ();
 FILLCELL_X32 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1121 ();
 FILLCELL_X32 FILLER_155_1153 ();
 FILLCELL_X32 FILLER_155_1185 ();
 FILLCELL_X32 FILLER_155_1217 ();
 FILLCELL_X8 FILLER_155_1249 ();
 FILLCELL_X4 FILLER_155_1257 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X32 FILLER_155_1584 ();
 FILLCELL_X32 FILLER_155_1616 ();
 FILLCELL_X32 FILLER_155_1648 ();
 FILLCELL_X32 FILLER_155_1680 ();
 FILLCELL_X32 FILLER_155_1712 ();
 FILLCELL_X32 FILLER_155_1744 ();
 FILLCELL_X32 FILLER_155_1776 ();
 FILLCELL_X32 FILLER_155_1808 ();
 FILLCELL_X32 FILLER_155_1840 ();
 FILLCELL_X16 FILLER_155_1872 ();
 FILLCELL_X8 FILLER_155_1888 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X32 FILLER_156_1080 ();
 FILLCELL_X32 FILLER_156_1112 ();
 FILLCELL_X32 FILLER_156_1144 ();
 FILLCELL_X32 FILLER_156_1176 ();
 FILLCELL_X32 FILLER_156_1208 ();
 FILLCELL_X32 FILLER_156_1240 ();
 FILLCELL_X32 FILLER_156_1272 ();
 FILLCELL_X32 FILLER_156_1304 ();
 FILLCELL_X32 FILLER_156_1336 ();
 FILLCELL_X32 FILLER_156_1368 ();
 FILLCELL_X32 FILLER_156_1400 ();
 FILLCELL_X32 FILLER_156_1432 ();
 FILLCELL_X32 FILLER_156_1464 ();
 FILLCELL_X32 FILLER_156_1496 ();
 FILLCELL_X32 FILLER_156_1528 ();
 FILLCELL_X32 FILLER_156_1560 ();
 FILLCELL_X32 FILLER_156_1592 ();
 FILLCELL_X32 FILLER_156_1624 ();
 FILLCELL_X32 FILLER_156_1656 ();
 FILLCELL_X32 FILLER_156_1688 ();
 FILLCELL_X32 FILLER_156_1720 ();
 FILLCELL_X32 FILLER_156_1752 ();
 FILLCELL_X32 FILLER_156_1784 ();
 FILLCELL_X32 FILLER_156_1816 ();
 FILLCELL_X32 FILLER_156_1848 ();
 FILLCELL_X8 FILLER_156_1880 ();
 FILLCELL_X4 FILLER_156_1888 ();
 FILLCELL_X2 FILLER_156_1892 ();
 FILLCELL_X1 FILLER_156_1895 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X32 FILLER_157_929 ();
 FILLCELL_X32 FILLER_157_961 ();
 FILLCELL_X32 FILLER_157_993 ();
 FILLCELL_X32 FILLER_157_1025 ();
 FILLCELL_X32 FILLER_157_1057 ();
 FILLCELL_X32 FILLER_157_1089 ();
 FILLCELL_X32 FILLER_157_1121 ();
 FILLCELL_X32 FILLER_157_1153 ();
 FILLCELL_X32 FILLER_157_1185 ();
 FILLCELL_X32 FILLER_157_1217 ();
 FILLCELL_X8 FILLER_157_1249 ();
 FILLCELL_X4 FILLER_157_1257 ();
 FILLCELL_X2 FILLER_157_1261 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X32 FILLER_157_1584 ();
 FILLCELL_X32 FILLER_157_1616 ();
 FILLCELL_X32 FILLER_157_1648 ();
 FILLCELL_X32 FILLER_157_1680 ();
 FILLCELL_X32 FILLER_157_1712 ();
 FILLCELL_X32 FILLER_157_1744 ();
 FILLCELL_X32 FILLER_157_1776 ();
 FILLCELL_X32 FILLER_157_1808 ();
 FILLCELL_X32 FILLER_157_1840 ();
 FILLCELL_X16 FILLER_157_1872 ();
 FILLCELL_X8 FILLER_157_1888 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X32 FILLER_158_1304 ();
 FILLCELL_X32 FILLER_158_1336 ();
 FILLCELL_X32 FILLER_158_1368 ();
 FILLCELL_X32 FILLER_158_1400 ();
 FILLCELL_X32 FILLER_158_1432 ();
 FILLCELL_X32 FILLER_158_1464 ();
 FILLCELL_X32 FILLER_158_1496 ();
 FILLCELL_X32 FILLER_158_1528 ();
 FILLCELL_X32 FILLER_158_1560 ();
 FILLCELL_X32 FILLER_158_1592 ();
 FILLCELL_X32 FILLER_158_1624 ();
 FILLCELL_X32 FILLER_158_1656 ();
 FILLCELL_X32 FILLER_158_1688 ();
 FILLCELL_X32 FILLER_158_1720 ();
 FILLCELL_X32 FILLER_158_1752 ();
 FILLCELL_X32 FILLER_158_1784 ();
 FILLCELL_X32 FILLER_158_1816 ();
 FILLCELL_X32 FILLER_158_1848 ();
 FILLCELL_X8 FILLER_158_1880 ();
 FILLCELL_X4 FILLER_158_1888 ();
 FILLCELL_X2 FILLER_158_1892 ();
 FILLCELL_X1 FILLER_158_1895 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X32 FILLER_159_929 ();
 FILLCELL_X32 FILLER_159_961 ();
 FILLCELL_X32 FILLER_159_993 ();
 FILLCELL_X32 FILLER_159_1025 ();
 FILLCELL_X32 FILLER_159_1057 ();
 FILLCELL_X32 FILLER_159_1089 ();
 FILLCELL_X32 FILLER_159_1121 ();
 FILLCELL_X32 FILLER_159_1153 ();
 FILLCELL_X32 FILLER_159_1185 ();
 FILLCELL_X32 FILLER_159_1217 ();
 FILLCELL_X8 FILLER_159_1249 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X32 FILLER_159_1584 ();
 FILLCELL_X32 FILLER_159_1616 ();
 FILLCELL_X32 FILLER_159_1648 ();
 FILLCELL_X32 FILLER_159_1680 ();
 FILLCELL_X32 FILLER_159_1712 ();
 FILLCELL_X32 FILLER_159_1744 ();
 FILLCELL_X32 FILLER_159_1776 ();
 FILLCELL_X32 FILLER_159_1808 ();
 FILLCELL_X32 FILLER_159_1840 ();
 FILLCELL_X16 FILLER_159_1872 ();
 FILLCELL_X8 FILLER_159_1888 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X32 FILLER_160_1304 ();
 FILLCELL_X32 FILLER_160_1336 ();
 FILLCELL_X32 FILLER_160_1368 ();
 FILLCELL_X32 FILLER_160_1400 ();
 FILLCELL_X32 FILLER_160_1432 ();
 FILLCELL_X32 FILLER_160_1464 ();
 FILLCELL_X32 FILLER_160_1496 ();
 FILLCELL_X32 FILLER_160_1528 ();
 FILLCELL_X32 FILLER_160_1560 ();
 FILLCELL_X32 FILLER_160_1592 ();
 FILLCELL_X32 FILLER_160_1624 ();
 FILLCELL_X32 FILLER_160_1656 ();
 FILLCELL_X32 FILLER_160_1688 ();
 FILLCELL_X32 FILLER_160_1720 ();
 FILLCELL_X32 FILLER_160_1752 ();
 FILLCELL_X32 FILLER_160_1784 ();
 FILLCELL_X32 FILLER_160_1816 ();
 FILLCELL_X32 FILLER_160_1848 ();
 FILLCELL_X8 FILLER_160_1880 ();
 FILLCELL_X4 FILLER_160_1888 ();
 FILLCELL_X2 FILLER_160_1892 ();
 FILLCELL_X1 FILLER_160_1895 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X32 FILLER_161_993 ();
 FILLCELL_X32 FILLER_161_1025 ();
 FILLCELL_X32 FILLER_161_1057 ();
 FILLCELL_X32 FILLER_161_1089 ();
 FILLCELL_X32 FILLER_161_1121 ();
 FILLCELL_X32 FILLER_161_1153 ();
 FILLCELL_X32 FILLER_161_1185 ();
 FILLCELL_X32 FILLER_161_1217 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X32 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1520 ();
 FILLCELL_X32 FILLER_161_1552 ();
 FILLCELL_X32 FILLER_161_1584 ();
 FILLCELL_X32 FILLER_161_1616 ();
 FILLCELL_X32 FILLER_161_1648 ();
 FILLCELL_X32 FILLER_161_1680 ();
 FILLCELL_X32 FILLER_161_1712 ();
 FILLCELL_X32 FILLER_161_1744 ();
 FILLCELL_X32 FILLER_161_1776 ();
 FILLCELL_X32 FILLER_161_1808 ();
 FILLCELL_X32 FILLER_161_1840 ();
 FILLCELL_X16 FILLER_161_1872 ();
 FILLCELL_X8 FILLER_161_1888 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X32 FILLER_162_1304 ();
 FILLCELL_X32 FILLER_162_1336 ();
 FILLCELL_X32 FILLER_162_1368 ();
 FILLCELL_X32 FILLER_162_1400 ();
 FILLCELL_X32 FILLER_162_1432 ();
 FILLCELL_X32 FILLER_162_1464 ();
 FILLCELL_X32 FILLER_162_1496 ();
 FILLCELL_X32 FILLER_162_1528 ();
 FILLCELL_X32 FILLER_162_1560 ();
 FILLCELL_X32 FILLER_162_1592 ();
 FILLCELL_X32 FILLER_162_1624 ();
 FILLCELL_X32 FILLER_162_1656 ();
 FILLCELL_X32 FILLER_162_1688 ();
 FILLCELL_X32 FILLER_162_1720 ();
 FILLCELL_X32 FILLER_162_1752 ();
 FILLCELL_X32 FILLER_162_1784 ();
 FILLCELL_X32 FILLER_162_1816 ();
 FILLCELL_X32 FILLER_162_1848 ();
 FILLCELL_X8 FILLER_162_1880 ();
 FILLCELL_X4 FILLER_162_1888 ();
 FILLCELL_X2 FILLER_162_1892 ();
 FILLCELL_X1 FILLER_162_1895 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X32 FILLER_163_961 ();
 FILLCELL_X32 FILLER_163_993 ();
 FILLCELL_X32 FILLER_163_1025 ();
 FILLCELL_X32 FILLER_163_1057 ();
 FILLCELL_X32 FILLER_163_1089 ();
 FILLCELL_X32 FILLER_163_1121 ();
 FILLCELL_X32 FILLER_163_1153 ();
 FILLCELL_X32 FILLER_163_1185 ();
 FILLCELL_X32 FILLER_163_1217 ();
 FILLCELL_X8 FILLER_163_1249 ();
 FILLCELL_X4 FILLER_163_1257 ();
 FILLCELL_X2 FILLER_163_1261 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X32 FILLER_163_1584 ();
 FILLCELL_X32 FILLER_163_1616 ();
 FILLCELL_X32 FILLER_163_1648 ();
 FILLCELL_X32 FILLER_163_1680 ();
 FILLCELL_X32 FILLER_163_1712 ();
 FILLCELL_X32 FILLER_163_1744 ();
 FILLCELL_X32 FILLER_163_1776 ();
 FILLCELL_X32 FILLER_163_1808 ();
 FILLCELL_X32 FILLER_163_1840 ();
 FILLCELL_X16 FILLER_163_1872 ();
 FILLCELL_X8 FILLER_163_1888 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X32 FILLER_164_1304 ();
 FILLCELL_X32 FILLER_164_1336 ();
 FILLCELL_X32 FILLER_164_1368 ();
 FILLCELL_X32 FILLER_164_1400 ();
 FILLCELL_X32 FILLER_164_1432 ();
 FILLCELL_X32 FILLER_164_1464 ();
 FILLCELL_X32 FILLER_164_1496 ();
 FILLCELL_X32 FILLER_164_1528 ();
 FILLCELL_X32 FILLER_164_1560 ();
 FILLCELL_X32 FILLER_164_1592 ();
 FILLCELL_X32 FILLER_164_1624 ();
 FILLCELL_X32 FILLER_164_1656 ();
 FILLCELL_X32 FILLER_164_1688 ();
 FILLCELL_X32 FILLER_164_1720 ();
 FILLCELL_X32 FILLER_164_1752 ();
 FILLCELL_X32 FILLER_164_1784 ();
 FILLCELL_X32 FILLER_164_1816 ();
 FILLCELL_X32 FILLER_164_1848 ();
 FILLCELL_X8 FILLER_164_1880 ();
 FILLCELL_X4 FILLER_164_1888 ();
 FILLCELL_X2 FILLER_164_1892 ();
 FILLCELL_X1 FILLER_164_1895 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X32 FILLER_165_993 ();
 FILLCELL_X32 FILLER_165_1025 ();
 FILLCELL_X32 FILLER_165_1057 ();
 FILLCELL_X32 FILLER_165_1089 ();
 FILLCELL_X32 FILLER_165_1121 ();
 FILLCELL_X32 FILLER_165_1153 ();
 FILLCELL_X32 FILLER_165_1185 ();
 FILLCELL_X32 FILLER_165_1217 ();
 FILLCELL_X8 FILLER_165_1249 ();
 FILLCELL_X4 FILLER_165_1257 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X32 FILLER_165_1584 ();
 FILLCELL_X32 FILLER_165_1616 ();
 FILLCELL_X32 FILLER_165_1648 ();
 FILLCELL_X32 FILLER_165_1680 ();
 FILLCELL_X32 FILLER_165_1712 ();
 FILLCELL_X32 FILLER_165_1744 ();
 FILLCELL_X32 FILLER_165_1776 ();
 FILLCELL_X32 FILLER_165_1808 ();
 FILLCELL_X32 FILLER_165_1840 ();
 FILLCELL_X16 FILLER_165_1872 ();
 FILLCELL_X8 FILLER_165_1888 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X32 FILLER_166_1048 ();
 FILLCELL_X32 FILLER_166_1080 ();
 FILLCELL_X32 FILLER_166_1112 ();
 FILLCELL_X32 FILLER_166_1144 ();
 FILLCELL_X32 FILLER_166_1176 ();
 FILLCELL_X32 FILLER_166_1208 ();
 FILLCELL_X32 FILLER_166_1240 ();
 FILLCELL_X32 FILLER_166_1272 ();
 FILLCELL_X32 FILLER_166_1304 ();
 FILLCELL_X32 FILLER_166_1336 ();
 FILLCELL_X32 FILLER_166_1368 ();
 FILLCELL_X32 FILLER_166_1400 ();
 FILLCELL_X32 FILLER_166_1432 ();
 FILLCELL_X32 FILLER_166_1464 ();
 FILLCELL_X32 FILLER_166_1496 ();
 FILLCELL_X32 FILLER_166_1528 ();
 FILLCELL_X32 FILLER_166_1560 ();
 FILLCELL_X32 FILLER_166_1592 ();
 FILLCELL_X32 FILLER_166_1624 ();
 FILLCELL_X32 FILLER_166_1656 ();
 FILLCELL_X32 FILLER_166_1688 ();
 FILLCELL_X32 FILLER_166_1720 ();
 FILLCELL_X32 FILLER_166_1752 ();
 FILLCELL_X32 FILLER_166_1784 ();
 FILLCELL_X32 FILLER_166_1816 ();
 FILLCELL_X32 FILLER_166_1848 ();
 FILLCELL_X8 FILLER_166_1880 ();
 FILLCELL_X4 FILLER_166_1888 ();
 FILLCELL_X2 FILLER_166_1892 ();
 FILLCELL_X1 FILLER_166_1895 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X32 FILLER_167_801 ();
 FILLCELL_X32 FILLER_167_833 ();
 FILLCELL_X32 FILLER_167_865 ();
 FILLCELL_X32 FILLER_167_897 ();
 FILLCELL_X32 FILLER_167_929 ();
 FILLCELL_X32 FILLER_167_961 ();
 FILLCELL_X32 FILLER_167_993 ();
 FILLCELL_X32 FILLER_167_1025 ();
 FILLCELL_X32 FILLER_167_1057 ();
 FILLCELL_X32 FILLER_167_1089 ();
 FILLCELL_X32 FILLER_167_1121 ();
 FILLCELL_X32 FILLER_167_1153 ();
 FILLCELL_X32 FILLER_167_1185 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X8 FILLER_167_1249 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X32 FILLER_167_1584 ();
 FILLCELL_X32 FILLER_167_1616 ();
 FILLCELL_X32 FILLER_167_1648 ();
 FILLCELL_X32 FILLER_167_1680 ();
 FILLCELL_X32 FILLER_167_1712 ();
 FILLCELL_X32 FILLER_167_1744 ();
 FILLCELL_X32 FILLER_167_1776 ();
 FILLCELL_X32 FILLER_167_1808 ();
 FILLCELL_X32 FILLER_167_1840 ();
 FILLCELL_X16 FILLER_167_1872 ();
 FILLCELL_X8 FILLER_167_1888 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X32 FILLER_168_1176 ();
 FILLCELL_X32 FILLER_168_1208 ();
 FILLCELL_X32 FILLER_168_1240 ();
 FILLCELL_X32 FILLER_168_1272 ();
 FILLCELL_X32 FILLER_168_1304 ();
 FILLCELL_X32 FILLER_168_1336 ();
 FILLCELL_X32 FILLER_168_1368 ();
 FILLCELL_X32 FILLER_168_1400 ();
 FILLCELL_X32 FILLER_168_1432 ();
 FILLCELL_X32 FILLER_168_1464 ();
 FILLCELL_X32 FILLER_168_1496 ();
 FILLCELL_X32 FILLER_168_1528 ();
 FILLCELL_X32 FILLER_168_1560 ();
 FILLCELL_X32 FILLER_168_1592 ();
 FILLCELL_X32 FILLER_168_1624 ();
 FILLCELL_X32 FILLER_168_1656 ();
 FILLCELL_X32 FILLER_168_1688 ();
 FILLCELL_X32 FILLER_168_1720 ();
 FILLCELL_X32 FILLER_168_1752 ();
 FILLCELL_X32 FILLER_168_1784 ();
 FILLCELL_X32 FILLER_168_1816 ();
 FILLCELL_X32 FILLER_168_1848 ();
 FILLCELL_X8 FILLER_168_1880 ();
 FILLCELL_X4 FILLER_168_1888 ();
 FILLCELL_X2 FILLER_168_1892 ();
 FILLCELL_X1 FILLER_168_1895 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X32 FILLER_169_577 ();
 FILLCELL_X32 FILLER_169_609 ();
 FILLCELL_X32 FILLER_169_641 ();
 FILLCELL_X32 FILLER_169_673 ();
 FILLCELL_X32 FILLER_169_705 ();
 FILLCELL_X32 FILLER_169_737 ();
 FILLCELL_X32 FILLER_169_769 ();
 FILLCELL_X32 FILLER_169_801 ();
 FILLCELL_X32 FILLER_169_833 ();
 FILLCELL_X32 FILLER_169_865 ();
 FILLCELL_X32 FILLER_169_897 ();
 FILLCELL_X32 FILLER_169_929 ();
 FILLCELL_X32 FILLER_169_961 ();
 FILLCELL_X32 FILLER_169_993 ();
 FILLCELL_X32 FILLER_169_1025 ();
 FILLCELL_X32 FILLER_169_1057 ();
 FILLCELL_X32 FILLER_169_1089 ();
 FILLCELL_X32 FILLER_169_1121 ();
 FILLCELL_X32 FILLER_169_1153 ();
 FILLCELL_X32 FILLER_169_1185 ();
 FILLCELL_X32 FILLER_169_1217 ();
 FILLCELL_X8 FILLER_169_1249 ();
 FILLCELL_X4 FILLER_169_1257 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X32 FILLER_169_1584 ();
 FILLCELL_X32 FILLER_169_1616 ();
 FILLCELL_X32 FILLER_169_1648 ();
 FILLCELL_X32 FILLER_169_1680 ();
 FILLCELL_X32 FILLER_169_1712 ();
 FILLCELL_X32 FILLER_169_1744 ();
 FILLCELL_X32 FILLER_169_1776 ();
 FILLCELL_X32 FILLER_169_1808 ();
 FILLCELL_X32 FILLER_169_1840 ();
 FILLCELL_X16 FILLER_169_1872 ();
 FILLCELL_X8 FILLER_169_1888 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X32 FILLER_170_1048 ();
 FILLCELL_X32 FILLER_170_1080 ();
 FILLCELL_X32 FILLER_170_1112 ();
 FILLCELL_X32 FILLER_170_1144 ();
 FILLCELL_X32 FILLER_170_1176 ();
 FILLCELL_X32 FILLER_170_1208 ();
 FILLCELL_X32 FILLER_170_1240 ();
 FILLCELL_X32 FILLER_170_1272 ();
 FILLCELL_X32 FILLER_170_1304 ();
 FILLCELL_X32 FILLER_170_1336 ();
 FILLCELL_X32 FILLER_170_1368 ();
 FILLCELL_X32 FILLER_170_1400 ();
 FILLCELL_X32 FILLER_170_1432 ();
 FILLCELL_X32 FILLER_170_1464 ();
 FILLCELL_X32 FILLER_170_1496 ();
 FILLCELL_X32 FILLER_170_1528 ();
 FILLCELL_X32 FILLER_170_1560 ();
 FILLCELL_X32 FILLER_170_1592 ();
 FILLCELL_X32 FILLER_170_1624 ();
 FILLCELL_X32 FILLER_170_1656 ();
 FILLCELL_X32 FILLER_170_1688 ();
 FILLCELL_X32 FILLER_170_1720 ();
 FILLCELL_X32 FILLER_170_1752 ();
 FILLCELL_X32 FILLER_170_1784 ();
 FILLCELL_X32 FILLER_170_1816 ();
 FILLCELL_X32 FILLER_170_1848 ();
 FILLCELL_X8 FILLER_170_1880 ();
 FILLCELL_X4 FILLER_170_1888 ();
 FILLCELL_X2 FILLER_170_1892 ();
 FILLCELL_X1 FILLER_170_1895 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X32 FILLER_171_353 ();
 FILLCELL_X32 FILLER_171_385 ();
 FILLCELL_X32 FILLER_171_417 ();
 FILLCELL_X32 FILLER_171_449 ();
 FILLCELL_X32 FILLER_171_481 ();
 FILLCELL_X32 FILLER_171_513 ();
 FILLCELL_X32 FILLER_171_545 ();
 FILLCELL_X32 FILLER_171_577 ();
 FILLCELL_X32 FILLER_171_609 ();
 FILLCELL_X32 FILLER_171_641 ();
 FILLCELL_X32 FILLER_171_673 ();
 FILLCELL_X32 FILLER_171_705 ();
 FILLCELL_X32 FILLER_171_737 ();
 FILLCELL_X32 FILLER_171_769 ();
 FILLCELL_X32 FILLER_171_801 ();
 FILLCELL_X32 FILLER_171_833 ();
 FILLCELL_X32 FILLER_171_865 ();
 FILLCELL_X32 FILLER_171_897 ();
 FILLCELL_X32 FILLER_171_929 ();
 FILLCELL_X32 FILLER_171_961 ();
 FILLCELL_X32 FILLER_171_993 ();
 FILLCELL_X32 FILLER_171_1025 ();
 FILLCELL_X32 FILLER_171_1057 ();
 FILLCELL_X32 FILLER_171_1089 ();
 FILLCELL_X32 FILLER_171_1121 ();
 FILLCELL_X32 FILLER_171_1153 ();
 FILLCELL_X32 FILLER_171_1185 ();
 FILLCELL_X32 FILLER_171_1217 ();
 FILLCELL_X8 FILLER_171_1249 ();
 FILLCELL_X4 FILLER_171_1257 ();
 FILLCELL_X2 FILLER_171_1261 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X32 FILLER_171_1584 ();
 FILLCELL_X32 FILLER_171_1616 ();
 FILLCELL_X32 FILLER_171_1648 ();
 FILLCELL_X32 FILLER_171_1680 ();
 FILLCELL_X32 FILLER_171_1712 ();
 FILLCELL_X32 FILLER_171_1744 ();
 FILLCELL_X32 FILLER_171_1776 ();
 FILLCELL_X32 FILLER_171_1808 ();
 FILLCELL_X32 FILLER_171_1840 ();
 FILLCELL_X16 FILLER_171_1872 ();
 FILLCELL_X8 FILLER_171_1888 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X32 FILLER_172_1080 ();
 FILLCELL_X32 FILLER_172_1112 ();
 FILLCELL_X32 FILLER_172_1144 ();
 FILLCELL_X32 FILLER_172_1176 ();
 FILLCELL_X32 FILLER_172_1208 ();
 FILLCELL_X32 FILLER_172_1240 ();
 FILLCELL_X32 FILLER_172_1272 ();
 FILLCELL_X32 FILLER_172_1304 ();
 FILLCELL_X32 FILLER_172_1336 ();
 FILLCELL_X32 FILLER_172_1368 ();
 FILLCELL_X32 FILLER_172_1400 ();
 FILLCELL_X32 FILLER_172_1432 ();
 FILLCELL_X32 FILLER_172_1464 ();
 FILLCELL_X32 FILLER_172_1496 ();
 FILLCELL_X32 FILLER_172_1528 ();
 FILLCELL_X32 FILLER_172_1560 ();
 FILLCELL_X32 FILLER_172_1592 ();
 FILLCELL_X32 FILLER_172_1624 ();
 FILLCELL_X32 FILLER_172_1656 ();
 FILLCELL_X32 FILLER_172_1688 ();
 FILLCELL_X32 FILLER_172_1720 ();
 FILLCELL_X32 FILLER_172_1752 ();
 FILLCELL_X32 FILLER_172_1784 ();
 FILLCELL_X32 FILLER_172_1816 ();
 FILLCELL_X32 FILLER_172_1848 ();
 FILLCELL_X8 FILLER_172_1880 ();
 FILLCELL_X4 FILLER_172_1888 ();
 FILLCELL_X2 FILLER_172_1892 ();
 FILLCELL_X1 FILLER_172_1895 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X32 FILLER_173_1089 ();
 FILLCELL_X32 FILLER_173_1121 ();
 FILLCELL_X32 FILLER_173_1153 ();
 FILLCELL_X32 FILLER_173_1185 ();
 FILLCELL_X32 FILLER_173_1217 ();
 FILLCELL_X8 FILLER_173_1249 ();
 FILLCELL_X4 FILLER_173_1257 ();
 FILLCELL_X2 FILLER_173_1261 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X32 FILLER_173_1584 ();
 FILLCELL_X32 FILLER_173_1616 ();
 FILLCELL_X32 FILLER_173_1648 ();
 FILLCELL_X32 FILLER_173_1680 ();
 FILLCELL_X32 FILLER_173_1712 ();
 FILLCELL_X32 FILLER_173_1744 ();
 FILLCELL_X32 FILLER_173_1776 ();
 FILLCELL_X32 FILLER_173_1808 ();
 FILLCELL_X32 FILLER_173_1840 ();
 FILLCELL_X16 FILLER_173_1872 ();
 FILLCELL_X8 FILLER_173_1888 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X32 FILLER_174_1304 ();
 FILLCELL_X32 FILLER_174_1336 ();
 FILLCELL_X32 FILLER_174_1368 ();
 FILLCELL_X32 FILLER_174_1400 ();
 FILLCELL_X32 FILLER_174_1432 ();
 FILLCELL_X32 FILLER_174_1464 ();
 FILLCELL_X32 FILLER_174_1496 ();
 FILLCELL_X32 FILLER_174_1528 ();
 FILLCELL_X32 FILLER_174_1560 ();
 FILLCELL_X32 FILLER_174_1592 ();
 FILLCELL_X32 FILLER_174_1624 ();
 FILLCELL_X32 FILLER_174_1656 ();
 FILLCELL_X32 FILLER_174_1688 ();
 FILLCELL_X32 FILLER_174_1720 ();
 FILLCELL_X32 FILLER_174_1752 ();
 FILLCELL_X32 FILLER_174_1784 ();
 FILLCELL_X32 FILLER_174_1816 ();
 FILLCELL_X32 FILLER_174_1848 ();
 FILLCELL_X8 FILLER_174_1880 ();
 FILLCELL_X4 FILLER_174_1888 ();
 FILLCELL_X2 FILLER_174_1892 ();
 FILLCELL_X1 FILLER_174_1895 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X32 FILLER_175_385 ();
 FILLCELL_X32 FILLER_175_417 ();
 FILLCELL_X32 FILLER_175_449 ();
 FILLCELL_X32 FILLER_175_481 ();
 FILLCELL_X32 FILLER_175_513 ();
 FILLCELL_X32 FILLER_175_545 ();
 FILLCELL_X32 FILLER_175_577 ();
 FILLCELL_X32 FILLER_175_609 ();
 FILLCELL_X32 FILLER_175_641 ();
 FILLCELL_X32 FILLER_175_673 ();
 FILLCELL_X32 FILLER_175_705 ();
 FILLCELL_X32 FILLER_175_737 ();
 FILLCELL_X32 FILLER_175_769 ();
 FILLCELL_X32 FILLER_175_801 ();
 FILLCELL_X32 FILLER_175_833 ();
 FILLCELL_X32 FILLER_175_865 ();
 FILLCELL_X32 FILLER_175_897 ();
 FILLCELL_X32 FILLER_175_929 ();
 FILLCELL_X32 FILLER_175_961 ();
 FILLCELL_X32 FILLER_175_993 ();
 FILLCELL_X32 FILLER_175_1025 ();
 FILLCELL_X32 FILLER_175_1057 ();
 FILLCELL_X32 FILLER_175_1089 ();
 FILLCELL_X32 FILLER_175_1121 ();
 FILLCELL_X32 FILLER_175_1153 ();
 FILLCELL_X32 FILLER_175_1185 ();
 FILLCELL_X32 FILLER_175_1217 ();
 FILLCELL_X8 FILLER_175_1249 ();
 FILLCELL_X4 FILLER_175_1257 ();
 FILLCELL_X2 FILLER_175_1261 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X32 FILLER_175_1584 ();
 FILLCELL_X32 FILLER_175_1616 ();
 FILLCELL_X32 FILLER_175_1648 ();
 FILLCELL_X32 FILLER_175_1680 ();
 FILLCELL_X32 FILLER_175_1712 ();
 FILLCELL_X32 FILLER_175_1744 ();
 FILLCELL_X32 FILLER_175_1776 ();
 FILLCELL_X32 FILLER_175_1808 ();
 FILLCELL_X32 FILLER_175_1840 ();
 FILLCELL_X16 FILLER_175_1872 ();
 FILLCELL_X8 FILLER_175_1888 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X32 FILLER_176_353 ();
 FILLCELL_X32 FILLER_176_385 ();
 FILLCELL_X32 FILLER_176_417 ();
 FILLCELL_X32 FILLER_176_449 ();
 FILLCELL_X32 FILLER_176_481 ();
 FILLCELL_X32 FILLER_176_513 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X32 FILLER_176_577 ();
 FILLCELL_X16 FILLER_176_609 ();
 FILLCELL_X4 FILLER_176_625 ();
 FILLCELL_X2 FILLER_176_629 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X32 FILLER_176_1112 ();
 FILLCELL_X32 FILLER_176_1144 ();
 FILLCELL_X32 FILLER_176_1176 ();
 FILLCELL_X32 FILLER_176_1208 ();
 FILLCELL_X32 FILLER_176_1240 ();
 FILLCELL_X32 FILLER_176_1272 ();
 FILLCELL_X32 FILLER_176_1304 ();
 FILLCELL_X32 FILLER_176_1336 ();
 FILLCELL_X32 FILLER_176_1368 ();
 FILLCELL_X32 FILLER_176_1400 ();
 FILLCELL_X32 FILLER_176_1432 ();
 FILLCELL_X32 FILLER_176_1464 ();
 FILLCELL_X32 FILLER_176_1496 ();
 FILLCELL_X32 FILLER_176_1528 ();
 FILLCELL_X32 FILLER_176_1560 ();
 FILLCELL_X32 FILLER_176_1592 ();
 FILLCELL_X32 FILLER_176_1624 ();
 FILLCELL_X32 FILLER_176_1656 ();
 FILLCELL_X32 FILLER_176_1688 ();
 FILLCELL_X32 FILLER_176_1720 ();
 FILLCELL_X32 FILLER_176_1752 ();
 FILLCELL_X32 FILLER_176_1784 ();
 FILLCELL_X32 FILLER_176_1816 ();
 FILLCELL_X32 FILLER_176_1848 ();
 FILLCELL_X8 FILLER_176_1880 ();
 FILLCELL_X4 FILLER_176_1888 ();
 FILLCELL_X2 FILLER_176_1892 ();
 FILLCELL_X1 FILLER_176_1895 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X32 FILLER_177_1089 ();
 FILLCELL_X32 FILLER_177_1121 ();
 FILLCELL_X32 FILLER_177_1153 ();
 FILLCELL_X32 FILLER_177_1185 ();
 FILLCELL_X32 FILLER_177_1217 ();
 FILLCELL_X8 FILLER_177_1249 ();
 FILLCELL_X4 FILLER_177_1257 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X32 FILLER_177_1584 ();
 FILLCELL_X32 FILLER_177_1616 ();
 FILLCELL_X32 FILLER_177_1648 ();
 FILLCELL_X32 FILLER_177_1680 ();
 FILLCELL_X32 FILLER_177_1712 ();
 FILLCELL_X32 FILLER_177_1744 ();
 FILLCELL_X32 FILLER_177_1776 ();
 FILLCELL_X32 FILLER_177_1808 ();
 FILLCELL_X32 FILLER_177_1840 ();
 FILLCELL_X16 FILLER_177_1872 ();
 FILLCELL_X8 FILLER_177_1888 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X32 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1144 ();
 FILLCELL_X32 FILLER_178_1176 ();
 FILLCELL_X32 FILLER_178_1208 ();
 FILLCELL_X32 FILLER_178_1240 ();
 FILLCELL_X32 FILLER_178_1272 ();
 FILLCELL_X32 FILLER_178_1304 ();
 FILLCELL_X32 FILLER_178_1336 ();
 FILLCELL_X32 FILLER_178_1368 ();
 FILLCELL_X32 FILLER_178_1400 ();
 FILLCELL_X32 FILLER_178_1432 ();
 FILLCELL_X32 FILLER_178_1464 ();
 FILLCELL_X32 FILLER_178_1496 ();
 FILLCELL_X32 FILLER_178_1528 ();
 FILLCELL_X32 FILLER_178_1560 ();
 FILLCELL_X32 FILLER_178_1592 ();
 FILLCELL_X32 FILLER_178_1624 ();
 FILLCELL_X32 FILLER_178_1656 ();
 FILLCELL_X32 FILLER_178_1688 ();
 FILLCELL_X32 FILLER_178_1720 ();
 FILLCELL_X32 FILLER_178_1752 ();
 FILLCELL_X32 FILLER_178_1784 ();
 FILLCELL_X32 FILLER_178_1816 ();
 FILLCELL_X32 FILLER_178_1848 ();
 FILLCELL_X8 FILLER_178_1880 ();
 FILLCELL_X4 FILLER_178_1888 ();
 FILLCELL_X2 FILLER_178_1892 ();
 FILLCELL_X1 FILLER_178_1895 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X32 FILLER_179_1089 ();
 FILLCELL_X32 FILLER_179_1121 ();
 FILLCELL_X32 FILLER_179_1153 ();
 FILLCELL_X32 FILLER_179_1185 ();
 FILLCELL_X32 FILLER_179_1217 ();
 FILLCELL_X8 FILLER_179_1249 ();
 FILLCELL_X4 FILLER_179_1257 ();
 FILLCELL_X2 FILLER_179_1261 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X32 FILLER_179_1584 ();
 FILLCELL_X32 FILLER_179_1616 ();
 FILLCELL_X32 FILLER_179_1648 ();
 FILLCELL_X32 FILLER_179_1680 ();
 FILLCELL_X32 FILLER_179_1712 ();
 FILLCELL_X32 FILLER_179_1744 ();
 FILLCELL_X32 FILLER_179_1776 ();
 FILLCELL_X32 FILLER_179_1808 ();
 FILLCELL_X32 FILLER_179_1840 ();
 FILLCELL_X16 FILLER_179_1872 ();
 FILLCELL_X8 FILLER_179_1888 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X32 FILLER_180_353 ();
 FILLCELL_X32 FILLER_180_385 ();
 FILLCELL_X32 FILLER_180_417 ();
 FILLCELL_X32 FILLER_180_449 ();
 FILLCELL_X32 FILLER_180_481 ();
 FILLCELL_X32 FILLER_180_513 ();
 FILLCELL_X32 FILLER_180_545 ();
 FILLCELL_X32 FILLER_180_577 ();
 FILLCELL_X16 FILLER_180_609 ();
 FILLCELL_X4 FILLER_180_625 ();
 FILLCELL_X2 FILLER_180_629 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X32 FILLER_180_1080 ();
 FILLCELL_X32 FILLER_180_1112 ();
 FILLCELL_X32 FILLER_180_1144 ();
 FILLCELL_X32 FILLER_180_1176 ();
 FILLCELL_X32 FILLER_180_1208 ();
 FILLCELL_X32 FILLER_180_1240 ();
 FILLCELL_X32 FILLER_180_1272 ();
 FILLCELL_X32 FILLER_180_1304 ();
 FILLCELL_X32 FILLER_180_1336 ();
 FILLCELL_X32 FILLER_180_1368 ();
 FILLCELL_X32 FILLER_180_1400 ();
 FILLCELL_X32 FILLER_180_1432 ();
 FILLCELL_X32 FILLER_180_1464 ();
 FILLCELL_X32 FILLER_180_1496 ();
 FILLCELL_X32 FILLER_180_1528 ();
 FILLCELL_X32 FILLER_180_1560 ();
 FILLCELL_X32 FILLER_180_1592 ();
 FILLCELL_X32 FILLER_180_1624 ();
 FILLCELL_X32 FILLER_180_1656 ();
 FILLCELL_X32 FILLER_180_1688 ();
 FILLCELL_X32 FILLER_180_1720 ();
 FILLCELL_X32 FILLER_180_1752 ();
 FILLCELL_X32 FILLER_180_1784 ();
 FILLCELL_X32 FILLER_180_1816 ();
 FILLCELL_X32 FILLER_180_1848 ();
 FILLCELL_X8 FILLER_180_1880 ();
 FILLCELL_X4 FILLER_180_1888 ();
 FILLCELL_X2 FILLER_180_1892 ();
 FILLCELL_X1 FILLER_180_1895 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X32 FILLER_181_1089 ();
 FILLCELL_X32 FILLER_181_1121 ();
 FILLCELL_X32 FILLER_181_1153 ();
 FILLCELL_X32 FILLER_181_1185 ();
 FILLCELL_X32 FILLER_181_1217 ();
 FILLCELL_X8 FILLER_181_1249 ();
 FILLCELL_X4 FILLER_181_1257 ();
 FILLCELL_X2 FILLER_181_1261 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X32 FILLER_181_1584 ();
 FILLCELL_X32 FILLER_181_1616 ();
 FILLCELL_X32 FILLER_181_1648 ();
 FILLCELL_X32 FILLER_181_1680 ();
 FILLCELL_X32 FILLER_181_1712 ();
 FILLCELL_X32 FILLER_181_1744 ();
 FILLCELL_X32 FILLER_181_1776 ();
 FILLCELL_X32 FILLER_181_1808 ();
 FILLCELL_X32 FILLER_181_1840 ();
 FILLCELL_X16 FILLER_181_1872 ();
 FILLCELL_X8 FILLER_181_1888 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X32 FILLER_182_1080 ();
 FILLCELL_X32 FILLER_182_1112 ();
 FILLCELL_X32 FILLER_182_1144 ();
 FILLCELL_X32 FILLER_182_1176 ();
 FILLCELL_X32 FILLER_182_1208 ();
 FILLCELL_X32 FILLER_182_1240 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X32 FILLER_182_1400 ();
 FILLCELL_X32 FILLER_182_1432 ();
 FILLCELL_X32 FILLER_182_1464 ();
 FILLCELL_X32 FILLER_182_1496 ();
 FILLCELL_X32 FILLER_182_1528 ();
 FILLCELL_X32 FILLER_182_1560 ();
 FILLCELL_X32 FILLER_182_1592 ();
 FILLCELL_X32 FILLER_182_1624 ();
 FILLCELL_X32 FILLER_182_1656 ();
 FILLCELL_X32 FILLER_182_1688 ();
 FILLCELL_X32 FILLER_182_1720 ();
 FILLCELL_X32 FILLER_182_1752 ();
 FILLCELL_X32 FILLER_182_1784 ();
 FILLCELL_X32 FILLER_182_1816 ();
 FILLCELL_X32 FILLER_182_1848 ();
 FILLCELL_X8 FILLER_182_1880 ();
 FILLCELL_X4 FILLER_182_1888 ();
 FILLCELL_X2 FILLER_182_1892 ();
 FILLCELL_X1 FILLER_182_1895 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X32 FILLER_183_1089 ();
 FILLCELL_X32 FILLER_183_1121 ();
 FILLCELL_X32 FILLER_183_1153 ();
 FILLCELL_X32 FILLER_183_1185 ();
 FILLCELL_X32 FILLER_183_1217 ();
 FILLCELL_X8 FILLER_183_1249 ();
 FILLCELL_X4 FILLER_183_1257 ();
 FILLCELL_X2 FILLER_183_1261 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X32 FILLER_183_1584 ();
 FILLCELL_X32 FILLER_183_1616 ();
 FILLCELL_X32 FILLER_183_1648 ();
 FILLCELL_X32 FILLER_183_1680 ();
 FILLCELL_X32 FILLER_183_1712 ();
 FILLCELL_X32 FILLER_183_1744 ();
 FILLCELL_X32 FILLER_183_1776 ();
 FILLCELL_X32 FILLER_183_1808 ();
 FILLCELL_X32 FILLER_183_1840 ();
 FILLCELL_X16 FILLER_183_1872 ();
 FILLCELL_X8 FILLER_183_1888 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X32 FILLER_184_1144 ();
 FILLCELL_X32 FILLER_184_1176 ();
 FILLCELL_X32 FILLER_184_1208 ();
 FILLCELL_X32 FILLER_184_1240 ();
 FILLCELL_X32 FILLER_184_1272 ();
 FILLCELL_X32 FILLER_184_1304 ();
 FILLCELL_X32 FILLER_184_1336 ();
 FILLCELL_X32 FILLER_184_1368 ();
 FILLCELL_X32 FILLER_184_1400 ();
 FILLCELL_X32 FILLER_184_1432 ();
 FILLCELL_X32 FILLER_184_1464 ();
 FILLCELL_X32 FILLER_184_1496 ();
 FILLCELL_X32 FILLER_184_1528 ();
 FILLCELL_X32 FILLER_184_1560 ();
 FILLCELL_X32 FILLER_184_1592 ();
 FILLCELL_X32 FILLER_184_1624 ();
 FILLCELL_X32 FILLER_184_1656 ();
 FILLCELL_X32 FILLER_184_1688 ();
 FILLCELL_X32 FILLER_184_1720 ();
 FILLCELL_X32 FILLER_184_1752 ();
 FILLCELL_X32 FILLER_184_1784 ();
 FILLCELL_X32 FILLER_184_1816 ();
 FILLCELL_X32 FILLER_184_1848 ();
 FILLCELL_X8 FILLER_184_1880 ();
 FILLCELL_X4 FILLER_184_1888 ();
 FILLCELL_X2 FILLER_184_1892 ();
 FILLCELL_X1 FILLER_184_1895 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X32 FILLER_185_1185 ();
 FILLCELL_X32 FILLER_185_1217 ();
 FILLCELL_X8 FILLER_185_1249 ();
 FILLCELL_X4 FILLER_185_1257 ();
 FILLCELL_X2 FILLER_185_1261 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X32 FILLER_185_1584 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X32 FILLER_185_1648 ();
 FILLCELL_X32 FILLER_185_1680 ();
 FILLCELL_X32 FILLER_185_1712 ();
 FILLCELL_X32 FILLER_185_1744 ();
 FILLCELL_X32 FILLER_185_1776 ();
 FILLCELL_X32 FILLER_185_1808 ();
 FILLCELL_X32 FILLER_185_1840 ();
 FILLCELL_X16 FILLER_185_1872 ();
 FILLCELL_X8 FILLER_185_1888 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X32 FILLER_186_1240 ();
 FILLCELL_X32 FILLER_186_1272 ();
 FILLCELL_X32 FILLER_186_1304 ();
 FILLCELL_X32 FILLER_186_1336 ();
 FILLCELL_X32 FILLER_186_1368 ();
 FILLCELL_X32 FILLER_186_1400 ();
 FILLCELL_X32 FILLER_186_1432 ();
 FILLCELL_X32 FILLER_186_1464 ();
 FILLCELL_X32 FILLER_186_1496 ();
 FILLCELL_X32 FILLER_186_1528 ();
 FILLCELL_X32 FILLER_186_1560 ();
 FILLCELL_X32 FILLER_186_1592 ();
 FILLCELL_X32 FILLER_186_1624 ();
 FILLCELL_X32 FILLER_186_1656 ();
 FILLCELL_X32 FILLER_186_1688 ();
 FILLCELL_X32 FILLER_186_1720 ();
 FILLCELL_X32 FILLER_186_1752 ();
 FILLCELL_X32 FILLER_186_1784 ();
 FILLCELL_X32 FILLER_186_1816 ();
 FILLCELL_X32 FILLER_186_1848 ();
 FILLCELL_X8 FILLER_186_1880 ();
 FILLCELL_X4 FILLER_186_1888 ();
 FILLCELL_X2 FILLER_186_1892 ();
 FILLCELL_X1 FILLER_186_1895 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X32 FILLER_187_1217 ();
 FILLCELL_X8 FILLER_187_1249 ();
 FILLCELL_X4 FILLER_187_1257 ();
 FILLCELL_X2 FILLER_187_1261 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X32 FILLER_187_1584 ();
 FILLCELL_X32 FILLER_187_1616 ();
 FILLCELL_X32 FILLER_187_1648 ();
 FILLCELL_X32 FILLER_187_1680 ();
 FILLCELL_X32 FILLER_187_1712 ();
 FILLCELL_X32 FILLER_187_1744 ();
 FILLCELL_X32 FILLER_187_1776 ();
 FILLCELL_X32 FILLER_187_1808 ();
 FILLCELL_X32 FILLER_187_1840 ();
 FILLCELL_X16 FILLER_187_1872 ();
 FILLCELL_X8 FILLER_187_1888 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X32 FILLER_188_1240 ();
 FILLCELL_X32 FILLER_188_1272 ();
 FILLCELL_X32 FILLER_188_1304 ();
 FILLCELL_X32 FILLER_188_1336 ();
 FILLCELL_X32 FILLER_188_1368 ();
 FILLCELL_X32 FILLER_188_1400 ();
 FILLCELL_X32 FILLER_188_1432 ();
 FILLCELL_X32 FILLER_188_1464 ();
 FILLCELL_X32 FILLER_188_1496 ();
 FILLCELL_X32 FILLER_188_1528 ();
 FILLCELL_X32 FILLER_188_1560 ();
 FILLCELL_X32 FILLER_188_1592 ();
 FILLCELL_X32 FILLER_188_1624 ();
 FILLCELL_X32 FILLER_188_1656 ();
 FILLCELL_X32 FILLER_188_1688 ();
 FILLCELL_X32 FILLER_188_1720 ();
 FILLCELL_X32 FILLER_188_1752 ();
 FILLCELL_X32 FILLER_188_1784 ();
 FILLCELL_X32 FILLER_188_1816 ();
 FILLCELL_X32 FILLER_188_1848 ();
 FILLCELL_X8 FILLER_188_1880 ();
 FILLCELL_X4 FILLER_188_1888 ();
 FILLCELL_X2 FILLER_188_1892 ();
 FILLCELL_X1 FILLER_188_1895 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X8 FILLER_189_1249 ();
 FILLCELL_X4 FILLER_189_1257 ();
 FILLCELL_X2 FILLER_189_1261 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X32 FILLER_189_1584 ();
 FILLCELL_X32 FILLER_189_1616 ();
 FILLCELL_X32 FILLER_189_1648 ();
 FILLCELL_X32 FILLER_189_1680 ();
 FILLCELL_X32 FILLER_189_1712 ();
 FILLCELL_X32 FILLER_189_1744 ();
 FILLCELL_X32 FILLER_189_1776 ();
 FILLCELL_X32 FILLER_189_1808 ();
 FILLCELL_X32 FILLER_189_1840 ();
 FILLCELL_X16 FILLER_189_1872 ();
 FILLCELL_X8 FILLER_189_1888 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X32 FILLER_190_1240 ();
 FILLCELL_X32 FILLER_190_1272 ();
 FILLCELL_X32 FILLER_190_1304 ();
 FILLCELL_X32 FILLER_190_1336 ();
 FILLCELL_X32 FILLER_190_1368 ();
 FILLCELL_X32 FILLER_190_1400 ();
 FILLCELL_X32 FILLER_190_1432 ();
 FILLCELL_X32 FILLER_190_1464 ();
 FILLCELL_X32 FILLER_190_1496 ();
 FILLCELL_X32 FILLER_190_1528 ();
 FILLCELL_X32 FILLER_190_1560 ();
 FILLCELL_X32 FILLER_190_1592 ();
 FILLCELL_X32 FILLER_190_1624 ();
 FILLCELL_X32 FILLER_190_1656 ();
 FILLCELL_X32 FILLER_190_1688 ();
 FILLCELL_X32 FILLER_190_1720 ();
 FILLCELL_X32 FILLER_190_1752 ();
 FILLCELL_X32 FILLER_190_1784 ();
 FILLCELL_X32 FILLER_190_1816 ();
 FILLCELL_X32 FILLER_190_1848 ();
 FILLCELL_X8 FILLER_190_1880 ();
 FILLCELL_X4 FILLER_190_1888 ();
 FILLCELL_X2 FILLER_190_1892 ();
 FILLCELL_X1 FILLER_190_1895 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X32 FILLER_191_1217 ();
 FILLCELL_X8 FILLER_191_1249 ();
 FILLCELL_X4 FILLER_191_1257 ();
 FILLCELL_X2 FILLER_191_1261 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X32 FILLER_191_1584 ();
 FILLCELL_X32 FILLER_191_1616 ();
 FILLCELL_X32 FILLER_191_1648 ();
 FILLCELL_X32 FILLER_191_1680 ();
 FILLCELL_X32 FILLER_191_1712 ();
 FILLCELL_X32 FILLER_191_1744 ();
 FILLCELL_X32 FILLER_191_1776 ();
 FILLCELL_X32 FILLER_191_1808 ();
 FILLCELL_X32 FILLER_191_1840 ();
 FILLCELL_X16 FILLER_191_1872 ();
 FILLCELL_X8 FILLER_191_1888 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X32 FILLER_192_1208 ();
 FILLCELL_X32 FILLER_192_1240 ();
 FILLCELL_X32 FILLER_192_1272 ();
 FILLCELL_X32 FILLER_192_1304 ();
 FILLCELL_X32 FILLER_192_1336 ();
 FILLCELL_X32 FILLER_192_1368 ();
 FILLCELL_X32 FILLER_192_1400 ();
 FILLCELL_X32 FILLER_192_1432 ();
 FILLCELL_X32 FILLER_192_1464 ();
 FILLCELL_X32 FILLER_192_1496 ();
 FILLCELL_X32 FILLER_192_1528 ();
 FILLCELL_X32 FILLER_192_1560 ();
 FILLCELL_X32 FILLER_192_1592 ();
 FILLCELL_X32 FILLER_192_1624 ();
 FILLCELL_X32 FILLER_192_1656 ();
 FILLCELL_X32 FILLER_192_1688 ();
 FILLCELL_X32 FILLER_192_1720 ();
 FILLCELL_X32 FILLER_192_1752 ();
 FILLCELL_X32 FILLER_192_1784 ();
 FILLCELL_X32 FILLER_192_1816 ();
 FILLCELL_X32 FILLER_192_1848 ();
 FILLCELL_X8 FILLER_192_1880 ();
 FILLCELL_X4 FILLER_192_1888 ();
 FILLCELL_X2 FILLER_192_1892 ();
 FILLCELL_X1 FILLER_192_1895 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X32 FILLER_193_1584 ();
 FILLCELL_X32 FILLER_193_1616 ();
 FILLCELL_X32 FILLER_193_1648 ();
 FILLCELL_X32 FILLER_193_1680 ();
 FILLCELL_X32 FILLER_193_1712 ();
 FILLCELL_X32 FILLER_193_1744 ();
 FILLCELL_X32 FILLER_193_1776 ();
 FILLCELL_X32 FILLER_193_1808 ();
 FILLCELL_X32 FILLER_193_1840 ();
 FILLCELL_X16 FILLER_193_1872 ();
 FILLCELL_X8 FILLER_193_1888 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X32 FILLER_194_1208 ();
 FILLCELL_X32 FILLER_194_1240 ();
 FILLCELL_X32 FILLER_194_1272 ();
 FILLCELL_X32 FILLER_194_1304 ();
 FILLCELL_X32 FILLER_194_1336 ();
 FILLCELL_X32 FILLER_194_1368 ();
 FILLCELL_X32 FILLER_194_1400 ();
 FILLCELL_X32 FILLER_194_1432 ();
 FILLCELL_X32 FILLER_194_1464 ();
 FILLCELL_X32 FILLER_194_1496 ();
 FILLCELL_X32 FILLER_194_1528 ();
 FILLCELL_X32 FILLER_194_1560 ();
 FILLCELL_X32 FILLER_194_1592 ();
 FILLCELL_X32 FILLER_194_1624 ();
 FILLCELL_X32 FILLER_194_1656 ();
 FILLCELL_X32 FILLER_194_1688 ();
 FILLCELL_X32 FILLER_194_1720 ();
 FILLCELL_X32 FILLER_194_1752 ();
 FILLCELL_X32 FILLER_194_1784 ();
 FILLCELL_X32 FILLER_194_1816 ();
 FILLCELL_X32 FILLER_194_1848 ();
 FILLCELL_X8 FILLER_194_1880 ();
 FILLCELL_X4 FILLER_194_1888 ();
 FILLCELL_X2 FILLER_194_1892 ();
 FILLCELL_X1 FILLER_194_1895 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X32 FILLER_195_1217 ();
 FILLCELL_X8 FILLER_195_1249 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X32 FILLER_195_1584 ();
 FILLCELL_X32 FILLER_195_1616 ();
 FILLCELL_X32 FILLER_195_1648 ();
 FILLCELL_X32 FILLER_195_1680 ();
 FILLCELL_X32 FILLER_195_1712 ();
 FILLCELL_X32 FILLER_195_1744 ();
 FILLCELL_X32 FILLER_195_1776 ();
 FILLCELL_X32 FILLER_195_1808 ();
 FILLCELL_X32 FILLER_195_1840 ();
 FILLCELL_X16 FILLER_195_1872 ();
 FILLCELL_X8 FILLER_195_1888 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X32 FILLER_196_1272 ();
 FILLCELL_X32 FILLER_196_1304 ();
 FILLCELL_X32 FILLER_196_1336 ();
 FILLCELL_X32 FILLER_196_1368 ();
 FILLCELL_X32 FILLER_196_1400 ();
 FILLCELL_X32 FILLER_196_1432 ();
 FILLCELL_X32 FILLER_196_1464 ();
 FILLCELL_X32 FILLER_196_1496 ();
 FILLCELL_X32 FILLER_196_1528 ();
 FILLCELL_X32 FILLER_196_1560 ();
 FILLCELL_X32 FILLER_196_1592 ();
 FILLCELL_X32 FILLER_196_1624 ();
 FILLCELL_X32 FILLER_196_1656 ();
 FILLCELL_X32 FILLER_196_1688 ();
 FILLCELL_X32 FILLER_196_1720 ();
 FILLCELL_X32 FILLER_196_1752 ();
 FILLCELL_X32 FILLER_196_1784 ();
 FILLCELL_X32 FILLER_196_1816 ();
 FILLCELL_X32 FILLER_196_1848 ();
 FILLCELL_X8 FILLER_196_1880 ();
 FILLCELL_X4 FILLER_196_1888 ();
 FILLCELL_X2 FILLER_196_1892 ();
 FILLCELL_X1 FILLER_196_1895 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X32 FILLER_197_1584 ();
 FILLCELL_X32 FILLER_197_1616 ();
 FILLCELL_X32 FILLER_197_1648 ();
 FILLCELL_X32 FILLER_197_1680 ();
 FILLCELL_X32 FILLER_197_1712 ();
 FILLCELL_X32 FILLER_197_1744 ();
 FILLCELL_X32 FILLER_197_1776 ();
 FILLCELL_X32 FILLER_197_1808 ();
 FILLCELL_X32 FILLER_197_1840 ();
 FILLCELL_X16 FILLER_197_1872 ();
 FILLCELL_X8 FILLER_197_1888 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X32 FILLER_198_1208 ();
 FILLCELL_X32 FILLER_198_1240 ();
 FILLCELL_X32 FILLER_198_1272 ();
 FILLCELL_X32 FILLER_198_1304 ();
 FILLCELL_X32 FILLER_198_1336 ();
 FILLCELL_X32 FILLER_198_1368 ();
 FILLCELL_X32 FILLER_198_1400 ();
 FILLCELL_X32 FILLER_198_1432 ();
 FILLCELL_X32 FILLER_198_1464 ();
 FILLCELL_X32 FILLER_198_1496 ();
 FILLCELL_X32 FILLER_198_1528 ();
 FILLCELL_X32 FILLER_198_1560 ();
 FILLCELL_X32 FILLER_198_1592 ();
 FILLCELL_X32 FILLER_198_1624 ();
 FILLCELL_X32 FILLER_198_1656 ();
 FILLCELL_X32 FILLER_198_1688 ();
 FILLCELL_X32 FILLER_198_1720 ();
 FILLCELL_X32 FILLER_198_1752 ();
 FILLCELL_X32 FILLER_198_1784 ();
 FILLCELL_X32 FILLER_198_1816 ();
 FILLCELL_X32 FILLER_198_1848 ();
 FILLCELL_X8 FILLER_198_1880 ();
 FILLCELL_X4 FILLER_198_1888 ();
 FILLCELL_X2 FILLER_198_1892 ();
 FILLCELL_X1 FILLER_198_1895 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X32 FILLER_199_1584 ();
 FILLCELL_X32 FILLER_199_1616 ();
 FILLCELL_X32 FILLER_199_1648 ();
 FILLCELL_X32 FILLER_199_1680 ();
 FILLCELL_X32 FILLER_199_1712 ();
 FILLCELL_X32 FILLER_199_1744 ();
 FILLCELL_X32 FILLER_199_1776 ();
 FILLCELL_X32 FILLER_199_1808 ();
 FILLCELL_X32 FILLER_199_1840 ();
 FILLCELL_X16 FILLER_199_1872 ();
 FILLCELL_X8 FILLER_199_1888 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X32 FILLER_200_1304 ();
 FILLCELL_X32 FILLER_200_1336 ();
 FILLCELL_X32 FILLER_200_1368 ();
 FILLCELL_X32 FILLER_200_1400 ();
 FILLCELL_X32 FILLER_200_1432 ();
 FILLCELL_X32 FILLER_200_1464 ();
 FILLCELL_X32 FILLER_200_1496 ();
 FILLCELL_X32 FILLER_200_1528 ();
 FILLCELL_X32 FILLER_200_1560 ();
 FILLCELL_X32 FILLER_200_1592 ();
 FILLCELL_X32 FILLER_200_1624 ();
 FILLCELL_X32 FILLER_200_1656 ();
 FILLCELL_X32 FILLER_200_1688 ();
 FILLCELL_X32 FILLER_200_1720 ();
 FILLCELL_X32 FILLER_200_1752 ();
 FILLCELL_X32 FILLER_200_1784 ();
 FILLCELL_X32 FILLER_200_1816 ();
 FILLCELL_X32 FILLER_200_1848 ();
 FILLCELL_X8 FILLER_200_1880 ();
 FILLCELL_X4 FILLER_200_1888 ();
 FILLCELL_X2 FILLER_200_1892 ();
 FILLCELL_X1 FILLER_200_1895 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X32 FILLER_201_1648 ();
 FILLCELL_X32 FILLER_201_1680 ();
 FILLCELL_X32 FILLER_201_1712 ();
 FILLCELL_X32 FILLER_201_1744 ();
 FILLCELL_X32 FILLER_201_1776 ();
 FILLCELL_X32 FILLER_201_1808 ();
 FILLCELL_X32 FILLER_201_1840 ();
 FILLCELL_X16 FILLER_201_1872 ();
 FILLCELL_X8 FILLER_201_1888 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X32 FILLER_202_1592 ();
 FILLCELL_X32 FILLER_202_1624 ();
 FILLCELL_X32 FILLER_202_1656 ();
 FILLCELL_X32 FILLER_202_1688 ();
 FILLCELL_X32 FILLER_202_1720 ();
 FILLCELL_X32 FILLER_202_1752 ();
 FILLCELL_X32 FILLER_202_1784 ();
 FILLCELL_X32 FILLER_202_1816 ();
 FILLCELL_X32 FILLER_202_1848 ();
 FILLCELL_X8 FILLER_202_1880 ();
 FILLCELL_X4 FILLER_202_1888 ();
 FILLCELL_X2 FILLER_202_1892 ();
 FILLCELL_X1 FILLER_202_1895 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X32 FILLER_203_1648 ();
 FILLCELL_X32 FILLER_203_1680 ();
 FILLCELL_X32 FILLER_203_1712 ();
 FILLCELL_X32 FILLER_203_1744 ();
 FILLCELL_X32 FILLER_203_1776 ();
 FILLCELL_X32 FILLER_203_1808 ();
 FILLCELL_X32 FILLER_203_1840 ();
 FILLCELL_X16 FILLER_203_1872 ();
 FILLCELL_X8 FILLER_203_1888 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X32 FILLER_204_1592 ();
 FILLCELL_X32 FILLER_204_1624 ();
 FILLCELL_X32 FILLER_204_1656 ();
 FILLCELL_X32 FILLER_204_1688 ();
 FILLCELL_X32 FILLER_204_1720 ();
 FILLCELL_X32 FILLER_204_1752 ();
 FILLCELL_X32 FILLER_204_1784 ();
 FILLCELL_X32 FILLER_204_1816 ();
 FILLCELL_X32 FILLER_204_1848 ();
 FILLCELL_X8 FILLER_204_1880 ();
 FILLCELL_X4 FILLER_204_1888 ();
 FILLCELL_X2 FILLER_204_1892 ();
 FILLCELL_X1 FILLER_204_1895 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X32 FILLER_205_1648 ();
 FILLCELL_X32 FILLER_205_1680 ();
 FILLCELL_X32 FILLER_205_1712 ();
 FILLCELL_X32 FILLER_205_1744 ();
 FILLCELL_X32 FILLER_205_1776 ();
 FILLCELL_X32 FILLER_205_1808 ();
 FILLCELL_X32 FILLER_205_1840 ();
 FILLCELL_X16 FILLER_205_1872 ();
 FILLCELL_X8 FILLER_205_1888 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X32 FILLER_206_1592 ();
 FILLCELL_X32 FILLER_206_1624 ();
 FILLCELL_X32 FILLER_206_1656 ();
 FILLCELL_X32 FILLER_206_1688 ();
 FILLCELL_X32 FILLER_206_1720 ();
 FILLCELL_X32 FILLER_206_1752 ();
 FILLCELL_X32 FILLER_206_1784 ();
 FILLCELL_X32 FILLER_206_1816 ();
 FILLCELL_X32 FILLER_206_1848 ();
 FILLCELL_X8 FILLER_206_1880 ();
 FILLCELL_X4 FILLER_206_1888 ();
 FILLCELL_X2 FILLER_206_1892 ();
 FILLCELL_X1 FILLER_206_1895 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X32 FILLER_207_1648 ();
 FILLCELL_X32 FILLER_207_1680 ();
 FILLCELL_X32 FILLER_207_1712 ();
 FILLCELL_X32 FILLER_207_1744 ();
 FILLCELL_X32 FILLER_207_1776 ();
 FILLCELL_X32 FILLER_207_1808 ();
 FILLCELL_X32 FILLER_207_1840 ();
 FILLCELL_X16 FILLER_207_1872 ();
 FILLCELL_X8 FILLER_207_1888 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X32 FILLER_208_1592 ();
 FILLCELL_X32 FILLER_208_1624 ();
 FILLCELL_X32 FILLER_208_1656 ();
 FILLCELL_X32 FILLER_208_1688 ();
 FILLCELL_X32 FILLER_208_1720 ();
 FILLCELL_X32 FILLER_208_1752 ();
 FILLCELL_X32 FILLER_208_1784 ();
 FILLCELL_X32 FILLER_208_1816 ();
 FILLCELL_X32 FILLER_208_1848 ();
 FILLCELL_X8 FILLER_208_1880 ();
 FILLCELL_X4 FILLER_208_1888 ();
 FILLCELL_X2 FILLER_208_1892 ();
 FILLCELL_X1 FILLER_208_1895 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X32 FILLER_209_1744 ();
 FILLCELL_X32 FILLER_209_1776 ();
 FILLCELL_X32 FILLER_209_1808 ();
 FILLCELL_X32 FILLER_209_1840 ();
 FILLCELL_X16 FILLER_209_1872 ();
 FILLCELL_X8 FILLER_209_1888 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X32 FILLER_210_1752 ();
 FILLCELL_X32 FILLER_210_1784 ();
 FILLCELL_X32 FILLER_210_1816 ();
 FILLCELL_X32 FILLER_210_1848 ();
 FILLCELL_X8 FILLER_210_1880 ();
 FILLCELL_X4 FILLER_210_1888 ();
 FILLCELL_X2 FILLER_210_1892 ();
 FILLCELL_X1 FILLER_210_1895 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X32 FILLER_211_1744 ();
 FILLCELL_X32 FILLER_211_1776 ();
 FILLCELL_X32 FILLER_211_1808 ();
 FILLCELL_X32 FILLER_211_1840 ();
 FILLCELL_X16 FILLER_211_1872 ();
 FILLCELL_X8 FILLER_211_1888 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X32 FILLER_212_1752 ();
 FILLCELL_X32 FILLER_212_1784 ();
 FILLCELL_X32 FILLER_212_1816 ();
 FILLCELL_X32 FILLER_212_1848 ();
 FILLCELL_X8 FILLER_212_1880 ();
 FILLCELL_X4 FILLER_212_1888 ();
 FILLCELL_X2 FILLER_212_1892 ();
 FILLCELL_X1 FILLER_212_1895 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X32 FILLER_213_1744 ();
 FILLCELL_X32 FILLER_213_1776 ();
 FILLCELL_X32 FILLER_213_1808 ();
 FILLCELL_X32 FILLER_213_1840 ();
 FILLCELL_X16 FILLER_213_1872 ();
 FILLCELL_X8 FILLER_213_1888 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X32 FILLER_214_1752 ();
 FILLCELL_X32 FILLER_214_1784 ();
 FILLCELL_X32 FILLER_214_1816 ();
 FILLCELL_X32 FILLER_214_1848 ();
 FILLCELL_X8 FILLER_214_1880 ();
 FILLCELL_X4 FILLER_214_1888 ();
 FILLCELL_X2 FILLER_214_1892 ();
 FILLCELL_X1 FILLER_214_1895 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X32 FILLER_215_1744 ();
 FILLCELL_X32 FILLER_215_1776 ();
 FILLCELL_X32 FILLER_215_1808 ();
 FILLCELL_X32 FILLER_215_1840 ();
 FILLCELL_X16 FILLER_215_1872 ();
 FILLCELL_X8 FILLER_215_1888 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X32 FILLER_216_1752 ();
 FILLCELL_X32 FILLER_216_1784 ();
 FILLCELL_X32 FILLER_216_1816 ();
 FILLCELL_X32 FILLER_216_1848 ();
 FILLCELL_X8 FILLER_216_1880 ();
 FILLCELL_X4 FILLER_216_1888 ();
 FILLCELL_X2 FILLER_216_1892 ();
 FILLCELL_X1 FILLER_216_1895 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X32 FILLER_217_1744 ();
 FILLCELL_X32 FILLER_217_1776 ();
 FILLCELL_X32 FILLER_217_1808 ();
 FILLCELL_X32 FILLER_217_1840 ();
 FILLCELL_X16 FILLER_217_1872 ();
 FILLCELL_X8 FILLER_217_1888 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X32 FILLER_218_1752 ();
 FILLCELL_X32 FILLER_218_1784 ();
 FILLCELL_X32 FILLER_218_1816 ();
 FILLCELL_X32 FILLER_218_1848 ();
 FILLCELL_X8 FILLER_218_1880 ();
 FILLCELL_X4 FILLER_218_1888 ();
 FILLCELL_X2 FILLER_218_1892 ();
 FILLCELL_X1 FILLER_218_1895 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X32 FILLER_219_1744 ();
 FILLCELL_X32 FILLER_219_1776 ();
 FILLCELL_X32 FILLER_219_1808 ();
 FILLCELL_X32 FILLER_219_1840 ();
 FILLCELL_X16 FILLER_219_1872 ();
 FILLCELL_X8 FILLER_219_1888 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X32 FILLER_220_1752 ();
 FILLCELL_X32 FILLER_220_1784 ();
 FILLCELL_X32 FILLER_220_1816 ();
 FILLCELL_X32 FILLER_220_1848 ();
 FILLCELL_X8 FILLER_220_1880 ();
 FILLCELL_X4 FILLER_220_1888 ();
 FILLCELL_X2 FILLER_220_1892 ();
 FILLCELL_X1 FILLER_220_1895 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X32 FILLER_221_1744 ();
 FILLCELL_X32 FILLER_221_1776 ();
 FILLCELL_X32 FILLER_221_1808 ();
 FILLCELL_X32 FILLER_221_1840 ();
 FILLCELL_X16 FILLER_221_1872 ();
 FILLCELL_X8 FILLER_221_1888 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X32 FILLER_222_1720 ();
 FILLCELL_X32 FILLER_222_1752 ();
 FILLCELL_X32 FILLER_222_1784 ();
 FILLCELL_X32 FILLER_222_1816 ();
 FILLCELL_X32 FILLER_222_1848 ();
 FILLCELL_X8 FILLER_222_1880 ();
 FILLCELL_X4 FILLER_222_1888 ();
 FILLCELL_X2 FILLER_222_1892 ();
 FILLCELL_X1 FILLER_222_1895 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X32 FILLER_223_1744 ();
 FILLCELL_X32 FILLER_223_1776 ();
 FILLCELL_X32 FILLER_223_1808 ();
 FILLCELL_X32 FILLER_223_1840 ();
 FILLCELL_X16 FILLER_223_1872 ();
 FILLCELL_X8 FILLER_223_1888 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X32 FILLER_224_1752 ();
 FILLCELL_X32 FILLER_224_1784 ();
 FILLCELL_X32 FILLER_224_1816 ();
 FILLCELL_X32 FILLER_224_1848 ();
 FILLCELL_X8 FILLER_224_1880 ();
 FILLCELL_X4 FILLER_224_1888 ();
 FILLCELL_X2 FILLER_224_1892 ();
 FILLCELL_X1 FILLER_224_1895 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X32 FILLER_225_1744 ();
 FILLCELL_X32 FILLER_225_1776 ();
 FILLCELL_X32 FILLER_225_1808 ();
 FILLCELL_X32 FILLER_225_1840 ();
 FILLCELL_X16 FILLER_225_1872 ();
 FILLCELL_X8 FILLER_225_1888 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X32 FILLER_226_1752 ();
 FILLCELL_X32 FILLER_226_1784 ();
 FILLCELL_X32 FILLER_226_1816 ();
 FILLCELL_X32 FILLER_226_1848 ();
 FILLCELL_X8 FILLER_226_1880 ();
 FILLCELL_X4 FILLER_226_1888 ();
 FILLCELL_X2 FILLER_226_1892 ();
 FILLCELL_X1 FILLER_226_1895 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X32 FILLER_227_1744 ();
 FILLCELL_X32 FILLER_227_1776 ();
 FILLCELL_X32 FILLER_227_1808 ();
 FILLCELL_X32 FILLER_227_1840 ();
 FILLCELL_X16 FILLER_227_1872 ();
 FILLCELL_X8 FILLER_227_1888 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X32 FILLER_228_1752 ();
 FILLCELL_X32 FILLER_228_1784 ();
 FILLCELL_X32 FILLER_228_1816 ();
 FILLCELL_X32 FILLER_228_1848 ();
 FILLCELL_X8 FILLER_228_1880 ();
 FILLCELL_X4 FILLER_228_1888 ();
 FILLCELL_X2 FILLER_228_1892 ();
 FILLCELL_X1 FILLER_228_1895 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X32 FILLER_229_1744 ();
 FILLCELL_X32 FILLER_229_1776 ();
 FILLCELL_X32 FILLER_229_1808 ();
 FILLCELL_X32 FILLER_229_1840 ();
 FILLCELL_X16 FILLER_229_1872 ();
 FILLCELL_X8 FILLER_229_1888 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X32 FILLER_230_1752 ();
 FILLCELL_X32 FILLER_230_1784 ();
 FILLCELL_X32 FILLER_230_1816 ();
 FILLCELL_X32 FILLER_230_1848 ();
 FILLCELL_X8 FILLER_230_1880 ();
 FILLCELL_X4 FILLER_230_1888 ();
 FILLCELL_X2 FILLER_230_1892 ();
 FILLCELL_X1 FILLER_230_1895 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X32 FILLER_231_1744 ();
 FILLCELL_X32 FILLER_231_1776 ();
 FILLCELL_X32 FILLER_231_1808 ();
 FILLCELL_X32 FILLER_231_1840 ();
 FILLCELL_X16 FILLER_231_1872 ();
 FILLCELL_X8 FILLER_231_1888 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X32 FILLER_232_1720 ();
 FILLCELL_X32 FILLER_232_1752 ();
 FILLCELL_X32 FILLER_232_1784 ();
 FILLCELL_X32 FILLER_232_1816 ();
 FILLCELL_X32 FILLER_232_1848 ();
 FILLCELL_X8 FILLER_232_1880 ();
 FILLCELL_X4 FILLER_232_1888 ();
 FILLCELL_X2 FILLER_232_1892 ();
 FILLCELL_X1 FILLER_232_1895 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X32 FILLER_233_1744 ();
 FILLCELL_X32 FILLER_233_1776 ();
 FILLCELL_X32 FILLER_233_1808 ();
 FILLCELL_X32 FILLER_233_1840 ();
 FILLCELL_X16 FILLER_233_1872 ();
 FILLCELL_X8 FILLER_233_1888 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X32 FILLER_234_1752 ();
 FILLCELL_X32 FILLER_234_1784 ();
 FILLCELL_X32 FILLER_234_1816 ();
 FILLCELL_X32 FILLER_234_1848 ();
 FILLCELL_X8 FILLER_234_1880 ();
 FILLCELL_X4 FILLER_234_1888 ();
 FILLCELL_X2 FILLER_234_1892 ();
 FILLCELL_X1 FILLER_234_1895 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X32 FILLER_235_1744 ();
 FILLCELL_X32 FILLER_235_1776 ();
 FILLCELL_X32 FILLER_235_1808 ();
 FILLCELL_X32 FILLER_235_1840 ();
 FILLCELL_X16 FILLER_235_1872 ();
 FILLCELL_X8 FILLER_235_1888 ();
 FILLCELL_X32 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_33 ();
 FILLCELL_X32 FILLER_236_65 ();
 FILLCELL_X32 FILLER_236_97 ();
 FILLCELL_X32 FILLER_236_129 ();
 FILLCELL_X32 FILLER_236_161 ();
 FILLCELL_X32 FILLER_236_193 ();
 FILLCELL_X32 FILLER_236_225 ();
 FILLCELL_X32 FILLER_236_257 ();
 FILLCELL_X32 FILLER_236_289 ();
 FILLCELL_X32 FILLER_236_321 ();
 FILLCELL_X32 FILLER_236_353 ();
 FILLCELL_X32 FILLER_236_385 ();
 FILLCELL_X32 FILLER_236_417 ();
 FILLCELL_X32 FILLER_236_449 ();
 FILLCELL_X32 FILLER_236_481 ();
 FILLCELL_X32 FILLER_236_513 ();
 FILLCELL_X32 FILLER_236_545 ();
 FILLCELL_X32 FILLER_236_577 ();
 FILLCELL_X16 FILLER_236_609 ();
 FILLCELL_X4 FILLER_236_625 ();
 FILLCELL_X2 FILLER_236_629 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X32 FILLER_236_1752 ();
 FILLCELL_X32 FILLER_236_1784 ();
 FILLCELL_X32 FILLER_236_1816 ();
 FILLCELL_X32 FILLER_236_1848 ();
 FILLCELL_X8 FILLER_236_1880 ();
 FILLCELL_X4 FILLER_236_1888 ();
 FILLCELL_X2 FILLER_236_1892 ();
 FILLCELL_X1 FILLER_236_1895 ();
 FILLCELL_X32 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_33 ();
 FILLCELL_X32 FILLER_237_65 ();
 FILLCELL_X32 FILLER_237_97 ();
 FILLCELL_X32 FILLER_237_129 ();
 FILLCELL_X32 FILLER_237_161 ();
 FILLCELL_X32 FILLER_237_193 ();
 FILLCELL_X32 FILLER_237_225 ();
 FILLCELL_X32 FILLER_237_257 ();
 FILLCELL_X32 FILLER_237_289 ();
 FILLCELL_X32 FILLER_237_321 ();
 FILLCELL_X32 FILLER_237_353 ();
 FILLCELL_X32 FILLER_237_385 ();
 FILLCELL_X32 FILLER_237_417 ();
 FILLCELL_X32 FILLER_237_449 ();
 FILLCELL_X32 FILLER_237_481 ();
 FILLCELL_X32 FILLER_237_513 ();
 FILLCELL_X32 FILLER_237_545 ();
 FILLCELL_X32 FILLER_237_577 ();
 FILLCELL_X32 FILLER_237_609 ();
 FILLCELL_X32 FILLER_237_641 ();
 FILLCELL_X32 FILLER_237_673 ();
 FILLCELL_X32 FILLER_237_705 ();
 FILLCELL_X32 FILLER_237_737 ();
 FILLCELL_X32 FILLER_237_769 ();
 FILLCELL_X32 FILLER_237_801 ();
 FILLCELL_X32 FILLER_237_833 ();
 FILLCELL_X32 FILLER_237_865 ();
 FILLCELL_X32 FILLER_237_897 ();
 FILLCELL_X32 FILLER_237_929 ();
 FILLCELL_X32 FILLER_237_961 ();
 FILLCELL_X32 FILLER_237_993 ();
 FILLCELL_X32 FILLER_237_1025 ();
 FILLCELL_X32 FILLER_237_1057 ();
 FILLCELL_X32 FILLER_237_1089 ();
 FILLCELL_X32 FILLER_237_1121 ();
 FILLCELL_X32 FILLER_237_1153 ();
 FILLCELL_X32 FILLER_237_1185 ();
 FILLCELL_X32 FILLER_237_1217 ();
 FILLCELL_X8 FILLER_237_1249 ();
 FILLCELL_X4 FILLER_237_1257 ();
 FILLCELL_X2 FILLER_237_1261 ();
 FILLCELL_X32 FILLER_237_1264 ();
 FILLCELL_X32 FILLER_237_1296 ();
 FILLCELL_X32 FILLER_237_1328 ();
 FILLCELL_X32 FILLER_237_1360 ();
 FILLCELL_X32 FILLER_237_1392 ();
 FILLCELL_X32 FILLER_237_1424 ();
 FILLCELL_X32 FILLER_237_1456 ();
 FILLCELL_X32 FILLER_237_1488 ();
 FILLCELL_X32 FILLER_237_1520 ();
 FILLCELL_X32 FILLER_237_1552 ();
 FILLCELL_X32 FILLER_237_1584 ();
 FILLCELL_X32 FILLER_237_1616 ();
 FILLCELL_X32 FILLER_237_1648 ();
 FILLCELL_X32 FILLER_237_1680 ();
 FILLCELL_X32 FILLER_237_1712 ();
 FILLCELL_X32 FILLER_237_1744 ();
 FILLCELL_X32 FILLER_237_1776 ();
 FILLCELL_X32 FILLER_237_1808 ();
 FILLCELL_X32 FILLER_237_1840 ();
 FILLCELL_X16 FILLER_237_1872 ();
 FILLCELL_X8 FILLER_237_1888 ();
 FILLCELL_X32 FILLER_238_1 ();
 FILLCELL_X32 FILLER_238_33 ();
 FILLCELL_X32 FILLER_238_65 ();
 FILLCELL_X32 FILLER_238_97 ();
 FILLCELL_X32 FILLER_238_129 ();
 FILLCELL_X32 FILLER_238_161 ();
 FILLCELL_X32 FILLER_238_193 ();
 FILLCELL_X32 FILLER_238_225 ();
 FILLCELL_X32 FILLER_238_257 ();
 FILLCELL_X32 FILLER_238_289 ();
 FILLCELL_X32 FILLER_238_321 ();
 FILLCELL_X32 FILLER_238_353 ();
 FILLCELL_X32 FILLER_238_385 ();
 FILLCELL_X32 FILLER_238_417 ();
 FILLCELL_X32 FILLER_238_449 ();
 FILLCELL_X32 FILLER_238_481 ();
 FILLCELL_X32 FILLER_238_513 ();
 FILLCELL_X32 FILLER_238_545 ();
 FILLCELL_X32 FILLER_238_577 ();
 FILLCELL_X16 FILLER_238_609 ();
 FILLCELL_X4 FILLER_238_625 ();
 FILLCELL_X2 FILLER_238_629 ();
 FILLCELL_X32 FILLER_238_632 ();
 FILLCELL_X32 FILLER_238_664 ();
 FILLCELL_X32 FILLER_238_696 ();
 FILLCELL_X32 FILLER_238_728 ();
 FILLCELL_X32 FILLER_238_760 ();
 FILLCELL_X32 FILLER_238_792 ();
 FILLCELL_X32 FILLER_238_824 ();
 FILLCELL_X32 FILLER_238_856 ();
 FILLCELL_X32 FILLER_238_888 ();
 FILLCELL_X32 FILLER_238_920 ();
 FILLCELL_X32 FILLER_238_952 ();
 FILLCELL_X32 FILLER_238_984 ();
 FILLCELL_X32 FILLER_238_1016 ();
 FILLCELL_X32 FILLER_238_1048 ();
 FILLCELL_X32 FILLER_238_1080 ();
 FILLCELL_X32 FILLER_238_1112 ();
 FILLCELL_X32 FILLER_238_1144 ();
 FILLCELL_X32 FILLER_238_1176 ();
 FILLCELL_X32 FILLER_238_1208 ();
 FILLCELL_X32 FILLER_238_1240 ();
 FILLCELL_X32 FILLER_238_1272 ();
 FILLCELL_X32 FILLER_238_1304 ();
 FILLCELL_X32 FILLER_238_1336 ();
 FILLCELL_X32 FILLER_238_1368 ();
 FILLCELL_X32 FILLER_238_1400 ();
 FILLCELL_X32 FILLER_238_1432 ();
 FILLCELL_X32 FILLER_238_1464 ();
 FILLCELL_X32 FILLER_238_1496 ();
 FILLCELL_X32 FILLER_238_1528 ();
 FILLCELL_X32 FILLER_238_1560 ();
 FILLCELL_X32 FILLER_238_1592 ();
 FILLCELL_X32 FILLER_238_1624 ();
 FILLCELL_X32 FILLER_238_1656 ();
 FILLCELL_X32 FILLER_238_1688 ();
 FILLCELL_X32 FILLER_238_1720 ();
 FILLCELL_X32 FILLER_238_1752 ();
 FILLCELL_X32 FILLER_238_1784 ();
 FILLCELL_X32 FILLER_238_1816 ();
 FILLCELL_X32 FILLER_238_1848 ();
 FILLCELL_X8 FILLER_238_1880 ();
 FILLCELL_X4 FILLER_238_1888 ();
 FILLCELL_X2 FILLER_238_1892 ();
 FILLCELL_X1 FILLER_238_1895 ();
 FILLCELL_X32 FILLER_239_1 ();
 FILLCELL_X32 FILLER_239_33 ();
 FILLCELL_X32 FILLER_239_65 ();
 FILLCELL_X32 FILLER_239_97 ();
 FILLCELL_X32 FILLER_239_129 ();
 FILLCELL_X32 FILLER_239_161 ();
 FILLCELL_X32 FILLER_239_193 ();
 FILLCELL_X32 FILLER_239_225 ();
 FILLCELL_X32 FILLER_239_257 ();
 FILLCELL_X32 FILLER_239_289 ();
 FILLCELL_X32 FILLER_239_321 ();
 FILLCELL_X32 FILLER_239_353 ();
 FILLCELL_X32 FILLER_239_385 ();
 FILLCELL_X32 FILLER_239_417 ();
 FILLCELL_X32 FILLER_239_449 ();
 FILLCELL_X32 FILLER_239_481 ();
 FILLCELL_X32 FILLER_239_513 ();
 FILLCELL_X32 FILLER_239_545 ();
 FILLCELL_X32 FILLER_239_577 ();
 FILLCELL_X32 FILLER_239_609 ();
 FILLCELL_X32 FILLER_239_641 ();
 FILLCELL_X32 FILLER_239_673 ();
 FILLCELL_X32 FILLER_239_705 ();
 FILLCELL_X32 FILLER_239_737 ();
 FILLCELL_X32 FILLER_239_769 ();
 FILLCELL_X32 FILLER_239_801 ();
 FILLCELL_X32 FILLER_239_833 ();
 FILLCELL_X32 FILLER_239_865 ();
 FILLCELL_X32 FILLER_239_897 ();
 FILLCELL_X32 FILLER_239_929 ();
 FILLCELL_X32 FILLER_239_961 ();
 FILLCELL_X32 FILLER_239_993 ();
 FILLCELL_X32 FILLER_239_1025 ();
 FILLCELL_X32 FILLER_239_1057 ();
 FILLCELL_X32 FILLER_239_1089 ();
 FILLCELL_X32 FILLER_239_1121 ();
 FILLCELL_X32 FILLER_239_1153 ();
 FILLCELL_X32 FILLER_239_1185 ();
 FILLCELL_X32 FILLER_239_1217 ();
 FILLCELL_X8 FILLER_239_1249 ();
 FILLCELL_X4 FILLER_239_1257 ();
 FILLCELL_X2 FILLER_239_1261 ();
 FILLCELL_X32 FILLER_239_1264 ();
 FILLCELL_X32 FILLER_239_1296 ();
 FILLCELL_X32 FILLER_239_1328 ();
 FILLCELL_X32 FILLER_239_1360 ();
 FILLCELL_X32 FILLER_239_1392 ();
 FILLCELL_X32 FILLER_239_1424 ();
 FILLCELL_X32 FILLER_239_1456 ();
 FILLCELL_X32 FILLER_239_1488 ();
 FILLCELL_X32 FILLER_239_1520 ();
 FILLCELL_X32 FILLER_239_1552 ();
 FILLCELL_X32 FILLER_239_1584 ();
 FILLCELL_X32 FILLER_239_1616 ();
 FILLCELL_X32 FILLER_239_1648 ();
 FILLCELL_X32 FILLER_239_1680 ();
 FILLCELL_X32 FILLER_239_1712 ();
 FILLCELL_X32 FILLER_239_1744 ();
 FILLCELL_X32 FILLER_239_1776 ();
 FILLCELL_X32 FILLER_239_1808 ();
 FILLCELL_X32 FILLER_239_1840 ();
 FILLCELL_X16 FILLER_239_1872 ();
 FILLCELL_X8 FILLER_239_1888 ();
 FILLCELL_X32 FILLER_240_1 ();
 FILLCELL_X32 FILLER_240_33 ();
 FILLCELL_X32 FILLER_240_65 ();
 FILLCELL_X32 FILLER_240_97 ();
 FILLCELL_X32 FILLER_240_129 ();
 FILLCELL_X32 FILLER_240_161 ();
 FILLCELL_X32 FILLER_240_193 ();
 FILLCELL_X32 FILLER_240_225 ();
 FILLCELL_X32 FILLER_240_257 ();
 FILLCELL_X32 FILLER_240_289 ();
 FILLCELL_X32 FILLER_240_321 ();
 FILLCELL_X32 FILLER_240_353 ();
 FILLCELL_X32 FILLER_240_385 ();
 FILLCELL_X32 FILLER_240_417 ();
 FILLCELL_X32 FILLER_240_449 ();
 FILLCELL_X32 FILLER_240_481 ();
 FILLCELL_X32 FILLER_240_513 ();
 FILLCELL_X32 FILLER_240_545 ();
 FILLCELL_X32 FILLER_240_577 ();
 FILLCELL_X16 FILLER_240_609 ();
 FILLCELL_X4 FILLER_240_625 ();
 FILLCELL_X2 FILLER_240_629 ();
 FILLCELL_X32 FILLER_240_632 ();
 FILLCELL_X32 FILLER_240_664 ();
 FILLCELL_X32 FILLER_240_696 ();
 FILLCELL_X32 FILLER_240_728 ();
 FILLCELL_X32 FILLER_240_760 ();
 FILLCELL_X32 FILLER_240_792 ();
 FILLCELL_X32 FILLER_240_824 ();
 FILLCELL_X32 FILLER_240_856 ();
 FILLCELL_X32 FILLER_240_888 ();
 FILLCELL_X32 FILLER_240_920 ();
 FILLCELL_X32 FILLER_240_952 ();
 FILLCELL_X32 FILLER_240_984 ();
 FILLCELL_X32 FILLER_240_1016 ();
 FILLCELL_X32 FILLER_240_1048 ();
 FILLCELL_X32 FILLER_240_1080 ();
 FILLCELL_X32 FILLER_240_1112 ();
 FILLCELL_X32 FILLER_240_1144 ();
 FILLCELL_X32 FILLER_240_1176 ();
 FILLCELL_X32 FILLER_240_1208 ();
 FILLCELL_X32 FILLER_240_1240 ();
 FILLCELL_X32 FILLER_240_1272 ();
 FILLCELL_X32 FILLER_240_1304 ();
 FILLCELL_X32 FILLER_240_1336 ();
 FILLCELL_X32 FILLER_240_1368 ();
 FILLCELL_X32 FILLER_240_1400 ();
 FILLCELL_X32 FILLER_240_1432 ();
 FILLCELL_X32 FILLER_240_1464 ();
 FILLCELL_X32 FILLER_240_1496 ();
 FILLCELL_X32 FILLER_240_1528 ();
 FILLCELL_X32 FILLER_240_1560 ();
 FILLCELL_X32 FILLER_240_1592 ();
 FILLCELL_X32 FILLER_240_1624 ();
 FILLCELL_X32 FILLER_240_1656 ();
 FILLCELL_X32 FILLER_240_1688 ();
 FILLCELL_X32 FILLER_240_1720 ();
 FILLCELL_X32 FILLER_240_1752 ();
 FILLCELL_X32 FILLER_240_1784 ();
 FILLCELL_X32 FILLER_240_1816 ();
 FILLCELL_X32 FILLER_240_1848 ();
 FILLCELL_X8 FILLER_240_1880 ();
 FILLCELL_X4 FILLER_240_1888 ();
 FILLCELL_X2 FILLER_240_1892 ();
 FILLCELL_X1 FILLER_240_1895 ();
 FILLCELL_X32 FILLER_241_1 ();
 FILLCELL_X32 FILLER_241_33 ();
 FILLCELL_X32 FILLER_241_65 ();
 FILLCELL_X32 FILLER_241_97 ();
 FILLCELL_X32 FILLER_241_129 ();
 FILLCELL_X32 FILLER_241_161 ();
 FILLCELL_X32 FILLER_241_193 ();
 FILLCELL_X32 FILLER_241_225 ();
 FILLCELL_X32 FILLER_241_257 ();
 FILLCELL_X32 FILLER_241_289 ();
 FILLCELL_X32 FILLER_241_321 ();
 FILLCELL_X32 FILLER_241_353 ();
 FILLCELL_X32 FILLER_241_385 ();
 FILLCELL_X32 FILLER_241_417 ();
 FILLCELL_X32 FILLER_241_449 ();
 FILLCELL_X32 FILLER_241_481 ();
 FILLCELL_X32 FILLER_241_513 ();
 FILLCELL_X32 FILLER_241_545 ();
 FILLCELL_X32 FILLER_241_577 ();
 FILLCELL_X32 FILLER_241_609 ();
 FILLCELL_X32 FILLER_241_641 ();
 FILLCELL_X32 FILLER_241_673 ();
 FILLCELL_X32 FILLER_241_705 ();
 FILLCELL_X32 FILLER_241_737 ();
 FILLCELL_X32 FILLER_241_769 ();
 FILLCELL_X32 FILLER_241_801 ();
 FILLCELL_X32 FILLER_241_833 ();
 FILLCELL_X32 FILLER_241_865 ();
 FILLCELL_X32 FILLER_241_897 ();
 FILLCELL_X32 FILLER_241_929 ();
 FILLCELL_X32 FILLER_241_961 ();
 FILLCELL_X32 FILLER_241_993 ();
 FILLCELL_X32 FILLER_241_1025 ();
 FILLCELL_X32 FILLER_241_1057 ();
 FILLCELL_X32 FILLER_241_1089 ();
 FILLCELL_X32 FILLER_241_1121 ();
 FILLCELL_X32 FILLER_241_1153 ();
 FILLCELL_X32 FILLER_241_1185 ();
 FILLCELL_X32 FILLER_241_1217 ();
 FILLCELL_X8 FILLER_241_1249 ();
 FILLCELL_X4 FILLER_241_1257 ();
 FILLCELL_X2 FILLER_241_1261 ();
 FILLCELL_X32 FILLER_241_1264 ();
 FILLCELL_X32 FILLER_241_1296 ();
 FILLCELL_X32 FILLER_241_1328 ();
 FILLCELL_X32 FILLER_241_1360 ();
 FILLCELL_X32 FILLER_241_1392 ();
 FILLCELL_X32 FILLER_241_1424 ();
 FILLCELL_X32 FILLER_241_1456 ();
 FILLCELL_X32 FILLER_241_1488 ();
 FILLCELL_X32 FILLER_241_1520 ();
 FILLCELL_X32 FILLER_241_1552 ();
 FILLCELL_X32 FILLER_241_1584 ();
 FILLCELL_X32 FILLER_241_1616 ();
 FILLCELL_X32 FILLER_241_1648 ();
 FILLCELL_X32 FILLER_241_1680 ();
 FILLCELL_X32 FILLER_241_1712 ();
 FILLCELL_X32 FILLER_241_1744 ();
 FILLCELL_X32 FILLER_241_1776 ();
 FILLCELL_X32 FILLER_241_1808 ();
 FILLCELL_X32 FILLER_241_1840 ();
 FILLCELL_X16 FILLER_241_1872 ();
 FILLCELL_X8 FILLER_241_1888 ();
 FILLCELL_X32 FILLER_242_1 ();
 FILLCELL_X32 FILLER_242_33 ();
 FILLCELL_X32 FILLER_242_65 ();
 FILLCELL_X32 FILLER_242_97 ();
 FILLCELL_X32 FILLER_242_129 ();
 FILLCELL_X32 FILLER_242_161 ();
 FILLCELL_X32 FILLER_242_193 ();
 FILLCELL_X32 FILLER_242_225 ();
 FILLCELL_X32 FILLER_242_257 ();
 FILLCELL_X32 FILLER_242_289 ();
 FILLCELL_X32 FILLER_242_321 ();
 FILLCELL_X32 FILLER_242_353 ();
 FILLCELL_X32 FILLER_242_385 ();
 FILLCELL_X32 FILLER_242_417 ();
 FILLCELL_X32 FILLER_242_449 ();
 FILLCELL_X32 FILLER_242_481 ();
 FILLCELL_X32 FILLER_242_513 ();
 FILLCELL_X32 FILLER_242_545 ();
 FILLCELL_X32 FILLER_242_577 ();
 FILLCELL_X16 FILLER_242_609 ();
 FILLCELL_X4 FILLER_242_625 ();
 FILLCELL_X2 FILLER_242_629 ();
 FILLCELL_X32 FILLER_242_632 ();
 FILLCELL_X32 FILLER_242_664 ();
 FILLCELL_X32 FILLER_242_696 ();
 FILLCELL_X32 FILLER_242_728 ();
 FILLCELL_X32 FILLER_242_760 ();
 FILLCELL_X32 FILLER_242_792 ();
 FILLCELL_X32 FILLER_242_824 ();
 FILLCELL_X32 FILLER_242_856 ();
 FILLCELL_X32 FILLER_242_888 ();
 FILLCELL_X32 FILLER_242_920 ();
 FILLCELL_X32 FILLER_242_952 ();
 FILLCELL_X32 FILLER_242_984 ();
 FILLCELL_X32 FILLER_242_1016 ();
 FILLCELL_X32 FILLER_242_1048 ();
 FILLCELL_X32 FILLER_242_1080 ();
 FILLCELL_X32 FILLER_242_1112 ();
 FILLCELL_X32 FILLER_242_1144 ();
 FILLCELL_X32 FILLER_242_1176 ();
 FILLCELL_X32 FILLER_242_1208 ();
 FILLCELL_X32 FILLER_242_1240 ();
 FILLCELL_X32 FILLER_242_1272 ();
 FILLCELL_X32 FILLER_242_1304 ();
 FILLCELL_X32 FILLER_242_1336 ();
 FILLCELL_X32 FILLER_242_1368 ();
 FILLCELL_X32 FILLER_242_1400 ();
 FILLCELL_X32 FILLER_242_1432 ();
 FILLCELL_X32 FILLER_242_1464 ();
 FILLCELL_X32 FILLER_242_1496 ();
 FILLCELL_X32 FILLER_242_1528 ();
 FILLCELL_X32 FILLER_242_1560 ();
 FILLCELL_X32 FILLER_242_1592 ();
 FILLCELL_X32 FILLER_242_1624 ();
 FILLCELL_X32 FILLER_242_1656 ();
 FILLCELL_X32 FILLER_242_1688 ();
 FILLCELL_X32 FILLER_242_1720 ();
 FILLCELL_X32 FILLER_242_1752 ();
 FILLCELL_X32 FILLER_242_1784 ();
 FILLCELL_X32 FILLER_242_1816 ();
 FILLCELL_X32 FILLER_242_1848 ();
 FILLCELL_X8 FILLER_242_1880 ();
 FILLCELL_X4 FILLER_242_1888 ();
 FILLCELL_X2 FILLER_242_1892 ();
 FILLCELL_X1 FILLER_242_1895 ();
 FILLCELL_X32 FILLER_243_1 ();
 FILLCELL_X32 FILLER_243_33 ();
 FILLCELL_X32 FILLER_243_65 ();
 FILLCELL_X32 FILLER_243_97 ();
 FILLCELL_X32 FILLER_243_129 ();
 FILLCELL_X32 FILLER_243_161 ();
 FILLCELL_X32 FILLER_243_193 ();
 FILLCELL_X32 FILLER_243_225 ();
 FILLCELL_X32 FILLER_243_257 ();
 FILLCELL_X32 FILLER_243_289 ();
 FILLCELL_X32 FILLER_243_321 ();
 FILLCELL_X32 FILLER_243_353 ();
 FILLCELL_X32 FILLER_243_385 ();
 FILLCELL_X32 FILLER_243_417 ();
 FILLCELL_X32 FILLER_243_449 ();
 FILLCELL_X32 FILLER_243_481 ();
 FILLCELL_X32 FILLER_243_513 ();
 FILLCELL_X32 FILLER_243_545 ();
 FILLCELL_X32 FILLER_243_577 ();
 FILLCELL_X32 FILLER_243_609 ();
 FILLCELL_X32 FILLER_243_641 ();
 FILLCELL_X32 FILLER_243_673 ();
 FILLCELL_X32 FILLER_243_705 ();
 FILLCELL_X32 FILLER_243_737 ();
 FILLCELL_X32 FILLER_243_769 ();
 FILLCELL_X32 FILLER_243_801 ();
 FILLCELL_X32 FILLER_243_833 ();
 FILLCELL_X32 FILLER_243_865 ();
 FILLCELL_X32 FILLER_243_897 ();
 FILLCELL_X32 FILLER_243_929 ();
 FILLCELL_X32 FILLER_243_961 ();
 FILLCELL_X32 FILLER_243_993 ();
 FILLCELL_X32 FILLER_243_1025 ();
 FILLCELL_X32 FILLER_243_1057 ();
 FILLCELL_X32 FILLER_243_1089 ();
 FILLCELL_X32 FILLER_243_1121 ();
 FILLCELL_X32 FILLER_243_1153 ();
 FILLCELL_X32 FILLER_243_1185 ();
 FILLCELL_X32 FILLER_243_1217 ();
 FILLCELL_X8 FILLER_243_1249 ();
 FILLCELL_X4 FILLER_243_1257 ();
 FILLCELL_X2 FILLER_243_1261 ();
 FILLCELL_X32 FILLER_243_1264 ();
 FILLCELL_X32 FILLER_243_1296 ();
 FILLCELL_X32 FILLER_243_1328 ();
 FILLCELL_X32 FILLER_243_1360 ();
 FILLCELL_X32 FILLER_243_1392 ();
 FILLCELL_X32 FILLER_243_1424 ();
 FILLCELL_X32 FILLER_243_1456 ();
 FILLCELL_X32 FILLER_243_1488 ();
 FILLCELL_X32 FILLER_243_1520 ();
 FILLCELL_X32 FILLER_243_1552 ();
 FILLCELL_X32 FILLER_243_1584 ();
 FILLCELL_X32 FILLER_243_1616 ();
 FILLCELL_X32 FILLER_243_1648 ();
 FILLCELL_X32 FILLER_243_1680 ();
 FILLCELL_X32 FILLER_243_1712 ();
 FILLCELL_X32 FILLER_243_1744 ();
 FILLCELL_X32 FILLER_243_1776 ();
 FILLCELL_X32 FILLER_243_1808 ();
 FILLCELL_X32 FILLER_243_1840 ();
 FILLCELL_X16 FILLER_243_1872 ();
 FILLCELL_X8 FILLER_243_1888 ();
 FILLCELL_X32 FILLER_244_1 ();
 FILLCELL_X32 FILLER_244_33 ();
 FILLCELL_X32 FILLER_244_65 ();
 FILLCELL_X32 FILLER_244_97 ();
 FILLCELL_X32 FILLER_244_129 ();
 FILLCELL_X32 FILLER_244_161 ();
 FILLCELL_X32 FILLER_244_193 ();
 FILLCELL_X32 FILLER_244_225 ();
 FILLCELL_X32 FILLER_244_257 ();
 FILLCELL_X32 FILLER_244_289 ();
 FILLCELL_X32 FILLER_244_321 ();
 FILLCELL_X32 FILLER_244_353 ();
 FILLCELL_X32 FILLER_244_385 ();
 FILLCELL_X32 FILLER_244_417 ();
 FILLCELL_X32 FILLER_244_449 ();
 FILLCELL_X32 FILLER_244_481 ();
 FILLCELL_X32 FILLER_244_513 ();
 FILLCELL_X32 FILLER_244_545 ();
 FILLCELL_X32 FILLER_244_577 ();
 FILLCELL_X16 FILLER_244_609 ();
 FILLCELL_X4 FILLER_244_625 ();
 FILLCELL_X2 FILLER_244_629 ();
 FILLCELL_X32 FILLER_244_632 ();
 FILLCELL_X32 FILLER_244_664 ();
 FILLCELL_X32 FILLER_244_696 ();
 FILLCELL_X32 FILLER_244_728 ();
 FILLCELL_X32 FILLER_244_760 ();
 FILLCELL_X32 FILLER_244_792 ();
 FILLCELL_X32 FILLER_244_824 ();
 FILLCELL_X32 FILLER_244_856 ();
 FILLCELL_X32 FILLER_244_888 ();
 FILLCELL_X32 FILLER_244_920 ();
 FILLCELL_X32 FILLER_244_952 ();
 FILLCELL_X32 FILLER_244_984 ();
 FILLCELL_X32 FILLER_244_1016 ();
 FILLCELL_X32 FILLER_244_1048 ();
 FILLCELL_X32 FILLER_244_1080 ();
 FILLCELL_X32 FILLER_244_1112 ();
 FILLCELL_X32 FILLER_244_1144 ();
 FILLCELL_X32 FILLER_244_1176 ();
 FILLCELL_X32 FILLER_244_1208 ();
 FILLCELL_X32 FILLER_244_1240 ();
 FILLCELL_X32 FILLER_244_1272 ();
 FILLCELL_X32 FILLER_244_1304 ();
 FILLCELL_X32 FILLER_244_1336 ();
 FILLCELL_X32 FILLER_244_1368 ();
 FILLCELL_X32 FILLER_244_1400 ();
 FILLCELL_X32 FILLER_244_1432 ();
 FILLCELL_X32 FILLER_244_1464 ();
 FILLCELL_X32 FILLER_244_1496 ();
 FILLCELL_X32 FILLER_244_1528 ();
 FILLCELL_X32 FILLER_244_1560 ();
 FILLCELL_X32 FILLER_244_1592 ();
 FILLCELL_X32 FILLER_244_1624 ();
 FILLCELL_X32 FILLER_244_1656 ();
 FILLCELL_X32 FILLER_244_1688 ();
 FILLCELL_X32 FILLER_244_1720 ();
 FILLCELL_X32 FILLER_244_1752 ();
 FILLCELL_X32 FILLER_244_1784 ();
 FILLCELL_X32 FILLER_244_1816 ();
 FILLCELL_X32 FILLER_244_1848 ();
 FILLCELL_X8 FILLER_244_1880 ();
 FILLCELL_X4 FILLER_244_1888 ();
 FILLCELL_X2 FILLER_244_1892 ();
 FILLCELL_X1 FILLER_244_1895 ();
 FILLCELL_X32 FILLER_245_1 ();
 FILLCELL_X32 FILLER_245_33 ();
 FILLCELL_X32 FILLER_245_65 ();
 FILLCELL_X32 FILLER_245_97 ();
 FILLCELL_X32 FILLER_245_129 ();
 FILLCELL_X32 FILLER_245_161 ();
 FILLCELL_X32 FILLER_245_193 ();
 FILLCELL_X32 FILLER_245_225 ();
 FILLCELL_X32 FILLER_245_257 ();
 FILLCELL_X32 FILLER_245_289 ();
 FILLCELL_X32 FILLER_245_321 ();
 FILLCELL_X32 FILLER_245_353 ();
 FILLCELL_X32 FILLER_245_385 ();
 FILLCELL_X32 FILLER_245_417 ();
 FILLCELL_X32 FILLER_245_449 ();
 FILLCELL_X32 FILLER_245_481 ();
 FILLCELL_X32 FILLER_245_513 ();
 FILLCELL_X32 FILLER_245_545 ();
 FILLCELL_X32 FILLER_245_577 ();
 FILLCELL_X32 FILLER_245_609 ();
 FILLCELL_X32 FILLER_245_641 ();
 FILLCELL_X32 FILLER_245_673 ();
 FILLCELL_X32 FILLER_245_705 ();
 FILLCELL_X32 FILLER_245_737 ();
 FILLCELL_X32 FILLER_245_769 ();
 FILLCELL_X32 FILLER_245_801 ();
 FILLCELL_X32 FILLER_245_833 ();
 FILLCELL_X32 FILLER_245_865 ();
 FILLCELL_X32 FILLER_245_897 ();
 FILLCELL_X32 FILLER_245_929 ();
 FILLCELL_X32 FILLER_245_961 ();
 FILLCELL_X32 FILLER_245_993 ();
 FILLCELL_X32 FILLER_245_1025 ();
 FILLCELL_X32 FILLER_245_1057 ();
 FILLCELL_X32 FILLER_245_1089 ();
 FILLCELL_X32 FILLER_245_1121 ();
 FILLCELL_X32 FILLER_245_1153 ();
 FILLCELL_X32 FILLER_245_1185 ();
 FILLCELL_X32 FILLER_245_1217 ();
 FILLCELL_X8 FILLER_245_1249 ();
 FILLCELL_X4 FILLER_245_1257 ();
 FILLCELL_X2 FILLER_245_1261 ();
 FILLCELL_X32 FILLER_245_1264 ();
 FILLCELL_X32 FILLER_245_1296 ();
 FILLCELL_X32 FILLER_245_1328 ();
 FILLCELL_X32 FILLER_245_1360 ();
 FILLCELL_X32 FILLER_245_1392 ();
 FILLCELL_X32 FILLER_245_1424 ();
 FILLCELL_X32 FILLER_245_1456 ();
 FILLCELL_X32 FILLER_245_1488 ();
 FILLCELL_X32 FILLER_245_1520 ();
 FILLCELL_X32 FILLER_245_1552 ();
 FILLCELL_X32 FILLER_245_1584 ();
 FILLCELL_X32 FILLER_245_1616 ();
 FILLCELL_X32 FILLER_245_1648 ();
 FILLCELL_X32 FILLER_245_1680 ();
 FILLCELL_X32 FILLER_245_1712 ();
 FILLCELL_X32 FILLER_245_1744 ();
 FILLCELL_X32 FILLER_245_1776 ();
 FILLCELL_X32 FILLER_245_1808 ();
 FILLCELL_X32 FILLER_245_1840 ();
 FILLCELL_X16 FILLER_245_1872 ();
 FILLCELL_X8 FILLER_245_1888 ();
 FILLCELL_X32 FILLER_246_1 ();
 FILLCELL_X32 FILLER_246_33 ();
 FILLCELL_X32 FILLER_246_65 ();
 FILLCELL_X32 FILLER_246_97 ();
 FILLCELL_X32 FILLER_246_129 ();
 FILLCELL_X32 FILLER_246_161 ();
 FILLCELL_X32 FILLER_246_193 ();
 FILLCELL_X32 FILLER_246_225 ();
 FILLCELL_X32 FILLER_246_257 ();
 FILLCELL_X32 FILLER_246_289 ();
 FILLCELL_X32 FILLER_246_321 ();
 FILLCELL_X32 FILLER_246_353 ();
 FILLCELL_X32 FILLER_246_385 ();
 FILLCELL_X32 FILLER_246_417 ();
 FILLCELL_X32 FILLER_246_449 ();
 FILLCELL_X32 FILLER_246_481 ();
 FILLCELL_X32 FILLER_246_513 ();
 FILLCELL_X32 FILLER_246_545 ();
 FILLCELL_X32 FILLER_246_577 ();
 FILLCELL_X16 FILLER_246_609 ();
 FILLCELL_X4 FILLER_246_625 ();
 FILLCELL_X2 FILLER_246_629 ();
 FILLCELL_X32 FILLER_246_632 ();
 FILLCELL_X32 FILLER_246_664 ();
 FILLCELL_X32 FILLER_246_696 ();
 FILLCELL_X32 FILLER_246_728 ();
 FILLCELL_X32 FILLER_246_760 ();
 FILLCELL_X32 FILLER_246_792 ();
 FILLCELL_X32 FILLER_246_824 ();
 FILLCELL_X32 FILLER_246_856 ();
 FILLCELL_X32 FILLER_246_888 ();
 FILLCELL_X32 FILLER_246_920 ();
 FILLCELL_X32 FILLER_246_952 ();
 FILLCELL_X32 FILLER_246_984 ();
 FILLCELL_X32 FILLER_246_1016 ();
 FILLCELL_X32 FILLER_246_1048 ();
 FILLCELL_X32 FILLER_246_1080 ();
 FILLCELL_X32 FILLER_246_1112 ();
 FILLCELL_X32 FILLER_246_1144 ();
 FILLCELL_X32 FILLER_246_1176 ();
 FILLCELL_X32 FILLER_246_1208 ();
 FILLCELL_X32 FILLER_246_1240 ();
 FILLCELL_X32 FILLER_246_1272 ();
 FILLCELL_X32 FILLER_246_1304 ();
 FILLCELL_X32 FILLER_246_1336 ();
 FILLCELL_X32 FILLER_246_1368 ();
 FILLCELL_X32 FILLER_246_1400 ();
 FILLCELL_X32 FILLER_246_1432 ();
 FILLCELL_X32 FILLER_246_1464 ();
 FILLCELL_X32 FILLER_246_1496 ();
 FILLCELL_X32 FILLER_246_1528 ();
 FILLCELL_X32 FILLER_246_1560 ();
 FILLCELL_X32 FILLER_246_1592 ();
 FILLCELL_X32 FILLER_246_1624 ();
 FILLCELL_X32 FILLER_246_1656 ();
 FILLCELL_X32 FILLER_246_1688 ();
 FILLCELL_X32 FILLER_246_1720 ();
 FILLCELL_X32 FILLER_246_1752 ();
 FILLCELL_X32 FILLER_246_1784 ();
 FILLCELL_X32 FILLER_246_1816 ();
 FILLCELL_X32 FILLER_246_1848 ();
 FILLCELL_X8 FILLER_246_1880 ();
 FILLCELL_X4 FILLER_246_1888 ();
 FILLCELL_X2 FILLER_246_1892 ();
 FILLCELL_X1 FILLER_246_1895 ();
 FILLCELL_X32 FILLER_247_1 ();
 FILLCELL_X32 FILLER_247_33 ();
 FILLCELL_X32 FILLER_247_65 ();
 FILLCELL_X32 FILLER_247_97 ();
 FILLCELL_X32 FILLER_247_129 ();
 FILLCELL_X32 FILLER_247_161 ();
 FILLCELL_X32 FILLER_247_193 ();
 FILLCELL_X32 FILLER_247_225 ();
 FILLCELL_X32 FILLER_247_257 ();
 FILLCELL_X32 FILLER_247_289 ();
 FILLCELL_X32 FILLER_247_321 ();
 FILLCELL_X32 FILLER_247_353 ();
 FILLCELL_X32 FILLER_247_385 ();
 FILLCELL_X32 FILLER_247_417 ();
 FILLCELL_X32 FILLER_247_449 ();
 FILLCELL_X32 FILLER_247_481 ();
 FILLCELL_X32 FILLER_247_513 ();
 FILLCELL_X32 FILLER_247_545 ();
 FILLCELL_X32 FILLER_247_577 ();
 FILLCELL_X32 FILLER_247_609 ();
 FILLCELL_X32 FILLER_247_641 ();
 FILLCELL_X32 FILLER_247_673 ();
 FILLCELL_X32 FILLER_247_705 ();
 FILLCELL_X32 FILLER_247_737 ();
 FILLCELL_X32 FILLER_247_769 ();
 FILLCELL_X32 FILLER_247_801 ();
 FILLCELL_X32 FILLER_247_833 ();
 FILLCELL_X32 FILLER_247_865 ();
 FILLCELL_X32 FILLER_247_897 ();
 FILLCELL_X32 FILLER_247_929 ();
 FILLCELL_X32 FILLER_247_961 ();
 FILLCELL_X32 FILLER_247_993 ();
 FILLCELL_X32 FILLER_247_1025 ();
 FILLCELL_X32 FILLER_247_1057 ();
 FILLCELL_X32 FILLER_247_1089 ();
 FILLCELL_X32 FILLER_247_1121 ();
 FILLCELL_X32 FILLER_247_1153 ();
 FILLCELL_X32 FILLER_247_1185 ();
 FILLCELL_X32 FILLER_247_1217 ();
 FILLCELL_X8 FILLER_247_1249 ();
 FILLCELL_X4 FILLER_247_1257 ();
 FILLCELL_X2 FILLER_247_1261 ();
 FILLCELL_X32 FILLER_247_1264 ();
 FILLCELL_X32 FILLER_247_1296 ();
 FILLCELL_X32 FILLER_247_1328 ();
 FILLCELL_X32 FILLER_247_1360 ();
 FILLCELL_X32 FILLER_247_1392 ();
 FILLCELL_X32 FILLER_247_1424 ();
 FILLCELL_X32 FILLER_247_1456 ();
 FILLCELL_X32 FILLER_247_1488 ();
 FILLCELL_X32 FILLER_247_1520 ();
 FILLCELL_X32 FILLER_247_1552 ();
 FILLCELL_X32 FILLER_247_1584 ();
 FILLCELL_X32 FILLER_247_1616 ();
 FILLCELL_X32 FILLER_247_1648 ();
 FILLCELL_X32 FILLER_247_1680 ();
 FILLCELL_X32 FILLER_247_1712 ();
 FILLCELL_X32 FILLER_247_1744 ();
 FILLCELL_X32 FILLER_247_1776 ();
 FILLCELL_X32 FILLER_247_1808 ();
 FILLCELL_X32 FILLER_247_1840 ();
 FILLCELL_X16 FILLER_247_1872 ();
 FILLCELL_X8 FILLER_247_1888 ();
 FILLCELL_X32 FILLER_248_1 ();
 FILLCELL_X32 FILLER_248_33 ();
 FILLCELL_X32 FILLER_248_65 ();
 FILLCELL_X32 FILLER_248_97 ();
 FILLCELL_X32 FILLER_248_129 ();
 FILLCELL_X32 FILLER_248_161 ();
 FILLCELL_X32 FILLER_248_193 ();
 FILLCELL_X32 FILLER_248_225 ();
 FILLCELL_X32 FILLER_248_257 ();
 FILLCELL_X32 FILLER_248_289 ();
 FILLCELL_X32 FILLER_248_321 ();
 FILLCELL_X32 FILLER_248_353 ();
 FILLCELL_X32 FILLER_248_385 ();
 FILLCELL_X32 FILLER_248_417 ();
 FILLCELL_X32 FILLER_248_449 ();
 FILLCELL_X32 FILLER_248_481 ();
 FILLCELL_X32 FILLER_248_513 ();
 FILLCELL_X32 FILLER_248_545 ();
 FILLCELL_X32 FILLER_248_577 ();
 FILLCELL_X16 FILLER_248_609 ();
 FILLCELL_X4 FILLER_248_625 ();
 FILLCELL_X2 FILLER_248_629 ();
 FILLCELL_X32 FILLER_248_632 ();
 FILLCELL_X32 FILLER_248_664 ();
 FILLCELL_X32 FILLER_248_696 ();
 FILLCELL_X32 FILLER_248_728 ();
 FILLCELL_X32 FILLER_248_760 ();
 FILLCELL_X32 FILLER_248_792 ();
 FILLCELL_X32 FILLER_248_824 ();
 FILLCELL_X32 FILLER_248_856 ();
 FILLCELL_X32 FILLER_248_888 ();
 FILLCELL_X32 FILLER_248_920 ();
 FILLCELL_X32 FILLER_248_952 ();
 FILLCELL_X32 FILLER_248_984 ();
 FILLCELL_X32 FILLER_248_1016 ();
 FILLCELL_X32 FILLER_248_1048 ();
 FILLCELL_X32 FILLER_248_1080 ();
 FILLCELL_X32 FILLER_248_1112 ();
 FILLCELL_X32 FILLER_248_1144 ();
 FILLCELL_X32 FILLER_248_1176 ();
 FILLCELL_X32 FILLER_248_1208 ();
 FILLCELL_X32 FILLER_248_1240 ();
 FILLCELL_X32 FILLER_248_1272 ();
 FILLCELL_X32 FILLER_248_1304 ();
 FILLCELL_X32 FILLER_248_1336 ();
 FILLCELL_X32 FILLER_248_1368 ();
 FILLCELL_X32 FILLER_248_1400 ();
 FILLCELL_X32 FILLER_248_1432 ();
 FILLCELL_X32 FILLER_248_1464 ();
 FILLCELL_X32 FILLER_248_1496 ();
 FILLCELL_X32 FILLER_248_1528 ();
 FILLCELL_X32 FILLER_248_1560 ();
 FILLCELL_X32 FILLER_248_1592 ();
 FILLCELL_X32 FILLER_248_1624 ();
 FILLCELL_X32 FILLER_248_1656 ();
 FILLCELL_X32 FILLER_248_1688 ();
 FILLCELL_X32 FILLER_248_1720 ();
 FILLCELL_X32 FILLER_248_1752 ();
 FILLCELL_X32 FILLER_248_1784 ();
 FILLCELL_X32 FILLER_248_1816 ();
 FILLCELL_X32 FILLER_248_1848 ();
 FILLCELL_X8 FILLER_248_1880 ();
 FILLCELL_X4 FILLER_248_1888 ();
 FILLCELL_X2 FILLER_248_1892 ();
 FILLCELL_X1 FILLER_248_1895 ();
 FILLCELL_X32 FILLER_249_1 ();
 FILLCELL_X32 FILLER_249_33 ();
 FILLCELL_X32 FILLER_249_65 ();
 FILLCELL_X32 FILLER_249_97 ();
 FILLCELL_X32 FILLER_249_129 ();
 FILLCELL_X32 FILLER_249_161 ();
 FILLCELL_X32 FILLER_249_193 ();
 FILLCELL_X32 FILLER_249_225 ();
 FILLCELL_X32 FILLER_249_257 ();
 FILLCELL_X32 FILLER_249_289 ();
 FILLCELL_X32 FILLER_249_321 ();
 FILLCELL_X32 FILLER_249_353 ();
 FILLCELL_X32 FILLER_249_385 ();
 FILLCELL_X32 FILLER_249_417 ();
 FILLCELL_X32 FILLER_249_449 ();
 FILLCELL_X32 FILLER_249_481 ();
 FILLCELL_X32 FILLER_249_513 ();
 FILLCELL_X32 FILLER_249_545 ();
 FILLCELL_X32 FILLER_249_577 ();
 FILLCELL_X32 FILLER_249_609 ();
 FILLCELL_X32 FILLER_249_641 ();
 FILLCELL_X32 FILLER_249_673 ();
 FILLCELL_X32 FILLER_249_705 ();
 FILLCELL_X32 FILLER_249_737 ();
 FILLCELL_X32 FILLER_249_769 ();
 FILLCELL_X32 FILLER_249_801 ();
 FILLCELL_X32 FILLER_249_833 ();
 FILLCELL_X32 FILLER_249_865 ();
 FILLCELL_X32 FILLER_249_897 ();
 FILLCELL_X32 FILLER_249_929 ();
 FILLCELL_X32 FILLER_249_961 ();
 FILLCELL_X32 FILLER_249_993 ();
 FILLCELL_X32 FILLER_249_1025 ();
 FILLCELL_X32 FILLER_249_1057 ();
 FILLCELL_X32 FILLER_249_1089 ();
 FILLCELL_X32 FILLER_249_1121 ();
 FILLCELL_X32 FILLER_249_1153 ();
 FILLCELL_X32 FILLER_249_1185 ();
 FILLCELL_X32 FILLER_249_1217 ();
 FILLCELL_X8 FILLER_249_1249 ();
 FILLCELL_X4 FILLER_249_1257 ();
 FILLCELL_X2 FILLER_249_1261 ();
 FILLCELL_X32 FILLER_249_1264 ();
 FILLCELL_X32 FILLER_249_1296 ();
 FILLCELL_X32 FILLER_249_1328 ();
 FILLCELL_X32 FILLER_249_1360 ();
 FILLCELL_X32 FILLER_249_1392 ();
 FILLCELL_X32 FILLER_249_1424 ();
 FILLCELL_X32 FILLER_249_1456 ();
 FILLCELL_X32 FILLER_249_1488 ();
 FILLCELL_X32 FILLER_249_1520 ();
 FILLCELL_X32 FILLER_249_1552 ();
 FILLCELL_X32 FILLER_249_1584 ();
 FILLCELL_X32 FILLER_249_1616 ();
 FILLCELL_X32 FILLER_249_1648 ();
 FILLCELL_X32 FILLER_249_1680 ();
 FILLCELL_X32 FILLER_249_1712 ();
 FILLCELL_X32 FILLER_249_1744 ();
 FILLCELL_X32 FILLER_249_1776 ();
 FILLCELL_X32 FILLER_249_1808 ();
 FILLCELL_X32 FILLER_249_1840 ();
 FILLCELL_X16 FILLER_249_1872 ();
 FILLCELL_X8 FILLER_249_1888 ();
 FILLCELL_X32 FILLER_250_1 ();
 FILLCELL_X32 FILLER_250_33 ();
 FILLCELL_X32 FILLER_250_65 ();
 FILLCELL_X32 FILLER_250_97 ();
 FILLCELL_X32 FILLER_250_129 ();
 FILLCELL_X32 FILLER_250_161 ();
 FILLCELL_X32 FILLER_250_193 ();
 FILLCELL_X32 FILLER_250_225 ();
 FILLCELL_X32 FILLER_250_257 ();
 FILLCELL_X32 FILLER_250_289 ();
 FILLCELL_X32 FILLER_250_321 ();
 FILLCELL_X32 FILLER_250_353 ();
 FILLCELL_X32 FILLER_250_385 ();
 FILLCELL_X32 FILLER_250_417 ();
 FILLCELL_X32 FILLER_250_449 ();
 FILLCELL_X32 FILLER_250_481 ();
 FILLCELL_X32 FILLER_250_513 ();
 FILLCELL_X32 FILLER_250_545 ();
 FILLCELL_X32 FILLER_250_577 ();
 FILLCELL_X16 FILLER_250_609 ();
 FILLCELL_X4 FILLER_250_625 ();
 FILLCELL_X2 FILLER_250_629 ();
 FILLCELL_X32 FILLER_250_632 ();
 FILLCELL_X32 FILLER_250_664 ();
 FILLCELL_X32 FILLER_250_696 ();
 FILLCELL_X32 FILLER_250_728 ();
 FILLCELL_X32 FILLER_250_760 ();
 FILLCELL_X32 FILLER_250_792 ();
 FILLCELL_X32 FILLER_250_824 ();
 FILLCELL_X32 FILLER_250_856 ();
 FILLCELL_X32 FILLER_250_888 ();
 FILLCELL_X32 FILLER_250_920 ();
 FILLCELL_X32 FILLER_250_952 ();
 FILLCELL_X32 FILLER_250_984 ();
 FILLCELL_X32 FILLER_250_1016 ();
 FILLCELL_X32 FILLER_250_1048 ();
 FILLCELL_X32 FILLER_250_1080 ();
 FILLCELL_X32 FILLER_250_1112 ();
 FILLCELL_X32 FILLER_250_1144 ();
 FILLCELL_X32 FILLER_250_1176 ();
 FILLCELL_X32 FILLER_250_1208 ();
 FILLCELL_X32 FILLER_250_1240 ();
 FILLCELL_X32 FILLER_250_1272 ();
 FILLCELL_X32 FILLER_250_1304 ();
 FILLCELL_X32 FILLER_250_1336 ();
 FILLCELL_X32 FILLER_250_1368 ();
 FILLCELL_X32 FILLER_250_1400 ();
 FILLCELL_X32 FILLER_250_1432 ();
 FILLCELL_X32 FILLER_250_1464 ();
 FILLCELL_X32 FILLER_250_1496 ();
 FILLCELL_X32 FILLER_250_1528 ();
 FILLCELL_X32 FILLER_250_1560 ();
 FILLCELL_X32 FILLER_250_1592 ();
 FILLCELL_X32 FILLER_250_1624 ();
 FILLCELL_X32 FILLER_250_1656 ();
 FILLCELL_X32 FILLER_250_1688 ();
 FILLCELL_X32 FILLER_250_1720 ();
 FILLCELL_X32 FILLER_250_1752 ();
 FILLCELL_X32 FILLER_250_1784 ();
 FILLCELL_X32 FILLER_250_1816 ();
 FILLCELL_X32 FILLER_250_1848 ();
 FILLCELL_X8 FILLER_250_1880 ();
 FILLCELL_X4 FILLER_250_1888 ();
 FILLCELL_X2 FILLER_250_1892 ();
 FILLCELL_X1 FILLER_250_1895 ();
 FILLCELL_X32 FILLER_251_1 ();
 FILLCELL_X32 FILLER_251_33 ();
 FILLCELL_X32 FILLER_251_65 ();
 FILLCELL_X32 FILLER_251_97 ();
 FILLCELL_X32 FILLER_251_129 ();
 FILLCELL_X32 FILLER_251_161 ();
 FILLCELL_X32 FILLER_251_193 ();
 FILLCELL_X32 FILLER_251_225 ();
 FILLCELL_X32 FILLER_251_257 ();
 FILLCELL_X32 FILLER_251_289 ();
 FILLCELL_X32 FILLER_251_321 ();
 FILLCELL_X32 FILLER_251_353 ();
 FILLCELL_X32 FILLER_251_385 ();
 FILLCELL_X32 FILLER_251_417 ();
 FILLCELL_X32 FILLER_251_449 ();
 FILLCELL_X32 FILLER_251_481 ();
 FILLCELL_X32 FILLER_251_513 ();
 FILLCELL_X32 FILLER_251_545 ();
 FILLCELL_X32 FILLER_251_577 ();
 FILLCELL_X32 FILLER_251_609 ();
 FILLCELL_X32 FILLER_251_641 ();
 FILLCELL_X32 FILLER_251_673 ();
 FILLCELL_X32 FILLER_251_705 ();
 FILLCELL_X32 FILLER_251_737 ();
 FILLCELL_X32 FILLER_251_769 ();
 FILLCELL_X32 FILLER_251_801 ();
 FILLCELL_X32 FILLER_251_833 ();
 FILLCELL_X32 FILLER_251_865 ();
 FILLCELL_X32 FILLER_251_897 ();
 FILLCELL_X32 FILLER_251_929 ();
 FILLCELL_X32 FILLER_251_961 ();
 FILLCELL_X32 FILLER_251_993 ();
 FILLCELL_X32 FILLER_251_1025 ();
 FILLCELL_X32 FILLER_251_1057 ();
 FILLCELL_X32 FILLER_251_1089 ();
 FILLCELL_X32 FILLER_251_1121 ();
 FILLCELL_X32 FILLER_251_1153 ();
 FILLCELL_X32 FILLER_251_1185 ();
 FILLCELL_X32 FILLER_251_1217 ();
 FILLCELL_X8 FILLER_251_1249 ();
 FILLCELL_X4 FILLER_251_1257 ();
 FILLCELL_X2 FILLER_251_1261 ();
 FILLCELL_X32 FILLER_251_1264 ();
 FILLCELL_X32 FILLER_251_1296 ();
 FILLCELL_X32 FILLER_251_1328 ();
 FILLCELL_X32 FILLER_251_1360 ();
 FILLCELL_X32 FILLER_251_1392 ();
 FILLCELL_X32 FILLER_251_1424 ();
 FILLCELL_X32 FILLER_251_1456 ();
 FILLCELL_X32 FILLER_251_1488 ();
 FILLCELL_X32 FILLER_251_1520 ();
 FILLCELL_X32 FILLER_251_1552 ();
 FILLCELL_X32 FILLER_251_1584 ();
 FILLCELL_X32 FILLER_251_1616 ();
 FILLCELL_X32 FILLER_251_1648 ();
 FILLCELL_X32 FILLER_251_1680 ();
 FILLCELL_X32 FILLER_251_1712 ();
 FILLCELL_X32 FILLER_251_1744 ();
 FILLCELL_X32 FILLER_251_1776 ();
 FILLCELL_X32 FILLER_251_1808 ();
 FILLCELL_X32 FILLER_251_1840 ();
 FILLCELL_X16 FILLER_251_1872 ();
 FILLCELL_X8 FILLER_251_1888 ();
 FILLCELL_X32 FILLER_252_1 ();
 FILLCELL_X32 FILLER_252_33 ();
 FILLCELL_X32 FILLER_252_65 ();
 FILLCELL_X32 FILLER_252_97 ();
 FILLCELL_X32 FILLER_252_129 ();
 FILLCELL_X32 FILLER_252_161 ();
 FILLCELL_X32 FILLER_252_193 ();
 FILLCELL_X32 FILLER_252_225 ();
 FILLCELL_X32 FILLER_252_257 ();
 FILLCELL_X32 FILLER_252_289 ();
 FILLCELL_X32 FILLER_252_321 ();
 FILLCELL_X32 FILLER_252_353 ();
 FILLCELL_X32 FILLER_252_385 ();
 FILLCELL_X32 FILLER_252_417 ();
 FILLCELL_X32 FILLER_252_449 ();
 FILLCELL_X32 FILLER_252_481 ();
 FILLCELL_X32 FILLER_252_513 ();
 FILLCELL_X32 FILLER_252_545 ();
 FILLCELL_X32 FILLER_252_577 ();
 FILLCELL_X16 FILLER_252_609 ();
 FILLCELL_X4 FILLER_252_625 ();
 FILLCELL_X2 FILLER_252_629 ();
 FILLCELL_X32 FILLER_252_632 ();
 FILLCELL_X32 FILLER_252_664 ();
 FILLCELL_X32 FILLER_252_696 ();
 FILLCELL_X32 FILLER_252_728 ();
 FILLCELL_X32 FILLER_252_760 ();
 FILLCELL_X32 FILLER_252_792 ();
 FILLCELL_X32 FILLER_252_824 ();
 FILLCELL_X32 FILLER_252_856 ();
 FILLCELL_X32 FILLER_252_888 ();
 FILLCELL_X32 FILLER_252_920 ();
 FILLCELL_X32 FILLER_252_952 ();
 FILLCELL_X32 FILLER_252_984 ();
 FILLCELL_X32 FILLER_252_1016 ();
 FILLCELL_X32 FILLER_252_1048 ();
 FILLCELL_X32 FILLER_252_1080 ();
 FILLCELL_X32 FILLER_252_1112 ();
 FILLCELL_X32 FILLER_252_1144 ();
 FILLCELL_X32 FILLER_252_1176 ();
 FILLCELL_X32 FILLER_252_1208 ();
 FILLCELL_X32 FILLER_252_1240 ();
 FILLCELL_X32 FILLER_252_1272 ();
 FILLCELL_X32 FILLER_252_1304 ();
 FILLCELL_X32 FILLER_252_1336 ();
 FILLCELL_X32 FILLER_252_1368 ();
 FILLCELL_X32 FILLER_252_1400 ();
 FILLCELL_X32 FILLER_252_1432 ();
 FILLCELL_X32 FILLER_252_1464 ();
 FILLCELL_X32 FILLER_252_1496 ();
 FILLCELL_X32 FILLER_252_1528 ();
 FILLCELL_X32 FILLER_252_1560 ();
 FILLCELL_X32 FILLER_252_1592 ();
 FILLCELL_X32 FILLER_252_1624 ();
 FILLCELL_X32 FILLER_252_1656 ();
 FILLCELL_X32 FILLER_252_1688 ();
 FILLCELL_X32 FILLER_252_1720 ();
 FILLCELL_X32 FILLER_252_1752 ();
 FILLCELL_X32 FILLER_252_1784 ();
 FILLCELL_X32 FILLER_252_1816 ();
 FILLCELL_X32 FILLER_252_1848 ();
 FILLCELL_X8 FILLER_252_1880 ();
 FILLCELL_X4 FILLER_252_1888 ();
 FILLCELL_X2 FILLER_252_1892 ();
 FILLCELL_X1 FILLER_252_1895 ();
 FILLCELL_X32 FILLER_253_1 ();
 FILLCELL_X32 FILLER_253_33 ();
 FILLCELL_X32 FILLER_253_65 ();
 FILLCELL_X32 FILLER_253_97 ();
 FILLCELL_X32 FILLER_253_129 ();
 FILLCELL_X32 FILLER_253_161 ();
 FILLCELL_X32 FILLER_253_193 ();
 FILLCELL_X32 FILLER_253_225 ();
 FILLCELL_X32 FILLER_253_257 ();
 FILLCELL_X32 FILLER_253_289 ();
 FILLCELL_X32 FILLER_253_321 ();
 FILLCELL_X32 FILLER_253_353 ();
 FILLCELL_X32 FILLER_253_385 ();
 FILLCELL_X32 FILLER_253_417 ();
 FILLCELL_X32 FILLER_253_449 ();
 FILLCELL_X32 FILLER_253_481 ();
 FILLCELL_X32 FILLER_253_513 ();
 FILLCELL_X32 FILLER_253_545 ();
 FILLCELL_X32 FILLER_253_577 ();
 FILLCELL_X32 FILLER_253_609 ();
 FILLCELL_X32 FILLER_253_641 ();
 FILLCELL_X32 FILLER_253_673 ();
 FILLCELL_X32 FILLER_253_705 ();
 FILLCELL_X32 FILLER_253_737 ();
 FILLCELL_X32 FILLER_253_769 ();
 FILLCELL_X32 FILLER_253_801 ();
 FILLCELL_X32 FILLER_253_833 ();
 FILLCELL_X32 FILLER_253_865 ();
 FILLCELL_X32 FILLER_253_897 ();
 FILLCELL_X32 FILLER_253_929 ();
 FILLCELL_X32 FILLER_253_961 ();
 FILLCELL_X32 FILLER_253_993 ();
 FILLCELL_X32 FILLER_253_1025 ();
 FILLCELL_X32 FILLER_253_1057 ();
 FILLCELL_X32 FILLER_253_1089 ();
 FILLCELL_X32 FILLER_253_1121 ();
 FILLCELL_X32 FILLER_253_1153 ();
 FILLCELL_X32 FILLER_253_1185 ();
 FILLCELL_X32 FILLER_253_1217 ();
 FILLCELL_X8 FILLER_253_1249 ();
 FILLCELL_X4 FILLER_253_1257 ();
 FILLCELL_X2 FILLER_253_1261 ();
 FILLCELL_X32 FILLER_253_1264 ();
 FILLCELL_X32 FILLER_253_1296 ();
 FILLCELL_X32 FILLER_253_1328 ();
 FILLCELL_X32 FILLER_253_1360 ();
 FILLCELL_X32 FILLER_253_1392 ();
 FILLCELL_X32 FILLER_253_1424 ();
 FILLCELL_X32 FILLER_253_1456 ();
 FILLCELL_X32 FILLER_253_1488 ();
 FILLCELL_X32 FILLER_253_1520 ();
 FILLCELL_X32 FILLER_253_1552 ();
 FILLCELL_X32 FILLER_253_1584 ();
 FILLCELL_X32 FILLER_253_1616 ();
 FILLCELL_X32 FILLER_253_1648 ();
 FILLCELL_X32 FILLER_253_1680 ();
 FILLCELL_X32 FILLER_253_1712 ();
 FILLCELL_X32 FILLER_253_1744 ();
 FILLCELL_X32 FILLER_253_1776 ();
 FILLCELL_X32 FILLER_253_1808 ();
 FILLCELL_X32 FILLER_253_1840 ();
 FILLCELL_X16 FILLER_253_1872 ();
 FILLCELL_X8 FILLER_253_1888 ();
 FILLCELL_X32 FILLER_254_1 ();
 FILLCELL_X32 FILLER_254_33 ();
 FILLCELL_X32 FILLER_254_65 ();
 FILLCELL_X32 FILLER_254_97 ();
 FILLCELL_X32 FILLER_254_129 ();
 FILLCELL_X32 FILLER_254_161 ();
 FILLCELL_X32 FILLER_254_193 ();
 FILLCELL_X32 FILLER_254_225 ();
 FILLCELL_X32 FILLER_254_257 ();
 FILLCELL_X32 FILLER_254_289 ();
 FILLCELL_X32 FILLER_254_321 ();
 FILLCELL_X32 FILLER_254_353 ();
 FILLCELL_X32 FILLER_254_385 ();
 FILLCELL_X32 FILLER_254_417 ();
 FILLCELL_X32 FILLER_254_449 ();
 FILLCELL_X32 FILLER_254_481 ();
 FILLCELL_X32 FILLER_254_513 ();
 FILLCELL_X32 FILLER_254_545 ();
 FILLCELL_X32 FILLER_254_577 ();
 FILLCELL_X16 FILLER_254_609 ();
 FILLCELL_X4 FILLER_254_625 ();
 FILLCELL_X2 FILLER_254_629 ();
 FILLCELL_X32 FILLER_254_632 ();
 FILLCELL_X32 FILLER_254_664 ();
 FILLCELL_X32 FILLER_254_696 ();
 FILLCELL_X32 FILLER_254_728 ();
 FILLCELL_X32 FILLER_254_760 ();
 FILLCELL_X32 FILLER_254_792 ();
 FILLCELL_X32 FILLER_254_824 ();
 FILLCELL_X32 FILLER_254_856 ();
 FILLCELL_X32 FILLER_254_888 ();
 FILLCELL_X32 FILLER_254_920 ();
 FILLCELL_X32 FILLER_254_952 ();
 FILLCELL_X32 FILLER_254_984 ();
 FILLCELL_X32 FILLER_254_1016 ();
 FILLCELL_X32 FILLER_254_1048 ();
 FILLCELL_X32 FILLER_254_1080 ();
 FILLCELL_X32 FILLER_254_1112 ();
 FILLCELL_X32 FILLER_254_1144 ();
 FILLCELL_X32 FILLER_254_1176 ();
 FILLCELL_X32 FILLER_254_1208 ();
 FILLCELL_X32 FILLER_254_1240 ();
 FILLCELL_X32 FILLER_254_1272 ();
 FILLCELL_X32 FILLER_254_1304 ();
 FILLCELL_X32 FILLER_254_1336 ();
 FILLCELL_X32 FILLER_254_1368 ();
 FILLCELL_X32 FILLER_254_1400 ();
 FILLCELL_X32 FILLER_254_1432 ();
 FILLCELL_X32 FILLER_254_1464 ();
 FILLCELL_X32 FILLER_254_1496 ();
 FILLCELL_X32 FILLER_254_1528 ();
 FILLCELL_X32 FILLER_254_1560 ();
 FILLCELL_X32 FILLER_254_1592 ();
 FILLCELL_X32 FILLER_254_1624 ();
 FILLCELL_X32 FILLER_254_1656 ();
 FILLCELL_X32 FILLER_254_1688 ();
 FILLCELL_X32 FILLER_254_1720 ();
 FILLCELL_X32 FILLER_254_1752 ();
 FILLCELL_X32 FILLER_254_1784 ();
 FILLCELL_X32 FILLER_254_1816 ();
 FILLCELL_X32 FILLER_254_1848 ();
 FILLCELL_X8 FILLER_254_1880 ();
 FILLCELL_X4 FILLER_254_1888 ();
 FILLCELL_X2 FILLER_254_1892 ();
 FILLCELL_X1 FILLER_254_1895 ();
 FILLCELL_X32 FILLER_255_1 ();
 FILLCELL_X32 FILLER_255_33 ();
 FILLCELL_X32 FILLER_255_65 ();
 FILLCELL_X32 FILLER_255_97 ();
 FILLCELL_X32 FILLER_255_129 ();
 FILLCELL_X32 FILLER_255_161 ();
 FILLCELL_X32 FILLER_255_193 ();
 FILLCELL_X32 FILLER_255_225 ();
 FILLCELL_X32 FILLER_255_257 ();
 FILLCELL_X32 FILLER_255_289 ();
 FILLCELL_X32 FILLER_255_321 ();
 FILLCELL_X32 FILLER_255_353 ();
 FILLCELL_X32 FILLER_255_385 ();
 FILLCELL_X32 FILLER_255_417 ();
 FILLCELL_X32 FILLER_255_449 ();
 FILLCELL_X32 FILLER_255_481 ();
 FILLCELL_X32 FILLER_255_513 ();
 FILLCELL_X32 FILLER_255_545 ();
 FILLCELL_X32 FILLER_255_577 ();
 FILLCELL_X32 FILLER_255_609 ();
 FILLCELL_X32 FILLER_255_641 ();
 FILLCELL_X32 FILLER_255_673 ();
 FILLCELL_X32 FILLER_255_705 ();
 FILLCELL_X32 FILLER_255_737 ();
 FILLCELL_X32 FILLER_255_769 ();
 FILLCELL_X32 FILLER_255_801 ();
 FILLCELL_X32 FILLER_255_833 ();
 FILLCELL_X32 FILLER_255_865 ();
 FILLCELL_X32 FILLER_255_897 ();
 FILLCELL_X32 FILLER_255_929 ();
 FILLCELL_X32 FILLER_255_961 ();
 FILLCELL_X32 FILLER_255_993 ();
 FILLCELL_X16 FILLER_255_1025 ();
 FILLCELL_X8 FILLER_255_1041 ();
 FILLCELL_X4 FILLER_255_1049 ();
 FILLCELL_X1 FILLER_255_1053 ();
 FILLCELL_X32 FILLER_255_1058 ();
 FILLCELL_X32 FILLER_255_1090 ();
 FILLCELL_X32 FILLER_255_1122 ();
 FILLCELL_X32 FILLER_255_1154 ();
 FILLCELL_X32 FILLER_255_1186 ();
 FILLCELL_X32 FILLER_255_1218 ();
 FILLCELL_X8 FILLER_255_1250 ();
 FILLCELL_X4 FILLER_255_1258 ();
 FILLCELL_X1 FILLER_255_1262 ();
 FILLCELL_X32 FILLER_255_1264 ();
 FILLCELL_X32 FILLER_255_1296 ();
 FILLCELL_X32 FILLER_255_1328 ();
 FILLCELL_X32 FILLER_255_1360 ();
 FILLCELL_X32 FILLER_255_1392 ();
 FILLCELL_X32 FILLER_255_1424 ();
 FILLCELL_X32 FILLER_255_1456 ();
 FILLCELL_X32 FILLER_255_1488 ();
 FILLCELL_X32 FILLER_255_1520 ();
 FILLCELL_X32 FILLER_255_1552 ();
 FILLCELL_X32 FILLER_255_1584 ();
 FILLCELL_X32 FILLER_255_1616 ();
 FILLCELL_X32 FILLER_255_1648 ();
 FILLCELL_X32 FILLER_255_1680 ();
 FILLCELL_X32 FILLER_255_1712 ();
 FILLCELL_X32 FILLER_255_1744 ();
 FILLCELL_X32 FILLER_255_1776 ();
 FILLCELL_X32 FILLER_255_1808 ();
 FILLCELL_X32 FILLER_255_1840 ();
 FILLCELL_X16 FILLER_255_1872 ();
 FILLCELL_X8 FILLER_255_1888 ();
 FILLCELL_X32 FILLER_256_1 ();
 FILLCELL_X32 FILLER_256_33 ();
 FILLCELL_X32 FILLER_256_65 ();
 FILLCELL_X32 FILLER_256_97 ();
 FILLCELL_X32 FILLER_256_129 ();
 FILLCELL_X32 FILLER_256_161 ();
 FILLCELL_X32 FILLER_256_193 ();
 FILLCELL_X32 FILLER_256_225 ();
 FILLCELL_X32 FILLER_256_257 ();
 FILLCELL_X32 FILLER_256_289 ();
 FILLCELL_X32 FILLER_256_321 ();
 FILLCELL_X32 FILLER_256_353 ();
 FILLCELL_X32 FILLER_256_385 ();
 FILLCELL_X32 FILLER_256_417 ();
 FILLCELL_X32 FILLER_256_449 ();
 FILLCELL_X32 FILLER_256_481 ();
 FILLCELL_X32 FILLER_256_513 ();
 FILLCELL_X32 FILLER_256_545 ();
 FILLCELL_X32 FILLER_256_577 ();
 FILLCELL_X16 FILLER_256_609 ();
 FILLCELL_X4 FILLER_256_625 ();
 FILLCELL_X2 FILLER_256_629 ();
 FILLCELL_X32 FILLER_256_632 ();
 FILLCELL_X32 FILLER_256_664 ();
 FILLCELL_X32 FILLER_256_696 ();
 FILLCELL_X32 FILLER_256_728 ();
 FILLCELL_X32 FILLER_256_760 ();
 FILLCELL_X32 FILLER_256_792 ();
 FILLCELL_X32 FILLER_256_824 ();
 FILLCELL_X32 FILLER_256_856 ();
 FILLCELL_X32 FILLER_256_888 ();
 FILLCELL_X8 FILLER_256_920 ();
 FILLCELL_X4 FILLER_256_928 ();
 FILLCELL_X16 FILLER_256_936 ();
 FILLCELL_X4 FILLER_256_952 ();
 FILLCELL_X2 FILLER_256_956 ();
 FILLCELL_X32 FILLER_256_961 ();
 FILLCELL_X32 FILLER_256_993 ();
 FILLCELL_X8 FILLER_256_1025 ();
 FILLCELL_X2 FILLER_256_1033 ();
 FILLCELL_X1 FILLER_256_1035 ();
 FILLCELL_X8 FILLER_256_1039 ();
 FILLCELL_X4 FILLER_256_1047 ();
 FILLCELL_X32 FILLER_256_1054 ();
 FILLCELL_X32 FILLER_256_1086 ();
 FILLCELL_X32 FILLER_256_1118 ();
 FILLCELL_X32 FILLER_256_1150 ();
 FILLCELL_X32 FILLER_256_1182 ();
 FILLCELL_X32 FILLER_256_1214 ();
 FILLCELL_X16 FILLER_256_1246 ();
 FILLCELL_X32 FILLER_256_1263 ();
 FILLCELL_X32 FILLER_256_1295 ();
 FILLCELL_X32 FILLER_256_1327 ();
 FILLCELL_X32 FILLER_256_1359 ();
 FILLCELL_X32 FILLER_256_1391 ();
 FILLCELL_X32 FILLER_256_1423 ();
 FILLCELL_X32 FILLER_256_1455 ();
 FILLCELL_X32 FILLER_256_1487 ();
 FILLCELL_X32 FILLER_256_1519 ();
 FILLCELL_X32 FILLER_256_1551 ();
 FILLCELL_X32 FILLER_256_1583 ();
 FILLCELL_X32 FILLER_256_1615 ();
 FILLCELL_X32 FILLER_256_1647 ();
 FILLCELL_X32 FILLER_256_1679 ();
 FILLCELL_X32 FILLER_256_1711 ();
 FILLCELL_X32 FILLER_256_1743 ();
 FILLCELL_X32 FILLER_256_1775 ();
 FILLCELL_X32 FILLER_256_1807 ();
 FILLCELL_X32 FILLER_256_1839 ();
 FILLCELL_X16 FILLER_256_1871 ();
 FILLCELL_X4 FILLER_256_1887 ();
 FILLCELL_X2 FILLER_256_1891 ();
 FILLCELL_X2 FILLER_256_1894 ();
endmodule
