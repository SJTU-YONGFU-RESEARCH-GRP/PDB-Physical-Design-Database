module multi_ported_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rst_n,
    data_count,
    rd_data,
    rd_en,
    rd_valid,
    wr_data,
    wr_en,
    wr_ready);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rst_n;
 output [4:0] data_count;
 output [63:0] rd_data;
 input [1:0] rd_en;
 output [1:0] rd_valid;
 input [63:0] wr_data;
 input [1:0] wr_en;
 output [1:0] wr_ready;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \next_count[0] ;
 wire \next_count[1] ;
 wire \next_count[2] ;
 wire \next_count[3] ;
 wire \next_count[4] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;

 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2762_ (.A1(_2116_),
    .A2(_2293_),
    .A3(_2300_),
    .A4(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2763_ (.I0(\mem[12][25] ),
    .I1(\mem[14][25] ),
    .S(_1994_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2764_ (.A1(_2203_),
    .A2(_1968_),
    .A3(_2306_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2765_ (.I(_1786_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2766_ (.A1(_2256_),
    .A2(_1586_),
    .A3(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2767_ (.I(_1803_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2768_ (.I0(\mem[9][25] ),
    .I1(\mem[11][25] ),
    .I2(\mem[13][25] ),
    .I3(\mem[15][25] ),
    .S0(_2079_),
    .S1(_2310_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2769_ (.I(_1376_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2770_ (.I0(_1585_),
    .I1(_1591_),
    .S(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2771_ (.I(_2712_),
    .Z(_2314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2772_ (.I0(\mem[8][25] ),
    .I1(\mem[10][25] ),
    .S(_2314_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2773_ (.A1(_2109_),
    .A2(_2315_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2774_ (.A1(_2030_),
    .A2(_1590_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2775_ (.I0(_2311_),
    .I1(_2313_),
    .I2(_2316_),
    .I3(_2317_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2776_ (.A1(_2133_),
    .A2(_2307_),
    .A3(_2309_),
    .A4(_2318_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2777_ (.A1(_2290_),
    .A2(_2305_),
    .A3(_2319_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2778_ (.A1(net132),
    .A2(_2186_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2779_ (.A1(_2061_),
    .A2(\mem[0][26] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][26] ),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2780_ (.A1(_2063_),
    .A2(\mem[2][26] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][26] ),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2781_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2321_),
    .A4(_2322_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2782_ (.I0(\mem[4][26] ),
    .I1(\mem[6][26] ),
    .S(_2294_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2783_ (.I0(_1596_),
    .I1(_2324_),
    .S(_2296_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2784_ (.I0(\mem[5][26] ),
    .I1(\mem[7][26] ),
    .S(_2013_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2785_ (.I0(_1595_),
    .I1(_2326_),
    .S(_2041_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2786_ (.A1(_2122_),
    .A2(_2325_),
    .B1(_2327_),
    .B2(_2097_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2787_ (.I(_1805_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2788_ (.I0(\mem[0][26] ),
    .I1(\mem[2][26] ),
    .S(_2197_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2789_ (.A1(_2329_),
    .A2(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2790_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1600_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2791_ (.A1(_2331_),
    .A2(_2332_),
    .B(_2251_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2792_ (.A1(_2116_),
    .A2(_2323_),
    .A3(_2328_),
    .A4(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2793_ (.I(_1818_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2794_ (.I0(\mem[12][26] ),
    .I1(\mem[14][26] ),
    .S(_1994_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2795_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2336_),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2796_ (.A1(_2256_),
    .A2(_1598_),
    .A3(_2308_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2797_ (.I0(\mem[9][26] ),
    .I1(\mem[11][26] ),
    .I2(\mem[13][26] ),
    .I3(\mem[15][26] ),
    .S0(_2079_),
    .S1(_2310_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2798_ (.I0(_1597_),
    .I1(_1604_),
    .S(_2312_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2799_ (.I0(\mem[8][26] ),
    .I1(\mem[10][26] ),
    .S(_2314_),
    .Z(_2341_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2800_ (.A1(_2109_),
    .A2(_2341_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2801_ (.A1(_2030_),
    .A2(_1603_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2802_ (.I0(_2339_),
    .I1(_2340_),
    .I2(_2342_),
    .I3(_2343_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2803_ (.A1(_2133_),
    .A2(_2337_),
    .A3(_2338_),
    .A4(_2344_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2804_ (.A1(_2320_),
    .A2(_2334_),
    .A3(_2345_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2805_ (.A1(net133),
    .A2(_2186_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2806_ (.A1(_2061_),
    .A2(\mem[0][27] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][27] ),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2807_ (.A1(_2063_),
    .A2(\mem[2][27] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][27] ),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2808_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2347_),
    .A4(_2348_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2809_ (.I0(\mem[4][27] ),
    .I1(\mem[6][27] ),
    .S(_2294_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2810_ (.I0(_1609_),
    .I1(_2350_),
    .S(_2296_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2811_ (.I0(\mem[5][27] ),
    .I1(\mem[7][27] ),
    .S(_2013_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2812_ (.I0(_1608_),
    .I1(_2352_),
    .S(_2041_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2813_ (.A1(_2122_),
    .A2(_2351_),
    .B1(_2353_),
    .B2(_2097_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2814_ (.I0(\mem[0][27] ),
    .I1(\mem[2][27] ),
    .S(_2197_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2815_ (.A1(_2329_),
    .A2(_2355_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2816_ (.I(_1732_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2817_ (.A1(_2357_),
    .A2(_2019_),
    .A3(_1614_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2818_ (.A1(_2356_),
    .A2(_2358_),
    .B(_2251_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2819_ (.A1(_2116_),
    .A2(_2349_),
    .A3(_2354_),
    .A4(_2359_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2820_ (.I(_1782_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2821_ (.I0(\mem[12][27] ),
    .I1(\mem[14][27] ),
    .S(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2822_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2362_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2823_ (.A1(_2256_),
    .A2(_1611_),
    .A3(_2308_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2824_ (.I0(\mem[9][27] ),
    .I1(\mem[11][27] ),
    .I2(\mem[13][27] ),
    .I3(\mem[15][27] ),
    .S0(_2079_),
    .S1(_2310_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2825_ (.I0(_1610_),
    .I1(_1618_),
    .S(_2312_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2826_ (.I0(\mem[8][27] ),
    .I1(\mem[10][27] ),
    .S(_2314_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2827_ (.A1(_2109_),
    .A2(_2367_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2828_ (.A1(_2030_),
    .A2(_1617_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2829_ (.I(_1534_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2830_ (.I0(_2365_),
    .I1(_2366_),
    .I2(_2368_),
    .I3(_2369_),
    .S0(_2057_),
    .S1(_2370_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2831_ (.A1(_2133_),
    .A2(_2363_),
    .A3(_2364_),
    .A4(_2371_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2832_ (.A1(_2346_),
    .A2(_2360_),
    .A3(_2372_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2833_ (.A1(net135),
    .A2(_2186_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2834_ (.A1(_2061_),
    .A2(\mem[0][28] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][28] ),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2835_ (.A1(_2063_),
    .A2(\mem[2][28] ),
    .A3(_2172_),
    .B1(_2090_),
    .B2(\mem[3][28] ),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2836_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2374_),
    .A4(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2837_ (.I0(\mem[4][28] ),
    .I1(\mem[6][28] ),
    .S(_2294_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2838_ (.I0(_1624_),
    .I1(_2377_),
    .S(_2296_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2839_ (.I0(\mem[5][28] ),
    .I1(\mem[7][28] ),
    .S(_2170_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2840_ (.I0(_1623_),
    .I1(_2379_),
    .S(_2041_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2841_ (.A1(_2122_),
    .A2(_2378_),
    .B1(_2380_),
    .B2(_2097_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2842_ (.I0(\mem[0][28] ),
    .I1(\mem[2][28] ),
    .S(_2197_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2843_ (.A1(_2329_),
    .A2(_2382_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2844_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1628_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2845_ (.A1(_2383_),
    .A2(_2384_),
    .B(_2251_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2846_ (.A1(_2116_),
    .A2(_2376_),
    .A3(_2381_),
    .A4(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2847_ (.I0(\mem[12][28] ),
    .I1(\mem[14][28] ),
    .S(_2361_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2848_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2387_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2849_ (.A1(_2256_),
    .A2(_1626_),
    .A3(_2308_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2850_ (.I0(\mem[9][28] ),
    .I1(\mem[11][28] ),
    .I2(\mem[13][28] ),
    .I3(\mem[15][28] ),
    .S0(_2079_),
    .S1(_2310_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2851_ (.I0(_1625_),
    .I1(_1631_),
    .S(_2312_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2852_ (.I0(\mem[8][28] ),
    .I1(\mem[10][28] ),
    .S(_2314_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2853_ (.A1(_2109_),
    .A2(_2392_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2854_ (.A1(_2152_),
    .A2(_1630_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2855_ (.I0(_2390_),
    .I1(_2391_),
    .I2(_2393_),
    .I3(_2394_),
    .S0(_2057_),
    .S1(_2370_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2856_ (.A1(_2133_),
    .A2(_2388_),
    .A3(_2389_),
    .A4(_2395_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2857_ (.A1(_2373_),
    .A2(_2386_),
    .A3(_2396_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2858_ (.A1(net136),
    .A2(_2186_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2859_ (.A1(_2061_),
    .A2(\mem[0][29] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][29] ),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2860_ (.A1(_2063_),
    .A2(\mem[2][29] ),
    .A3(_2172_),
    .B1(_2090_),
    .B2(\mem[3][29] ),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2861_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2398_),
    .A4(_2399_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2862_ (.I0(\mem[4][29] ),
    .I1(\mem[6][29] ),
    .S(_2294_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2863_ (.I0(_1635_),
    .I1(_2401_),
    .S(_2296_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2864_ (.I0(\mem[5][29] ),
    .I1(\mem[7][29] ),
    .S(_2170_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2865_ (.I0(_1634_),
    .I1(_2403_),
    .S(_1771_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2866_ (.A1(_2122_),
    .A2(_2402_),
    .B1(_2404_),
    .B2(_2097_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2867_ (.I0(\mem[0][29] ),
    .I1(\mem[2][29] ),
    .S(_2197_),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2868_ (.A1(_2329_),
    .A2(_2406_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2869_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1639_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2870_ (.A1(_2407_),
    .A2(_2408_),
    .B(_2251_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2871_ (.A1(_2116_),
    .A2(_2400_),
    .A3(_2405_),
    .A4(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2872_ (.I0(\mem[12][29] ),
    .I1(\mem[14][29] ),
    .S(_2361_),
    .Z(_2411_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2873_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2411_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2874_ (.A1(_2256_),
    .A2(_1637_),
    .A3(_2308_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2875_ (.I0(\mem[9][29] ),
    .I1(\mem[11][29] ),
    .I2(\mem[13][29] ),
    .I3(\mem[15][29] ),
    .S0(_2079_),
    .S1(_2310_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2876_ (.I0(_1636_),
    .I1(_1642_),
    .S(_2312_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2877_ (.I0(\mem[8][29] ),
    .I1(\mem[10][29] ),
    .S(_2314_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2878_ (.A1(_2109_),
    .A2(_2416_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2879_ (.A1(_2152_),
    .A2(_1641_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2880_ (.I0(_2414_),
    .I1(_2415_),
    .I2(_2417_),
    .I3(_2418_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2881_ (.A1(_2133_),
    .A2(_2412_),
    .A3(_2413_),
    .A4(_2419_),
    .Z(_2420_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2882_ (.A1(_2397_),
    .A2(_2410_),
    .A3(_2420_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2883_ (.A1(net106),
    .A2(_2186_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2884_ (.A1(_2162_),
    .A2(\mem[0][2] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][2] ),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2885_ (.A1(_2166_),
    .A2(\mem[2][2] ),
    .A3(_2172_),
    .B1(_2090_),
    .B2(\mem[3][2] ),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2886_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2422_),
    .A4(_2423_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2887_ (.I0(\mem[4][2] ),
    .I1(\mem[6][2] ),
    .S(_2294_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2888_ (.I0(_1646_),
    .I1(_2425_),
    .S(_2296_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2889_ (.I0(\mem[5][2] ),
    .I1(\mem[7][2] ),
    .S(_2170_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2890_ (.I0(_1645_),
    .I1(_2427_),
    .S(_1771_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2891_ (.A1(_2122_),
    .A2(_2426_),
    .B1(_2428_),
    .B2(_2097_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2892_ (.I0(\mem[0][2] ),
    .I1(\mem[2][2] ),
    .S(_2197_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2893_ (.A1(_2329_),
    .A2(_2430_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2894_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1650_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2895_ (.A1(_2431_),
    .A2(_2432_),
    .B(_2251_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2896_ (.A1(_2116_),
    .A2(_2424_),
    .A3(_2429_),
    .A4(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2897_ (.I0(\mem[12][2] ),
    .I1(\mem[14][2] ),
    .S(_2361_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2898_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2435_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2899_ (.A1(_2256_),
    .A2(_1648_),
    .A3(_2308_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2900_ (.I0(\mem[9][2] ),
    .I1(\mem[11][2] ),
    .I2(\mem[13][2] ),
    .I3(\mem[15][2] ),
    .S0(_1800_),
    .S1(_2310_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2901_ (.I0(_1647_),
    .I1(_1653_),
    .S(_2312_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2902_ (.I0(\mem[8][2] ),
    .I1(\mem[10][2] ),
    .S(_2314_),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2903_ (.A1(_2109_),
    .A2(_2440_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2904_ (.A1(_2152_),
    .A2(_1652_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2905_ (.I0(_2438_),
    .I1(_2439_),
    .I2(_2441_),
    .I3(_2442_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2443_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2906_ (.A1(_2133_),
    .A2(_2436_),
    .A3(_2437_),
    .A4(_2443_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2907_ (.A1(_2421_),
    .A2(_2434_),
    .A3(_2444_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2908_ (.A1(net137),
    .A2(_2186_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2909_ (.A1(_2162_),
    .A2(\mem[0][30] ),
    .A3(_2188_),
    .B1(_2164_),
    .B2(\mem[1][30] ),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2910_ (.A1(_2166_),
    .A2(\mem[2][30] ),
    .A3(_2172_),
    .B1(_2167_),
    .B2(\mem[3][30] ),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2911_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2446_),
    .A4(_2447_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2912_ (.I0(\mem[4][30] ),
    .I1(\mem[6][30] ),
    .S(_2294_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2913_ (.I0(_1657_),
    .I1(_2449_),
    .S(_2296_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2914_ (.I0(\mem[5][30] ),
    .I1(\mem[7][30] ),
    .S(_2170_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2915_ (.I0(_1656_),
    .I1(_2451_),
    .S(_1771_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2916_ (.A1(_2122_),
    .A2(_2450_),
    .B1(_2452_),
    .B2(_2178_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2917_ (.I0(\mem[0][30] ),
    .I1(\mem[2][30] ),
    .S(_2197_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2918_ (.A1(_2329_),
    .A2(_2454_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2919_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1661_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2920_ (.A1(_2455_),
    .A2(_2456_),
    .B(_2251_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2921_ (.A1(_2116_),
    .A2(_2448_),
    .A3(_2453_),
    .A4(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2922_ (.I0(\mem[12][30] ),
    .I1(\mem[14][30] ),
    .S(_2361_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2923_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2459_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2924_ (.A1(_2256_),
    .A2(_1659_),
    .A3(_2308_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2925_ (.I0(\mem[9][30] ),
    .I1(\mem[11][30] ),
    .I2(\mem[13][30] ),
    .I3(\mem[15][30] ),
    .S0(_1800_),
    .S1(_2310_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2926_ (.I0(_1658_),
    .I1(_1664_),
    .S(_2312_),
    .Z(_2463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2927_ (.I0(\mem[8][30] ),
    .I1(\mem[10][30] ),
    .S(_2314_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2928_ (.A1(_1826_),
    .A2(_2464_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2929_ (.A1(_2152_),
    .A2(_1663_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2930_ (.I0(_2462_),
    .I1(_2463_),
    .I2(_2465_),
    .I3(_2466_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2931_ (.A1(_2133_),
    .A2(_2460_),
    .A3(_2461_),
    .A4(_2467_),
    .Z(_2468_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2932_ (.A1(_2445_),
    .A2(_2458_),
    .A3(_2468_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2933_ (.A1(net138),
    .A2(_2186_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2934_ (.A1(_2162_),
    .A2(\mem[0][31] ),
    .A3(_2188_),
    .B1(_2164_),
    .B2(\mem[1][31] ),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2935_ (.A1(_2166_),
    .A2(\mem[2][31] ),
    .A3(_2172_),
    .B1(_2167_),
    .B2(\mem[3][31] ),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2936_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2470_),
    .A4(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2937_ (.I0(\mem[4][31] ),
    .I1(\mem[6][31] ),
    .S(_2294_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2938_ (.I0(_1668_),
    .I1(_2473_),
    .S(_2296_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2939_ (.I0(\mem[5][31] ),
    .I1(\mem[7][31] ),
    .S(_2170_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2940_ (.I0(_1667_),
    .I1(_2475_),
    .S(_1771_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2941_ (.A1(_1790_),
    .A2(_2474_),
    .B1(_2476_),
    .B2(_2178_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2942_ (.I0(\mem[0][31] ),
    .I1(\mem[2][31] ),
    .S(_2197_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2943_ (.A1(_2329_),
    .A2(_2478_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2944_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1672_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2945_ (.A1(_2479_),
    .A2(_2480_),
    .B(_2251_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2946_ (.A1(_2144_),
    .A2(_2472_),
    .A3(_2477_),
    .A4(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2947_ (.I0(\mem[12][31] ),
    .I1(\mem[14][31] ),
    .S(_2361_),
    .Z(_2483_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2948_ (.A1(_2203_),
    .A2(_2335_),
    .A3(_2483_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2949_ (.A1(_2256_),
    .A2(_1670_),
    .A3(_2308_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2950_ (.I0(\mem[9][31] ),
    .I1(\mem[11][31] ),
    .I2(\mem[13][31] ),
    .I3(\mem[15][31] ),
    .S0(_1800_),
    .S1(_2310_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2951_ (.I0(_1669_),
    .I1(_1675_),
    .S(_2312_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2952_ (.I0(\mem[8][31] ),
    .I1(\mem[10][31] ),
    .S(_2314_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2953_ (.A1(_1826_),
    .A2(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2954_ (.A1(_2152_),
    .A2(_1674_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2955_ (.I0(_2486_),
    .I1(_2487_),
    .I2(_2489_),
    .I3(_2490_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2956_ (.A1(_1855_),
    .A2(_2484_),
    .A3(_2485_),
    .A4(_2491_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2957_ (.A1(_2469_),
    .A2(_2482_),
    .A3(_2492_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2958_ (.A1(net107),
    .A2(_0611_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2959_ (.A1(_2162_),
    .A2(\mem[0][3] ),
    .A3(_1840_),
    .B1(_2164_),
    .B2(\mem[1][3] ),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2960_ (.A1(_2166_),
    .A2(\mem[2][3] ),
    .A3(_2172_),
    .B1(_2167_),
    .B2(\mem[3][3] ),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2961_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2494_),
    .A4(_2495_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2962_ (.I0(\mem[4][3] ),
    .I1(\mem[6][3] ),
    .S(_2294_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2963_ (.I0(_1679_),
    .I1(_2497_),
    .S(_2296_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2964_ (.I0(\mem[5][3] ),
    .I1(\mem[7][3] ),
    .S(_2170_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2965_ (.I0(_1678_),
    .I1(_2499_),
    .S(_1771_),
    .Z(_2500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2966_ (.A1(_1790_),
    .A2(_2498_),
    .B1(_2500_),
    .B2(_2178_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2967_ (.I0(\mem[0][3] ),
    .I1(\mem[2][3] ),
    .S(_1816_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2968_ (.A1(_2329_),
    .A2(_2502_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2969_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1683_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2970_ (.A1(_2503_),
    .A2(_2504_),
    .B(_2251_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2971_ (.A1(_2144_),
    .A2(_2496_),
    .A3(_2501_),
    .A4(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2972_ (.I0(\mem[12][3] ),
    .I1(\mem[14][3] ),
    .S(_2361_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2973_ (.A1(_1735_),
    .A2(_2335_),
    .A3(_2507_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2974_ (.A1(_2256_),
    .A2(_1681_),
    .A3(_2308_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2975_ (.I0(\mem[9][3] ),
    .I1(\mem[11][3] ),
    .I2(\mem[13][3] ),
    .I3(\mem[15][3] ),
    .S0(_1800_),
    .S1(_2310_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2976_ (.I0(_1680_),
    .I1(_1686_),
    .S(_2312_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2977_ (.I0(\mem[8][3] ),
    .I1(\mem[10][3] ),
    .S(_2314_),
    .Z(_2512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2978_ (.A1(_1826_),
    .A2(_2512_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2979_ (.A1(_2152_),
    .A2(_1685_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2980_ (.I0(_2510_),
    .I1(_2511_),
    .I2(_2513_),
    .I3(_2514_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2981_ (.A1(_1855_),
    .A2(_2508_),
    .A3(_2509_),
    .A4(_2515_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2982_ (.A1(_2493_),
    .A2(_2506_),
    .A3(_2516_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2983_ (.I0(\mem[4][4] ),
    .I1(\mem[6][4] ),
    .S(_2145_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2984_ (.A1(_1736_),
    .A2(_1857_),
    .A3(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2985_ (.A1(_2729_),
    .A2(_1689_),
    .A3(_1820_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2986_ (.A1(_2144_),
    .A2(_2518_),
    .A3(_2519_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2987_ (.I0(\mem[1][4] ),
    .I1(\mem[3][4] ),
    .I2(\mem[5][4] ),
    .I3(\mem[7][4] ),
    .S0(_1801_),
    .S1(_1823_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2988_ (.I0(_1690_),
    .I1(_1694_),
    .S(_1377_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2989_ (.A1(_2182_),
    .A2(_2522_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2990_ (.A1(_0604_),
    .A2(_2521_),
    .B(_2523_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2991_ (.I0(\mem[0][4] ),
    .I1(\mem[2][4] ),
    .S(_2145_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2992_ (.A1(_1695_),
    .A2(_2156_),
    .B1(_2525_),
    .B2(_1849_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2993_ (.I0(_2524_),
    .I1(_2526_),
    .S(_1811_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2994_ (.A1(net108),
    .A2(_2731_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2995_ (.A1(_1391_),
    .A2(\mem[8][4] ),
    .A3(_2163_),
    .B1(_2164_),
    .B2(\mem[9][4] ),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _2996_ (.A1(_0614_),
    .A2(\mem[10][4] ),
    .A3(_0603_),
    .B1(_2167_),
    .B2(\mem[11][4] ),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2997_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2529_),
    .A4(_2530_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2998_ (.I0(\mem[12][4] ),
    .I1(\mem[14][4] ),
    .S(_2174_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2999_ (.I0(_1691_),
    .I1(_2532_),
    .S(_2176_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3000_ (.I0(\mem[13][4] ),
    .I1(\mem[15][4] ),
    .S(_2174_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3001_ (.I0(_1692_),
    .I1(_2534_),
    .S(_2176_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3002_ (.A1(_1790_),
    .A2(_2533_),
    .B1(_2535_),
    .B2(_2178_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3003_ (.I0(\mem[8][4] ),
    .I1(\mem[10][4] ),
    .S(_1783_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3004_ (.A1(_1806_),
    .A2(_2537_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3005_ (.A1(_1378_),
    .A2(_2182_),
    .A3(_1697_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3006_ (.A1(_2538_),
    .A2(_2539_),
    .B(_1760_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3007_ (.A1(_1799_),
    .A2(_2531_),
    .A3(_2536_),
    .A4(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3008_ (.A1(_2520_),
    .A2(_2527_),
    .B(_2528_),
    .C(_2541_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3009_ (.A1(net109),
    .A2(_0611_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3010_ (.A1(_2162_),
    .A2(\mem[0][5] ),
    .A3(_1840_),
    .B1(_2164_),
    .B2(\mem[1][5] ),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3011_ (.A1(_2166_),
    .A2(\mem[2][5] ),
    .A3(_2172_),
    .B1(_2167_),
    .B2(\mem[3][5] ),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3012_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2543_),
    .A4(_2544_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3013_ (.I0(\mem[4][5] ),
    .I1(\mem[6][5] ),
    .S(_2294_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3014_ (.I0(_1701_),
    .I1(_2546_),
    .S(_2296_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3015_ (.I0(\mem[5][5] ),
    .I1(\mem[7][5] ),
    .S(_2170_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3016_ (.I0(_1700_),
    .I1(_2548_),
    .S(_1771_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3017_ (.A1(_1790_),
    .A2(_2547_),
    .B1(_2549_),
    .B2(_2178_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3018_ (.I0(\mem[0][5] ),
    .I1(\mem[2][5] ),
    .S(_1816_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3019_ (.A1(_2329_),
    .A2(_2551_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3020_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1705_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3021_ (.A1(_2552_),
    .A2(_2553_),
    .B(_1760_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3022_ (.A1(_2144_),
    .A2(_2545_),
    .A3(_2550_),
    .A4(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3023_ (.I0(\mem[12][5] ),
    .I1(\mem[14][5] ),
    .S(_2361_),
    .Z(_2556_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3024_ (.A1(_1735_),
    .A2(_2335_),
    .A3(_2556_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3025_ (.A1(_1808_),
    .A2(_1703_),
    .A3(_2308_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3026_ (.I0(\mem[9][5] ),
    .I1(\mem[11][5] ),
    .I2(\mem[13][5] ),
    .I3(\mem[15][5] ),
    .S0(_1800_),
    .S1(_2310_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3027_ (.I0(_1702_),
    .I1(_1708_),
    .S(_2312_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3028_ (.I0(\mem[8][5] ),
    .I1(\mem[10][5] ),
    .S(_2314_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3029_ (.A1(_1826_),
    .A2(_2561_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3030_ (.A1(_2152_),
    .A2(_1707_),
    .Z(_2563_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3031_ (.I0(_2559_),
    .I1(_2560_),
    .I2(_2562_),
    .I3(_2563_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3032_ (.A1(_1855_),
    .A2(_2557_),
    .A3(_2558_),
    .A4(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3033_ (.A1(_2542_),
    .A2(_2555_),
    .A3(_2565_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3034_ (.I0(\mem[4][6] ),
    .I1(\mem[6][6] ),
    .S(_2145_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3035_ (.A1(_1736_),
    .A2(_1857_),
    .A3(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3036_ (.A1(_2729_),
    .A2(_1711_),
    .A3(_1820_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3037_ (.A1(_2144_),
    .A2(_2567_),
    .A3(_2568_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3038_ (.I0(\mem[1][6] ),
    .I1(\mem[3][6] ),
    .I2(\mem[5][6] ),
    .I3(\mem[7][6] ),
    .S0(_1801_),
    .S1(_1823_),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3039_ (.I0(_1712_),
    .I1(_1716_),
    .S(_1377_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3040_ (.A1(_2182_),
    .A2(_2571_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3041_ (.A1(_0604_),
    .A2(_2570_),
    .B(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3042_ (.I0(\mem[0][6] ),
    .I1(\mem[2][6] ),
    .S(_1801_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3043_ (.A1(_1717_),
    .A2(_2156_),
    .B1(_2574_),
    .B2(_1849_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3044_ (.I0(_2573_),
    .I1(_2575_),
    .S(_1811_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3045_ (.A1(net110),
    .A2(_2731_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3046_ (.A1(_1391_),
    .A2(\mem[8][6] ),
    .A3(_2163_),
    .B1(_1773_),
    .B2(\mem[9][6] ),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3047_ (.A1(_0614_),
    .A2(\mem[10][6] ),
    .A3(_0603_),
    .B1(_1762_),
    .B2(\mem[11][6] ),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3048_ (.A1(_2161_),
    .A2(_1768_),
    .A3(_2578_),
    .A4(_2579_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3049_ (.I0(\mem[12][6] ),
    .I1(\mem[14][6] ),
    .S(_2174_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3050_ (.I0(_1713_),
    .I1(_2581_),
    .S(_2176_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3051_ (.I0(\mem[13][6] ),
    .I1(\mem[15][6] ),
    .S(_2174_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3052_ (.I0(_1714_),
    .I1(_2583_),
    .S(_2176_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3053_ (.A1(_1789_),
    .A2(_2582_),
    .B1(_2584_),
    .B2(_1780_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3054_ (.I0(\mem[8][6] ),
    .I1(\mem[10][6] ),
    .S(_1783_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3055_ (.A1(_1806_),
    .A2(_2586_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3056_ (.A1(_1378_),
    .A2(_2182_),
    .A3(_1719_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3057_ (.A1(_2587_),
    .A2(_2588_),
    .B(_1760_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3058_ (.A1(_1799_),
    .A2(_2580_),
    .A3(_2585_),
    .A4(_2589_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3059_ (.A1(_2569_),
    .A2(_2576_),
    .B(_2577_),
    .C(_2590_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3060_ (.A1(net111),
    .A2(_0611_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3061_ (.A1(_2162_),
    .A2(\mem[0][7] ),
    .A3(_1840_),
    .B1(_2164_),
    .B2(\mem[1][7] ),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3062_ (.A1(_2166_),
    .A2(\mem[2][7] ),
    .A3(_2172_),
    .B1(_2167_),
    .B2(\mem[3][7] ),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3063_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2592_),
    .A4(_2593_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3064_ (.I0(\mem[4][7] ),
    .I1(\mem[6][7] ),
    .S(_1791_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3065_ (.I0(_1723_),
    .I1(_2595_),
    .S(_1793_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3066_ (.I0(\mem[5][7] ),
    .I1(\mem[7][7] ),
    .S(_2170_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3067_ (.I0(_1722_),
    .I1(_2597_),
    .S(_1771_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3068_ (.A1(_1790_),
    .A2(_2596_),
    .B1(_2598_),
    .B2(_2178_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3069_ (.I0(\mem[0][7] ),
    .I1(\mem[2][7] ),
    .S(_1816_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3070_ (.A1(_2329_),
    .A2(_2600_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3071_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1727_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3072_ (.A1(_2601_),
    .A2(_2602_),
    .B(_1760_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3073_ (.A1(_2144_),
    .A2(_2594_),
    .A3(_2599_),
    .A4(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3074_ (.I0(\mem[12][7] ),
    .I1(\mem[14][7] ),
    .S(_2361_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3075_ (.A1(_1735_),
    .A2(_2335_),
    .A3(_2605_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3076_ (.A1(_1808_),
    .A2(_1725_),
    .A3(_1786_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3077_ (.I0(\mem[9][7] ),
    .I1(\mem[11][7] ),
    .I2(\mem[13][7] ),
    .I3(\mem[15][7] ),
    .S0(_1800_),
    .S1(_1803_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3078_ (.I0(_1724_),
    .I1(_1730_),
    .S(_1376_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3079_ (.I0(\mem[8][7] ),
    .I1(\mem[10][7] ),
    .S(_1761_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3080_ (.A1(_1826_),
    .A2(_2610_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3081_ (.A1(_2152_),
    .A2(_1729_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3082_ (.I0(_2608_),
    .I1(_2609_),
    .I2(_2611_),
    .I3(_2612_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3083_ (.A1(_1855_),
    .A2(_2606_),
    .A3(_2607_),
    .A4(_2613_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3084_ (.A1(_2591_),
    .A2(_2604_),
    .A3(_2614_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3085_ (.I0(\mem[4][8] ),
    .I1(\mem[6][8] ),
    .S(_2145_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3086_ (.A1(_1736_),
    .A2(_1857_),
    .A3(_2615_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3087_ (.A1(_2729_),
    .A2(_1737_),
    .A3(_1820_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3088_ (.A1(_1835_),
    .A2(_2616_),
    .A3(_2617_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3089_ (.I0(\mem[1][8] ),
    .I1(\mem[3][8] ),
    .I2(\mem[5][8] ),
    .I3(\mem[7][8] ),
    .S0(_1801_),
    .S1(_1823_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3090_ (.I0(_1738_),
    .I1(_1742_),
    .S(_1377_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3091_ (.A1(_2182_),
    .A2(_2620_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3092_ (.A1(_0604_),
    .A2(_2619_),
    .B(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3093_ (.I0(\mem[0][8] ),
    .I1(\mem[2][8] ),
    .S(_1801_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3094_ (.A1(_1743_),
    .A2(_2156_),
    .B1(_2623_),
    .B2(_1849_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3095_ (.I0(_2622_),
    .I1(_2624_),
    .S(_1811_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3096_ (.A1(net113),
    .A2(_2731_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3097_ (.A1(_1391_),
    .A2(\mem[8][8] ),
    .A3(_2163_),
    .B1(_1773_),
    .B2(\mem[9][8] ),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3098_ (.A1(_0614_),
    .A2(\mem[10][8] ),
    .A3(_0603_),
    .B1(_1762_),
    .B2(\mem[11][8] ),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3099_ (.A1(_1810_),
    .A2(_1768_),
    .A3(_2627_),
    .A4(_2628_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3100_ (.I0(\mem[12][8] ),
    .I1(\mem[14][8] ),
    .S(_2174_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3101_ (.I0(_1739_),
    .I1(_2630_),
    .S(_2176_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3102_ (.I0(\mem[13][8] ),
    .I1(\mem[15][8] ),
    .S(_1822_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3103_ (.I0(_1740_),
    .I1(_2632_),
    .S(_2163_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3104_ (.A1(_1789_),
    .A2(_2631_),
    .B1(_2633_),
    .B2(_1780_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3105_ (.I0(\mem[8][8] ),
    .I1(\mem[10][8] ),
    .S(_1783_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3106_ (.A1(_1806_),
    .A2(_2635_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3107_ (.A1(_1378_),
    .A2(_1831_),
    .A3(_1745_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3108_ (.A1(_2636_),
    .A2(_2637_),
    .B(_1760_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3109_ (.A1(_1799_),
    .A2(_2629_),
    .A3(_2634_),
    .A4(_2638_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3110_ (.A1(_2618_),
    .A2(_2625_),
    .B(_2626_),
    .C(_2639_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3111_ (.A1(net114),
    .A2(_0611_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3112_ (.A1(_2162_),
    .A2(\mem[0][9] ),
    .A3(_1840_),
    .B1(_2164_),
    .B2(\mem[1][9] ),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _3113_ (.A1(_2166_),
    .A2(\mem[2][9] ),
    .A3(_2172_),
    .B1(_2167_),
    .B2(\mem[3][9] ),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3114_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2641_),
    .A4(_2642_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3115_ (.I0(\mem[4][9] ),
    .I1(\mem[6][9] ),
    .S(_1791_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3116_ (.I0(_1749_),
    .I1(_2644_),
    .S(_1793_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3117_ (.I0(\mem[5][9] ),
    .I1(\mem[7][9] ),
    .S(_2170_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3118_ (.I0(_1748_),
    .I1(_2646_),
    .S(_1771_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3119_ (.A1(_1790_),
    .A2(_2645_),
    .B1(_2647_),
    .B2(_2178_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3120_ (.I0(\mem[0][9] ),
    .I1(\mem[2][9] ),
    .S(_1816_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3121_ (.A1(_1806_),
    .A2(_2649_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3122_ (.A1(_2357_),
    .A2(_2151_),
    .A3(_1753_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3123_ (.A1(_2650_),
    .A2(_2651_),
    .B(_1760_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3124_ (.A1(_2144_),
    .A2(_2643_),
    .A3(_2648_),
    .A4(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3125_ (.I0(\mem[12][9] ),
    .I1(\mem[14][9] ),
    .S(_2361_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3126_ (.A1(_1735_),
    .A2(_1818_),
    .A3(_2654_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3127_ (.A1(_1808_),
    .A2(_1751_),
    .A3(_1786_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3128_ (.I0(\mem[9][9] ),
    .I1(\mem[11][9] ),
    .I2(\mem[13][9] ),
    .I3(\mem[15][9] ),
    .S0(_1800_),
    .S1(_1803_),
    .Z(_2657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3129_ (.I0(_1750_),
    .I1(_1756_),
    .S(_1376_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3130_ (.I0(\mem[8][9] ),
    .I1(\mem[10][9] ),
    .S(_1761_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3131_ (.A1(_1826_),
    .A2(_2659_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3132_ (.A1(_2152_),
    .A2(_1755_),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _3133_ (.I0(_2657_),
    .I1(_2658_),
    .I2(_2660_),
    .I3(_2661_),
    .S0(_1913_),
    .S1(_2370_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _3134_ (.A1(_1855_),
    .A2(_2655_),
    .A3(_2656_),
    .A4(_2662_),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3135_ (.A1(_2640_),
    .A2(_2653_),
    .A3(_2663_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3136_ (.I0(_0005_),
    .I1(_1811_),
    .S(_0000_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3137_ (.I0(_0006_),
    .I1(_1770_),
    .S(_0000_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3138_ (.A1(_2689_),
    .A2(_0000_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3139_ (.A1(_1379_),
    .A2(_2664_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3140_ (.A1(_2733_),
    .A2(_2727_),
    .B(_2726_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3141_ (.A1(_1733_),
    .A2(_0000_),
    .A3(_2665_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3142_ (.A1(_1364_),
    .A2(_2666_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3143_ (.I0(_0003_),
    .I1(\wr_ptr[0] ),
    .S(_0002_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3144_ (.I0(_0004_),
    .I1(\wr_ptr[1] ),
    .S(_0002_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3145_ (.A1(\wr_ptr[1] ),
    .A2(_2715_),
    .B(_2724_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3146_ (.A1(_0002_),
    .A2(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3147_ (.A1(_0620_),
    .A2(_2668_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3148_ (.I(_2717_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3149_ (.A1(_2669_),
    .A2(_2722_),
    .B(_2715_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3150_ (.A1(_2717_),
    .A2(_2722_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3151_ (.I0(_2670_),
    .I1(_2671_),
    .S(_2695_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3152_ (.A1(_0620_),
    .A2(_0002_),
    .A3(_2672_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3153_ (.A1(\wr_ptr[3] ),
    .A2(_2673_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3154_ (.A1(_2704_),
    .A2(_2742_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3155_ (.A1(_2740_),
    .A2(_2751_),
    .B1(_2674_),
    .B2(net73),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3156_ (.A1(_0615_),
    .A2(_2675_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3157_ (.A1(net72),
    .A2(net74),
    .A3(_0600_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3158_ (.A1(_2708_),
    .A2(_2704_),
    .A3(_2746_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3159_ (.A1(_2676_),
    .A2(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _3160_ (.A1(_2757_),
    .A2(_2751_),
    .B1(_2678_),
    .B2(_0607_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3161_ (.A1(_0607_),
    .A2(_2708_),
    .A3(_2674_),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3162_ (.A1(_2750_),
    .A2(_2693_),
    .Z(\next_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3163_ (.A1(_2690_),
    .A2(_2737_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3164_ (.A1(_2736_),
    .A2(_2679_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3165_ (.A1(_2750_),
    .A2(_2680_),
    .B(_2749_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3166_ (.A1(_2743_),
    .A2(_2681_),
    .Z(\next_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3167_ (.A1(_2750_),
    .A2(_2693_),
    .B(_2749_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3168_ (.I(_2744_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3169_ (.A1(_2743_),
    .A2(_2682_),
    .B(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3170_ (.A1(_2752_),
    .A2(_2684_),
    .ZN(\next_count[4] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3171_ (.A1(_2706_),
    .A2(_0594_),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3172_ (.A1(net74),
    .A2(_2759_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _3173_ (.A1(_2685_),
    .A2(_0615_),
    .B(_2707_),
    .C(net78),
    .ZN(net146));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3174_ (.I(_2706_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3175_ (.I(net72),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3176_ (.A1(net68),
    .A2(_2706_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3177_ (.I(_2755_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _3178_ (.A1(net73),
    .A2(net72),
    .A3(net74),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _3179_ (.A1(_2742_),
    .A2(_0592_),
    .A3(_0593_),
    .B(net76),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3180_ (.A1(_0591_),
    .A2(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3181_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3182_ (.I(_0596_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3183_ (.I(_2714_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3184_ (.I(\wr_ptr[1] ),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3185_ (.A1(net74),
    .A2(_2759_),
    .B(_2746_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3186_ (.A1(net73),
    .A2(net72),
    .A3(net68),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3187_ (.A1(net69),
    .A2(_2706_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _3188_ (.I(net76),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _3189_ (.A1(_0597_),
    .A2(_0598_),
    .B(_0599_),
    .C(_2704_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _3190_ (.I(_2751_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _3191_ (.A1(_0600_),
    .A2(_0593_),
    .B(net2),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _3192_ (.I(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3193_ (.I(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3194_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3195_ (.I(_0604_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3196_ (.I(_2709_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _3197_ (.A1(net73),
    .A2(net74),
    .A3(_0605_),
    .B(_2751_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3198_ (.I(net73),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3199_ (.A1(_0607_),
    .A2(_2704_),
    .A3(_2710_),
    .A4(_2742_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3200_ (.I(net3),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _3201_ (.A1(_2753_),
    .A2(_0606_),
    .B(_0608_),
    .C(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3202_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3203_ (.I(_0611_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3204_ (.I(\rd_ptr[1] ),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3205_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _3206_ (.I(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3207_ (.I(_0614_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3208_ (.I(_2733_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3209_ (.I(\wr_ptr[0] ),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3210_ (.I(_2731_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3211_ (.A1(net73),
    .A2(_2717_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3212_ (.I(_2738_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3213_ (.I(net74),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3214_ (.I(net75),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3215_ (.I(_2739_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3216_ (.A1(net73),
    .A2(net72),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3217_ (.A1(_2746_),
    .A2(_0615_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3218_ (.I(_2719_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3219_ (.A1(\wr_ptr[1] ),
    .A2(_2717_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3220_ (.I(_0601_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3221_ (.I(_2725_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3222_ (.A1(net73),
    .A2(_2715_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3223_ (.A1(_2735_),
    .A2(_0616_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3224_ (.I(net29),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3225_ (.I(net4),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3226_ (.I(\wr_ptr[3] ),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3227_ (.I(\wr_ptr[2] ),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3228_ (.A1(_0619_),
    .A2(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _3229_ (.A1(_2696_),
    .A2(_2714_),
    .A3(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3230_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3231_ (.I0(\mem[0][0] ),
    .I1(_0618_),
    .S(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3232_ (.A1(_2694_),
    .A2(_2695_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3233_ (.I(_2697_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3234_ (.A1(\wr_ptr[0] ),
    .A2(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _3235_ (.I0(_0625_),
    .I1(_0627_),
    .S(_0596_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3236_ (.A1(\wr_ptr[3] ),
    .A2(_2719_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3237_ (.A1(_0619_),
    .A2(_2719_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3238_ (.A1(\wr_ptr[0] ),
    .A2(\wr_ptr[1] ),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3239_ (.A1(\wr_ptr[2] ),
    .A2(_0591_),
    .A3(_0594_),
    .A4(_0631_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3240_ (.I0(_0629_),
    .I1(_0630_),
    .S(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3241_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3242_ (.A1(_2702_),
    .A2(_0591_),
    .A3(_0594_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3243_ (.A1(\wr_ptr[2] ),
    .A2(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3244_ (.I(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3245_ (.A1(_0628_),
    .A2(_0634_),
    .A3(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3246_ (.I(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3247_ (.I0(_0617_),
    .I1(_0624_),
    .S(_0639_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3248_ (.I(net40),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3249_ (.I(net5),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3250_ (.I0(\mem[0][10] ),
    .I1(_0641_),
    .S(_0623_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3251_ (.I0(_0640_),
    .I1(_0642_),
    .S(_0639_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3252_ (.I(net41),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3253_ (.I(net6),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3254_ (.I0(\mem[0][11] ),
    .I1(_0644_),
    .S(_0623_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3255_ (.I0(_0643_),
    .I1(_0645_),
    .S(_0639_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3256_ (.I(net42),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3257_ (.I(net7),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3258_ (.I0(\mem[0][12] ),
    .I1(_0647_),
    .S(_0623_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3259_ (.I0(_0646_),
    .I1(_0648_),
    .S(_0639_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3260_ (.I(net43),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3261_ (.I(net8),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3262_ (.I0(\mem[0][13] ),
    .I1(_0650_),
    .S(_0623_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3263_ (.I0(_0649_),
    .I1(_0651_),
    .S(_0639_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3264_ (.I(net44),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3265_ (.I(net9),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3266_ (.I0(\mem[0][14] ),
    .I1(_0653_),
    .S(_0623_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3267_ (.I0(_0652_),
    .I1(_0654_),
    .S(_0639_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3268_ (.I(net45),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3269_ (.I(net10),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3270_ (.I0(\mem[0][15] ),
    .I1(_0656_),
    .S(_0623_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3271_ (.I0(_0655_),
    .I1(_0657_),
    .S(_0639_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3272_ (.I(net46),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3273_ (.I(net11),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3274_ (.I0(\mem[0][16] ),
    .I1(_0659_),
    .S(_0623_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3275_ (.I0(_0658_),
    .I1(_0660_),
    .S(_0639_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3276_ (.I(net47),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3277_ (.I(net12),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3278_ (.I0(\mem[0][17] ),
    .I1(_0662_),
    .S(_0623_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3279_ (.I0(_0661_),
    .I1(_0663_),
    .S(_0639_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3280_ (.I(net49),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3281_ (.I(net13),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3282_ (.I0(\mem[0][18] ),
    .I1(_0665_),
    .S(_0623_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3283_ (.I0(_0664_),
    .I1(_0666_),
    .S(_0639_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3284_ (.I(net50),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3285_ (.I(net14),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3286_ (.I(_0622_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3287_ (.I0(\mem[0][19] ),
    .I1(_0668_),
    .S(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3288_ (.I(_0638_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3289_ (.I0(_0667_),
    .I1(_0670_),
    .S(_0671_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3290_ (.I(net30),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3291_ (.I(net15),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3292_ (.I0(\mem[0][1] ),
    .I1(_0673_),
    .S(_0669_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3293_ (.I0(_0672_),
    .I1(_0674_),
    .S(_0671_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3294_ (.I(net51),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3295_ (.I(net16),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3296_ (.I0(\mem[0][20] ),
    .I1(_0676_),
    .S(_0669_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3297_ (.I0(_0675_),
    .I1(_0677_),
    .S(_0671_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3298_ (.I(net52),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3299_ (.I(net17),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3300_ (.I0(\mem[0][21] ),
    .I1(_0679_),
    .S(_0669_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3301_ (.I0(_0678_),
    .I1(_0680_),
    .S(_0671_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3302_ (.I(net53),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3303_ (.I(net18),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3304_ (.I0(\mem[0][22] ),
    .I1(_0682_),
    .S(_0669_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3305_ (.I0(_0681_),
    .I1(_0683_),
    .S(_0671_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3306_ (.I(net54),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3307_ (.I(net19),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3308_ (.I0(\mem[0][23] ),
    .I1(_0685_),
    .S(_0669_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3309_ (.I0(_0684_),
    .I1(_0686_),
    .S(_0671_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3310_ (.I(net55),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3311_ (.I(net20),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3312_ (.I0(\mem[0][24] ),
    .I1(_0688_),
    .S(_0669_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3313_ (.I0(_0687_),
    .I1(_0689_),
    .S(_0671_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3314_ (.I(net56),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3315_ (.I(net21),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3316_ (.I0(\mem[0][25] ),
    .I1(_0691_),
    .S(_0669_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3317_ (.I0(_0690_),
    .I1(_0692_),
    .S(_0671_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3318_ (.I(net57),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3319_ (.I(net22),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3320_ (.I0(\mem[0][26] ),
    .I1(_0694_),
    .S(_0669_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3321_ (.I0(_0693_),
    .I1(_0695_),
    .S(_0671_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3322_ (.I(net58),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3323_ (.I(net23),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3324_ (.I0(\mem[0][27] ),
    .I1(_0697_),
    .S(_0669_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3325_ (.I0(_0696_),
    .I1(_0698_),
    .S(_0671_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3326_ (.I(net60),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3327_ (.I(net24),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3328_ (.I(_0622_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3329_ (.I0(\mem[0][28] ),
    .I1(_0700_),
    .S(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3330_ (.I(_0638_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3331_ (.I0(_0699_),
    .I1(_0702_),
    .S(_0703_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3332_ (.I(net61),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3333_ (.I(net25),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3334_ (.I0(\mem[0][29] ),
    .I1(_0705_),
    .S(_0701_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3335_ (.I0(_0704_),
    .I1(_0706_),
    .S(_0703_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3336_ (.I(net31),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3337_ (.I(net26),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3338_ (.I0(\mem[0][2] ),
    .I1(_0708_),
    .S(_0701_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3339_ (.I0(_0707_),
    .I1(_0709_),
    .S(_0703_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3340_ (.I(net62),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3341_ (.I(net27),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3342_ (.I0(\mem[0][30] ),
    .I1(_0711_),
    .S(_0701_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3343_ (.I0(_0710_),
    .I1(_0712_),
    .S(_0703_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3344_ (.I(net63),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3345_ (.I(net28),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3346_ (.I0(\mem[0][31] ),
    .I1(_0714_),
    .S(_0701_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3347_ (.I0(_0713_),
    .I1(_0715_),
    .S(_0703_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3348_ (.I(net32),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3349_ (.I(net37),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3350_ (.I0(\mem[0][3] ),
    .I1(_0717_),
    .S(_0701_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3351_ (.I0(_0716_),
    .I1(_0718_),
    .S(_0703_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3352_ (.I(net33),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3353_ (.I(net48),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3354_ (.I0(\mem[0][4] ),
    .I1(_0720_),
    .S(_0701_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3355_ (.I0(_0719_),
    .I1(_0721_),
    .S(_0703_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3356_ (.I(net34),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3357_ (.I(net59),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3358_ (.I0(\mem[0][5] ),
    .I1(_0723_),
    .S(_0701_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3359_ (.I0(_0722_),
    .I1(_0724_),
    .S(_0703_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3360_ (.I(net35),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _3361_ (.I(net64),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3362_ (.I0(\mem[0][6] ),
    .I1(_0726_),
    .S(_0701_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3363_ (.I0(_0725_),
    .I1(_0727_),
    .S(_0703_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3364_ (.I(net36),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3365_ (.I(net65),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3366_ (.I0(\mem[0][7] ),
    .I1(_0729_),
    .S(_0701_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3367_ (.I0(_0728_),
    .I1(_0730_),
    .S(_0703_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3368_ (.I(net38),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3369_ (.I(net66),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3370_ (.I0(\mem[0][8] ),
    .I1(_0732_),
    .S(_0622_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3371_ (.I0(_0731_),
    .I1(_0733_),
    .S(_0638_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3372_ (.I(net39),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _3373_ (.I(net67),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3374_ (.I0(\mem[0][9] ),
    .I1(_0735_),
    .S(_0622_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3375_ (.I0(_0734_),
    .I1(_0736_),
    .S(_0638_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3376_ (.A1(\wr_ptr[3] ),
    .A2(_0620_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _3377_ (.A1(_2698_),
    .A2(_2714_),
    .A3(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3378_ (.I(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3379_ (.I0(\mem[10][0] ),
    .I1(_0618_),
    .S(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3380_ (.A1(_2694_),
    .A2(\wr_ptr[1] ),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3381_ (.A1(\wr_ptr[0] ),
    .A2(_2697_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _3382_ (.I0(_0741_),
    .I1(_0742_),
    .S(_0596_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3383_ (.I0(_0630_),
    .I1(_0629_),
    .S(_0632_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3384_ (.I(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3385_ (.A1(_0637_),
    .A2(_0743_),
    .A3(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3386_ (.I(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3387_ (.I0(_0617_),
    .I1(_0740_),
    .S(_0747_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3388_ (.I0(\mem[10][10] ),
    .I1(_0641_),
    .S(_0739_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3389_ (.I0(_0640_),
    .I1(_0748_),
    .S(_0747_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3390_ (.I0(\mem[10][11] ),
    .I1(_0644_),
    .S(_0739_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3391_ (.I0(_0643_),
    .I1(_0749_),
    .S(_0747_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3392_ (.I0(\mem[10][12] ),
    .I1(_0647_),
    .S(_0739_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3393_ (.I0(_0646_),
    .I1(_0750_),
    .S(_0747_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3394_ (.I0(\mem[10][13] ),
    .I1(_0650_),
    .S(_0739_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3395_ (.I0(_0649_),
    .I1(_0751_),
    .S(_0747_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3396_ (.I0(\mem[10][14] ),
    .I1(_0653_),
    .S(_0739_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3397_ (.I0(_0652_),
    .I1(_0752_),
    .S(_0747_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3398_ (.I0(\mem[10][15] ),
    .I1(_0656_),
    .S(_0739_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3399_ (.I0(_0655_),
    .I1(_0753_),
    .S(_0747_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3400_ (.I0(\mem[10][16] ),
    .I1(_0659_),
    .S(_0739_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3401_ (.I0(_0658_),
    .I1(_0754_),
    .S(_0747_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3402_ (.I0(\mem[10][17] ),
    .I1(_0662_),
    .S(_0739_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3403_ (.I0(_0661_),
    .I1(_0755_),
    .S(_0747_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3404_ (.I0(\mem[10][18] ),
    .I1(_0665_),
    .S(_0739_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3405_ (.I0(_0664_),
    .I1(_0756_),
    .S(_0747_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3406_ (.I(_0738_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3407_ (.I0(\mem[10][19] ),
    .I1(_0668_),
    .S(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3408_ (.I(_0746_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3409_ (.I0(_0667_),
    .I1(_0758_),
    .S(_0759_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3410_ (.I0(\mem[10][1] ),
    .I1(_0673_),
    .S(_0757_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3411_ (.I0(_0672_),
    .I1(_0760_),
    .S(_0759_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3412_ (.I0(\mem[10][20] ),
    .I1(_0676_),
    .S(_0757_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3413_ (.I0(_0675_),
    .I1(_0761_),
    .S(_0759_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3414_ (.I0(\mem[10][21] ),
    .I1(_0679_),
    .S(_0757_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3415_ (.I0(_0678_),
    .I1(_0762_),
    .S(_0759_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3416_ (.I0(\mem[10][22] ),
    .I1(_0682_),
    .S(_0757_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3417_ (.I0(_0681_),
    .I1(_0763_),
    .S(_0759_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3418_ (.I0(\mem[10][23] ),
    .I1(_0685_),
    .S(_0757_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3419_ (.I0(_0684_),
    .I1(_0764_),
    .S(_0759_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3420_ (.I0(\mem[10][24] ),
    .I1(_0688_),
    .S(_0757_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3421_ (.I0(_0687_),
    .I1(_0765_),
    .S(_0759_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3422_ (.I0(\mem[10][25] ),
    .I1(_0691_),
    .S(_0757_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3423_ (.I0(_0690_),
    .I1(_0766_),
    .S(_0759_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3424_ (.I0(\mem[10][26] ),
    .I1(_0694_),
    .S(_0757_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3425_ (.I0(_0693_),
    .I1(_0767_),
    .S(_0759_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3426_ (.I0(\mem[10][27] ),
    .I1(_0697_),
    .S(_0757_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3427_ (.I0(_0696_),
    .I1(_0768_),
    .S(_0759_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3428_ (.I(_0738_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3429_ (.I0(\mem[10][28] ),
    .I1(_0700_),
    .S(_0769_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3430_ (.I(_0746_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3431_ (.I0(_0699_),
    .I1(_0770_),
    .S(_0771_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3432_ (.I0(\mem[10][29] ),
    .I1(_0705_),
    .S(_0769_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3433_ (.I0(_0704_),
    .I1(_0772_),
    .S(_0771_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3434_ (.I0(\mem[10][2] ),
    .I1(_0708_),
    .S(_0769_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3435_ (.I0(_0707_),
    .I1(_0773_),
    .S(_0771_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3436_ (.I0(\mem[10][30] ),
    .I1(_0711_),
    .S(_0769_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3437_ (.I0(_0710_),
    .I1(_0774_),
    .S(_0771_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3438_ (.I0(\mem[10][31] ),
    .I1(_0714_),
    .S(_0769_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3439_ (.I0(_0713_),
    .I1(_0775_),
    .S(_0771_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3440_ (.I0(\mem[10][3] ),
    .I1(_0717_),
    .S(_0769_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3441_ (.I0(_0716_),
    .I1(_0776_),
    .S(_0771_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3442_ (.I0(\mem[10][4] ),
    .I1(_0720_),
    .S(_0769_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3443_ (.I0(_0719_),
    .I1(_0777_),
    .S(_0771_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3444_ (.I0(\mem[10][5] ),
    .I1(_0723_),
    .S(_0769_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3445_ (.I0(_0722_),
    .I1(_0778_),
    .S(_0771_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3446_ (.I0(\mem[10][6] ),
    .I1(_0726_),
    .S(_0769_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3447_ (.I0(_0725_),
    .I1(_0779_),
    .S(_0771_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3448_ (.I0(\mem[10][7] ),
    .I1(_0729_),
    .S(_0769_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3449_ (.I0(_0728_),
    .I1(_0780_),
    .S(_0771_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3450_ (.I0(\mem[10][8] ),
    .I1(_0732_),
    .S(_0738_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3451_ (.I0(_0731_),
    .I1(_0781_),
    .S(_0746_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3452_ (.I0(\mem[10][9] ),
    .I1(_0735_),
    .S(_0738_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3453_ (.I0(_0734_),
    .I1(_0782_),
    .S(_0746_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _3454_ (.A1(_0635_),
    .A2(_0737_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3455_ (.I(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3456_ (.I0(\mem[11][0] ),
    .I1(_0618_),
    .S(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3457_ (.A1(_2694_),
    .A2(_2697_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _3458_ (.I0(_0631_),
    .I1(_0786_),
    .S(_0596_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3459_ (.A1(_0637_),
    .A2(_0745_),
    .A3(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3460_ (.I(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3461_ (.I0(_0617_),
    .I1(_0785_),
    .S(_0789_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3462_ (.I0(\mem[11][10] ),
    .I1(_0641_),
    .S(_0784_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3463_ (.I0(_0640_),
    .I1(_0790_),
    .S(_0789_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3464_ (.I0(\mem[11][11] ),
    .I1(_0644_),
    .S(_0784_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3465_ (.I0(_0643_),
    .I1(_0791_),
    .S(_0789_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3466_ (.I0(\mem[11][12] ),
    .I1(_0647_),
    .S(_0784_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3467_ (.I0(_0646_),
    .I1(_0792_),
    .S(_0789_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3468_ (.I0(\mem[11][13] ),
    .I1(_0650_),
    .S(_0784_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3469_ (.I0(_0649_),
    .I1(_0793_),
    .S(_0789_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3470_ (.I0(\mem[11][14] ),
    .I1(_0653_),
    .S(_0784_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3471_ (.I0(_0652_),
    .I1(_0794_),
    .S(_0789_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3472_ (.I0(\mem[11][15] ),
    .I1(_0656_),
    .S(_0784_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3473_ (.I0(_0655_),
    .I1(_0795_),
    .S(_0789_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3474_ (.I0(\mem[11][16] ),
    .I1(_0659_),
    .S(_0784_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3475_ (.I0(_0658_),
    .I1(_0796_),
    .S(_0789_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3476_ (.I0(\mem[11][17] ),
    .I1(_0662_),
    .S(_0784_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3477_ (.I0(_0661_),
    .I1(_0797_),
    .S(_0789_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3478_ (.I0(\mem[11][18] ),
    .I1(_0665_),
    .S(_0784_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3479_ (.I0(_0664_),
    .I1(_0798_),
    .S(_0789_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3480_ (.I(_0783_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3481_ (.I0(\mem[11][19] ),
    .I1(_0668_),
    .S(_0799_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3482_ (.I(_0788_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3483_ (.I0(_0667_),
    .I1(_0800_),
    .S(_0801_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3484_ (.I0(\mem[11][1] ),
    .I1(_0673_),
    .S(_0799_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3485_ (.I0(_0672_),
    .I1(_0802_),
    .S(_0801_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3486_ (.I0(\mem[11][20] ),
    .I1(_0676_),
    .S(_0799_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3487_ (.I0(_0675_),
    .I1(_0803_),
    .S(_0801_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3488_ (.I0(\mem[11][21] ),
    .I1(_0679_),
    .S(_0799_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3489_ (.I0(_0678_),
    .I1(_0804_),
    .S(_0801_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3490_ (.I0(\mem[11][22] ),
    .I1(_0682_),
    .S(_0799_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3491_ (.I0(_0681_),
    .I1(_0805_),
    .S(_0801_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3492_ (.I0(\mem[11][23] ),
    .I1(_0685_),
    .S(_0799_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3493_ (.I0(_0684_),
    .I1(_0806_),
    .S(_0801_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3494_ (.I0(\mem[11][24] ),
    .I1(_0688_),
    .S(_0799_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3495_ (.I0(_0687_),
    .I1(_0807_),
    .S(_0801_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3496_ (.I0(\mem[11][25] ),
    .I1(_0691_),
    .S(_0799_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3497_ (.I0(_0690_),
    .I1(_0808_),
    .S(_0801_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3498_ (.I0(\mem[11][26] ),
    .I1(_0694_),
    .S(_0799_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3499_ (.I0(_0693_),
    .I1(_0809_),
    .S(_0801_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3500_ (.I0(\mem[11][27] ),
    .I1(_0697_),
    .S(_0799_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3501_ (.I0(_0696_),
    .I1(_0810_),
    .S(_0801_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3502_ (.I(_0783_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3503_ (.I0(\mem[11][28] ),
    .I1(_0700_),
    .S(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3504_ (.I(_0788_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3505_ (.I0(_0699_),
    .I1(_0812_),
    .S(_0813_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3506_ (.I0(\mem[11][29] ),
    .I1(_0705_),
    .S(_0811_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3507_ (.I0(_0704_),
    .I1(_0814_),
    .S(_0813_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3508_ (.I0(\mem[11][2] ),
    .I1(_0708_),
    .S(_0811_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3509_ (.I0(_0707_),
    .I1(_0815_),
    .S(_0813_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3510_ (.I0(\mem[11][30] ),
    .I1(_0711_),
    .S(_0811_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3511_ (.I0(_0710_),
    .I1(_0816_),
    .S(_0813_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3512_ (.I0(\mem[11][31] ),
    .I1(_0714_),
    .S(_0811_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3513_ (.I0(_0713_),
    .I1(_0817_),
    .S(_0813_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3514_ (.I0(\mem[11][3] ),
    .I1(_0717_),
    .S(_0811_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3515_ (.I0(_0716_),
    .I1(_0818_),
    .S(_0813_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3516_ (.I0(\mem[11][4] ),
    .I1(_0720_),
    .S(_0811_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3517_ (.I0(_0719_),
    .I1(_0819_),
    .S(_0813_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3518_ (.I0(\mem[11][5] ),
    .I1(_0723_),
    .S(_0811_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3519_ (.I0(_0722_),
    .I1(_0820_),
    .S(_0813_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3520_ (.I0(\mem[11][6] ),
    .I1(_0726_),
    .S(_0811_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3521_ (.I0(_0725_),
    .I1(_0821_),
    .S(_0813_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3522_ (.I0(\mem[11][7] ),
    .I1(_0729_),
    .S(_0811_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3523_ (.I0(_0728_),
    .I1(_0822_),
    .S(_0813_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3524_ (.I0(\mem[11][8] ),
    .I1(_0732_),
    .S(_0783_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3525_ (.I0(_0731_),
    .I1(_0823_),
    .S(_0788_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3526_ (.I0(\mem[11][9] ),
    .I1(_0735_),
    .S(_0783_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3527_ (.I0(_0734_),
    .I1(_0824_),
    .S(_0788_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _3528_ (.A1(\wr_ptr[3] ),
    .A2(\wr_ptr[2] ),
    .A3(_2696_),
    .A4(_0596_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3529_ (.I(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3530_ (.I0(\mem[12][0] ),
    .I1(_0618_),
    .S(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3531_ (.A1(_0620_),
    .A2(_0635_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3532_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3533_ (.A1(_0628_),
    .A2(_0829_),
    .A3(_0745_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3534_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3535_ (.I0(_0617_),
    .I1(_0827_),
    .S(_0831_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3536_ (.I0(\mem[12][10] ),
    .I1(_0641_),
    .S(_0826_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3537_ (.I0(_0640_),
    .I1(_0832_),
    .S(_0831_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3538_ (.I0(\mem[12][11] ),
    .I1(_0644_),
    .S(_0826_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3539_ (.I0(_0643_),
    .I1(_0833_),
    .S(_0831_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3540_ (.I0(\mem[12][12] ),
    .I1(_0647_),
    .S(_0826_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3541_ (.I0(_0646_),
    .I1(_0834_),
    .S(_0831_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3542_ (.I0(\mem[12][13] ),
    .I1(_0650_),
    .S(_0826_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3543_ (.I0(_0649_),
    .I1(_0835_),
    .S(_0831_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3544_ (.I0(\mem[12][14] ),
    .I1(_0653_),
    .S(_0826_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3545_ (.I0(_0652_),
    .I1(_0836_),
    .S(_0831_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3546_ (.I0(\mem[12][15] ),
    .I1(_0656_),
    .S(_0826_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3547_ (.I0(_0655_),
    .I1(_0837_),
    .S(_0831_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3548_ (.I0(\mem[12][16] ),
    .I1(_0659_),
    .S(_0826_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3549_ (.I0(_0658_),
    .I1(_0838_),
    .S(_0831_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3550_ (.I0(\mem[12][17] ),
    .I1(_0662_),
    .S(_0826_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3551_ (.I0(_0661_),
    .I1(_0839_),
    .S(_0831_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3552_ (.I0(\mem[12][18] ),
    .I1(_0665_),
    .S(_0826_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3553_ (.I0(_0664_),
    .I1(_0840_),
    .S(_0831_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3554_ (.I(_0825_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3555_ (.I0(\mem[12][19] ),
    .I1(_0668_),
    .S(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3556_ (.I(_0830_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3557_ (.I0(_0667_),
    .I1(_0842_),
    .S(_0843_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3558_ (.I0(\mem[12][1] ),
    .I1(_0673_),
    .S(_0841_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3559_ (.I0(_0672_),
    .I1(_0844_),
    .S(_0843_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3560_ (.I0(\mem[12][20] ),
    .I1(_0676_),
    .S(_0841_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3561_ (.I0(_0675_),
    .I1(_0845_),
    .S(_0843_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3562_ (.I0(\mem[12][21] ),
    .I1(_0679_),
    .S(_0841_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3563_ (.I0(_0678_),
    .I1(_0846_),
    .S(_0843_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3564_ (.I0(\mem[12][22] ),
    .I1(_0682_),
    .S(_0841_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3565_ (.I0(_0681_),
    .I1(_0847_),
    .S(_0843_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3566_ (.I0(\mem[12][23] ),
    .I1(_0685_),
    .S(_0841_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3567_ (.I0(_0684_),
    .I1(_0848_),
    .S(_0843_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3568_ (.I0(\mem[12][24] ),
    .I1(_0688_),
    .S(_0841_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3569_ (.I0(_0687_),
    .I1(_0849_),
    .S(_0843_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3570_ (.I0(\mem[12][25] ),
    .I1(_0691_),
    .S(_0841_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3571_ (.I0(_0690_),
    .I1(_0850_),
    .S(_0843_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3572_ (.I0(\mem[12][26] ),
    .I1(_0694_),
    .S(_0841_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3573_ (.I0(_0693_),
    .I1(_0851_),
    .S(_0843_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3574_ (.I0(\mem[12][27] ),
    .I1(_0697_),
    .S(_0841_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3575_ (.I0(_0696_),
    .I1(_0852_),
    .S(_0843_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3576_ (.I(_0825_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3577_ (.I0(\mem[12][28] ),
    .I1(_0700_),
    .S(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3578_ (.I(_0830_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3579_ (.I0(_0699_),
    .I1(_0854_),
    .S(_0855_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3580_ (.I0(\mem[12][29] ),
    .I1(_0705_),
    .S(_0853_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3581_ (.I0(_0704_),
    .I1(_0856_),
    .S(_0855_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3582_ (.I0(\mem[12][2] ),
    .I1(_0708_),
    .S(_0853_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3583_ (.I0(_0707_),
    .I1(_0857_),
    .S(_0855_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3584_ (.I0(\mem[12][30] ),
    .I1(_0711_),
    .S(_0853_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3585_ (.I0(_0710_),
    .I1(_0858_),
    .S(_0855_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3586_ (.I0(\mem[12][31] ),
    .I1(_0714_),
    .S(_0853_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3587_ (.I0(_0713_),
    .I1(_0859_),
    .S(_0855_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3588_ (.I0(\mem[12][3] ),
    .I1(_0717_),
    .S(_0853_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3589_ (.I0(_0716_),
    .I1(_0860_),
    .S(_0855_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3590_ (.I0(\mem[12][4] ),
    .I1(_0720_),
    .S(_0853_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3591_ (.I0(_0719_),
    .I1(_0861_),
    .S(_0855_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3592_ (.I0(\mem[12][5] ),
    .I1(_0723_),
    .S(_0853_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3593_ (.I0(_0722_),
    .I1(_0862_),
    .S(_0855_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3594_ (.I0(\mem[12][6] ),
    .I1(_0726_),
    .S(_0853_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3595_ (.I0(_0725_),
    .I1(_0863_),
    .S(_0855_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3596_ (.I0(\mem[12][7] ),
    .I1(_0729_),
    .S(_0853_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3597_ (.I0(_0728_),
    .I1(_0864_),
    .S(_0855_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3598_ (.I0(\mem[12][8] ),
    .I1(_0732_),
    .S(_0825_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3599_ (.I0(_0731_),
    .I1(_0865_),
    .S(_0830_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3600_ (.I0(\mem[12][9] ),
    .I1(_0735_),
    .S(_0825_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3601_ (.I0(_0734_),
    .I1(_0866_),
    .S(_0830_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _3602_ (.A1(\wr_ptr[3] ),
    .A2(\wr_ptr[2] ),
    .A3(_2700_),
    .A4(_0596_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3603_ (.I(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3604_ (.I0(\mem[13][0] ),
    .I1(_0618_),
    .S(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3605_ (.A1(\wr_ptr[0] ),
    .A2(_2695_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3606_ (.A1(_2694_),
    .A2(_0626_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _3607_ (.I0(_0870_),
    .I1(_0871_),
    .S(_0596_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3608_ (.A1(_0829_),
    .A2(_0745_),
    .A3(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3609_ (.I(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3610_ (.I0(_0617_),
    .I1(_0869_),
    .S(_0874_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3611_ (.I0(\mem[13][10] ),
    .I1(_0641_),
    .S(_0868_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3612_ (.I0(_0640_),
    .I1(_0875_),
    .S(_0874_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3613_ (.I0(\mem[13][11] ),
    .I1(_0644_),
    .S(_0868_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3614_ (.I0(_0643_),
    .I1(_0876_),
    .S(_0874_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3615_ (.I0(\mem[13][12] ),
    .I1(_0647_),
    .S(_0868_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3616_ (.I0(_0646_),
    .I1(_0877_),
    .S(_0874_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3617_ (.I0(\mem[13][13] ),
    .I1(_0650_),
    .S(_0868_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3618_ (.I0(_0649_),
    .I1(_0878_),
    .S(_0874_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3619_ (.I0(\mem[13][14] ),
    .I1(_0653_),
    .S(_0868_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3620_ (.I0(_0652_),
    .I1(_0879_),
    .S(_0874_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3621_ (.I0(\mem[13][15] ),
    .I1(_0656_),
    .S(_0868_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3622_ (.I0(_0655_),
    .I1(_0880_),
    .S(_0874_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3623_ (.I0(\mem[13][16] ),
    .I1(_0659_),
    .S(_0868_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3624_ (.I0(_0658_),
    .I1(_0881_),
    .S(_0874_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3625_ (.I0(\mem[13][17] ),
    .I1(_0662_),
    .S(_0868_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3626_ (.I0(_0661_),
    .I1(_0882_),
    .S(_0874_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3627_ (.I0(\mem[13][18] ),
    .I1(_0665_),
    .S(_0868_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3628_ (.I0(_0664_),
    .I1(_0883_),
    .S(_0874_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3629_ (.I(_0867_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3630_ (.I0(\mem[13][19] ),
    .I1(_0668_),
    .S(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3631_ (.I(_0873_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3632_ (.I0(_0667_),
    .I1(_0885_),
    .S(_0886_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3633_ (.I0(\mem[13][1] ),
    .I1(_0673_),
    .S(_0884_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3634_ (.I0(_0672_),
    .I1(_0887_),
    .S(_0886_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3635_ (.I0(\mem[13][20] ),
    .I1(_0676_),
    .S(_0884_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3636_ (.I0(_0675_),
    .I1(_0888_),
    .S(_0886_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3637_ (.I0(\mem[13][21] ),
    .I1(_0679_),
    .S(_0884_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3638_ (.I0(_0678_),
    .I1(_0889_),
    .S(_0886_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3639_ (.I0(\mem[13][22] ),
    .I1(_0682_),
    .S(_0884_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3640_ (.I0(_0681_),
    .I1(_0890_),
    .S(_0886_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3641_ (.I0(\mem[13][23] ),
    .I1(_0685_),
    .S(_0884_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3642_ (.I0(_0684_),
    .I1(_0891_),
    .S(_0886_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3643_ (.I0(\mem[13][24] ),
    .I1(_0688_),
    .S(_0884_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3644_ (.I0(_0687_),
    .I1(_0892_),
    .S(_0886_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3645_ (.I0(\mem[13][25] ),
    .I1(_0691_),
    .S(_0884_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3646_ (.I0(_0690_),
    .I1(_0893_),
    .S(_0886_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3647_ (.I0(\mem[13][26] ),
    .I1(_0694_),
    .S(_0884_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3648_ (.I0(_0693_),
    .I1(_0894_),
    .S(_0886_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3649_ (.I0(\mem[13][27] ),
    .I1(_0697_),
    .S(_0884_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3650_ (.I0(_0696_),
    .I1(_0895_),
    .S(_0886_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3651_ (.I(_0867_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3652_ (.I0(\mem[13][28] ),
    .I1(_0700_),
    .S(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3653_ (.I(_0873_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3654_ (.I0(_0699_),
    .I1(_0897_),
    .S(_0898_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3655_ (.I0(\mem[13][29] ),
    .I1(_0705_),
    .S(_0896_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3656_ (.I0(_0704_),
    .I1(_0899_),
    .S(_0898_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3657_ (.I0(\mem[13][2] ),
    .I1(_0708_),
    .S(_0896_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3658_ (.I0(_0707_),
    .I1(_0900_),
    .S(_0898_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3659_ (.I0(\mem[13][30] ),
    .I1(_0711_),
    .S(_0896_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3660_ (.I0(_0710_),
    .I1(_0901_),
    .S(_0898_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3661_ (.I0(\mem[13][31] ),
    .I1(_0714_),
    .S(_0896_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3662_ (.I0(_0713_),
    .I1(_0902_),
    .S(_0898_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3663_ (.I0(\mem[13][3] ),
    .I1(_0717_),
    .S(_0896_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3664_ (.I0(_0716_),
    .I1(_0903_),
    .S(_0898_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3665_ (.I0(\mem[13][4] ),
    .I1(_0720_),
    .S(_0896_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3666_ (.I0(_0719_),
    .I1(_0904_),
    .S(_0898_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3667_ (.I0(\mem[13][5] ),
    .I1(_0723_),
    .S(_0896_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3668_ (.I0(_0722_),
    .I1(_0905_),
    .S(_0898_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3669_ (.I0(\mem[13][6] ),
    .I1(_0726_),
    .S(_0896_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3670_ (.I0(_0725_),
    .I1(_0906_),
    .S(_0898_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3671_ (.I0(\mem[13][7] ),
    .I1(_0729_),
    .S(_0896_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3672_ (.I0(_0728_),
    .I1(_0907_),
    .S(_0898_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3673_ (.I0(\mem[13][8] ),
    .I1(_0732_),
    .S(_0867_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3674_ (.I0(_0731_),
    .I1(_0908_),
    .S(_0873_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3675_ (.I0(\mem[13][9] ),
    .I1(_0735_),
    .S(_0867_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3676_ (.I0(_0734_),
    .I1(_0909_),
    .S(_0873_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _3677_ (.A1(\wr_ptr[3] ),
    .A2(\wr_ptr[2] ),
    .A3(_2698_),
    .A4(_0596_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3678_ (.I(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3679_ (.I0(\mem[14][0] ),
    .I1(_0618_),
    .S(_0911_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3680_ (.A1(_0829_),
    .A2(_0743_),
    .A3(_0745_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3681_ (.I(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3682_ (.I0(_0617_),
    .I1(_0912_),
    .S(_0914_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3683_ (.I0(\mem[14][10] ),
    .I1(_0641_),
    .S(_0911_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3684_ (.I0(_0640_),
    .I1(_0915_),
    .S(_0914_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3685_ (.I0(\mem[14][11] ),
    .I1(_0644_),
    .S(_0911_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3686_ (.I0(_0643_),
    .I1(_0916_),
    .S(_0914_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3687_ (.I0(\mem[14][12] ),
    .I1(_0647_),
    .S(_0911_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3688_ (.I0(_0646_),
    .I1(_0917_),
    .S(_0914_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3689_ (.I0(\mem[14][13] ),
    .I1(_0650_),
    .S(_0911_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3690_ (.I0(_0649_),
    .I1(_0918_),
    .S(_0914_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3691_ (.I0(\mem[14][14] ),
    .I1(_0653_),
    .S(_0911_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3692_ (.I0(_0652_),
    .I1(_0919_),
    .S(_0914_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3693_ (.I0(\mem[14][15] ),
    .I1(_0656_),
    .S(_0911_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3694_ (.I0(_0655_),
    .I1(_0920_),
    .S(_0914_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3695_ (.I0(\mem[14][16] ),
    .I1(_0659_),
    .S(_0911_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3696_ (.I0(_0658_),
    .I1(_0921_),
    .S(_0914_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3697_ (.I0(\mem[14][17] ),
    .I1(_0662_),
    .S(_0911_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3698_ (.I0(_0661_),
    .I1(_0922_),
    .S(_0914_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3699_ (.I0(\mem[14][18] ),
    .I1(_0665_),
    .S(_0911_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3700_ (.I0(_0664_),
    .I1(_0923_),
    .S(_0914_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3701_ (.I(_0910_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3702_ (.I0(\mem[14][19] ),
    .I1(_0668_),
    .S(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3703_ (.I(_0913_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3704_ (.I0(_0667_),
    .I1(_0925_),
    .S(_0926_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3705_ (.I0(\mem[14][1] ),
    .I1(_0673_),
    .S(_0924_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3706_ (.I0(_0672_),
    .I1(_0927_),
    .S(_0926_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3707_ (.I0(\mem[14][20] ),
    .I1(_0676_),
    .S(_0924_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3708_ (.I0(_0675_),
    .I1(_0928_),
    .S(_0926_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3709_ (.I0(\mem[14][21] ),
    .I1(_0679_),
    .S(_0924_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3710_ (.I0(_0678_),
    .I1(_0929_),
    .S(_0926_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3711_ (.I0(\mem[14][22] ),
    .I1(_0682_),
    .S(_0924_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3712_ (.I0(_0681_),
    .I1(_0930_),
    .S(_0926_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3713_ (.I0(\mem[14][23] ),
    .I1(_0685_),
    .S(_0924_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3714_ (.I0(_0684_),
    .I1(_0931_),
    .S(_0926_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3715_ (.I0(\mem[14][24] ),
    .I1(_0688_),
    .S(_0924_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3716_ (.I0(_0687_),
    .I1(_0932_),
    .S(_0926_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3717_ (.I0(\mem[14][25] ),
    .I1(_0691_),
    .S(_0924_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3718_ (.I0(_0690_),
    .I1(_0933_),
    .S(_0926_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3719_ (.I0(\mem[14][26] ),
    .I1(_0694_),
    .S(_0924_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3720_ (.I0(_0693_),
    .I1(_0934_),
    .S(_0926_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3721_ (.I0(\mem[14][27] ),
    .I1(_0697_),
    .S(_0924_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3722_ (.I0(_0696_),
    .I1(_0935_),
    .S(_0926_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3723_ (.I(_0910_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3724_ (.I0(\mem[14][28] ),
    .I1(_0700_),
    .S(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3725_ (.I(_0913_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3726_ (.I0(_0699_),
    .I1(_0937_),
    .S(_0938_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3727_ (.I0(\mem[14][29] ),
    .I1(_0705_),
    .S(_0936_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3728_ (.I0(_0704_),
    .I1(_0939_),
    .S(_0938_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3729_ (.I0(\mem[14][2] ),
    .I1(_0708_),
    .S(_0936_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3730_ (.I0(_0707_),
    .I1(_0940_),
    .S(_0938_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3731_ (.I0(\mem[14][30] ),
    .I1(_0711_),
    .S(_0936_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3732_ (.I0(_0710_),
    .I1(_0941_),
    .S(_0938_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3733_ (.I0(\mem[14][31] ),
    .I1(_0714_),
    .S(_0936_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3734_ (.I0(_0713_),
    .I1(_0942_),
    .S(_0938_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3735_ (.I0(\mem[14][3] ),
    .I1(_0717_),
    .S(_0936_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3736_ (.I0(_0716_),
    .I1(_0943_),
    .S(_0938_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3737_ (.I0(\mem[14][4] ),
    .I1(_0720_),
    .S(_0936_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3738_ (.I0(_0719_),
    .I1(_0944_),
    .S(_0938_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3739_ (.I0(\mem[14][5] ),
    .I1(_0723_),
    .S(_0936_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3740_ (.I0(_0722_),
    .I1(_0945_),
    .S(_0938_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3741_ (.I0(\mem[14][6] ),
    .I1(_0726_),
    .S(_0936_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3742_ (.I0(_0725_),
    .I1(_0946_),
    .S(_0938_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3743_ (.I0(\mem[14][7] ),
    .I1(_0729_),
    .S(_0936_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3744_ (.I0(_0728_),
    .I1(_0947_),
    .S(_0938_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3745_ (.I0(\mem[14][8] ),
    .I1(_0732_),
    .S(_0910_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3746_ (.I0(_0731_),
    .I1(_0948_),
    .S(_0913_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3747_ (.I0(\mem[14][9] ),
    .I1(_0735_),
    .S(_0910_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3748_ (.I0(_0734_),
    .I1(_0949_),
    .S(_0913_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _3749_ (.A1(\wr_ptr[3] ),
    .A2(\wr_ptr[2] ),
    .A3(_0635_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3750_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3751_ (.I0(\mem[15][0] ),
    .I1(_0618_),
    .S(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3752_ (.A1(_0829_),
    .A2(_0745_),
    .A3(_0787_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3753_ (.I(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3754_ (.I0(_0617_),
    .I1(_0952_),
    .S(_0954_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3755_ (.I0(\mem[15][10] ),
    .I1(_0641_),
    .S(_0951_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3756_ (.I0(_0640_),
    .I1(_0955_),
    .S(_0954_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3757_ (.I0(\mem[15][11] ),
    .I1(_0644_),
    .S(_0951_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3758_ (.I0(_0643_),
    .I1(_0956_),
    .S(_0954_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3759_ (.I0(\mem[15][12] ),
    .I1(_0647_),
    .S(_0951_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3760_ (.I0(_0646_),
    .I1(_0957_),
    .S(_0954_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3761_ (.I0(\mem[15][13] ),
    .I1(_0650_),
    .S(_0951_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3762_ (.I0(_0649_),
    .I1(_0958_),
    .S(_0954_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3763_ (.I0(\mem[15][14] ),
    .I1(_0653_),
    .S(_0951_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3764_ (.I0(_0652_),
    .I1(_0959_),
    .S(_0954_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3765_ (.I0(\mem[15][15] ),
    .I1(_0656_),
    .S(_0951_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3766_ (.I0(_0655_),
    .I1(_0960_),
    .S(_0954_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3767_ (.I0(\mem[15][16] ),
    .I1(_0659_),
    .S(_0951_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3768_ (.I0(_0658_),
    .I1(_0961_),
    .S(_0954_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3769_ (.I0(\mem[15][17] ),
    .I1(_0662_),
    .S(_0951_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3770_ (.I0(_0661_),
    .I1(_0962_),
    .S(_0954_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3771_ (.I0(\mem[15][18] ),
    .I1(_0665_),
    .S(_0951_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3772_ (.I0(_0664_),
    .I1(_0963_),
    .S(_0954_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3773_ (.I(_0950_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3774_ (.I0(\mem[15][19] ),
    .I1(_0668_),
    .S(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3775_ (.I(_0953_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3776_ (.I0(_0667_),
    .I1(_0965_),
    .S(_0966_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3777_ (.I0(\mem[15][1] ),
    .I1(_0673_),
    .S(_0964_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3778_ (.I0(_0672_),
    .I1(_0967_),
    .S(_0966_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3779_ (.I0(\mem[15][20] ),
    .I1(_0676_),
    .S(_0964_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3780_ (.I0(_0675_),
    .I1(_0968_),
    .S(_0966_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3781_ (.I0(\mem[15][21] ),
    .I1(_0679_),
    .S(_0964_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3782_ (.I0(_0678_),
    .I1(_0969_),
    .S(_0966_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3783_ (.I0(\mem[15][22] ),
    .I1(_0682_),
    .S(_0964_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3784_ (.I0(_0681_),
    .I1(_0970_),
    .S(_0966_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3785_ (.I0(\mem[15][23] ),
    .I1(_0685_),
    .S(_0964_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3786_ (.I0(_0684_),
    .I1(_0971_),
    .S(_0966_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3787_ (.I0(\mem[15][24] ),
    .I1(_0688_),
    .S(_0964_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3788_ (.I0(_0687_),
    .I1(_0972_),
    .S(_0966_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3789_ (.I0(\mem[15][25] ),
    .I1(_0691_),
    .S(_0964_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3790_ (.I0(_0690_),
    .I1(_0973_),
    .S(_0966_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3791_ (.I0(\mem[15][26] ),
    .I1(_0694_),
    .S(_0964_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3792_ (.I0(_0693_),
    .I1(_0974_),
    .S(_0966_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3793_ (.I0(\mem[15][27] ),
    .I1(_0697_),
    .S(_0964_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3794_ (.I0(_0696_),
    .I1(_0975_),
    .S(_0966_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3795_ (.I(_0950_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3796_ (.I0(\mem[15][28] ),
    .I1(_0700_),
    .S(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3797_ (.I(_0953_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3798_ (.I0(_0699_),
    .I1(_0977_),
    .S(_0978_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3799_ (.I0(\mem[15][29] ),
    .I1(_0705_),
    .S(_0976_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3800_ (.I0(_0704_),
    .I1(_0979_),
    .S(_0978_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3801_ (.I0(\mem[15][2] ),
    .I1(_0708_),
    .S(_0976_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3802_ (.I0(_0707_),
    .I1(_0980_),
    .S(_0978_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3803_ (.I0(\mem[15][30] ),
    .I1(_0711_),
    .S(_0976_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3804_ (.I0(_0710_),
    .I1(_0981_),
    .S(_0978_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3805_ (.I0(\mem[15][31] ),
    .I1(_0714_),
    .S(_0976_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3806_ (.I0(_0713_),
    .I1(_0982_),
    .S(_0978_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3807_ (.I0(\mem[15][3] ),
    .I1(_0717_),
    .S(_0976_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3808_ (.I0(_0716_),
    .I1(_0983_),
    .S(_0978_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3809_ (.I0(\mem[15][4] ),
    .I1(_0720_),
    .S(_0976_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3810_ (.I0(_0719_),
    .I1(_0984_),
    .S(_0978_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3811_ (.I0(\mem[15][5] ),
    .I1(_0723_),
    .S(_0976_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3812_ (.I0(_0722_),
    .I1(_0985_),
    .S(_0978_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3813_ (.I0(\mem[15][6] ),
    .I1(_0726_),
    .S(_0976_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3814_ (.I0(_0725_),
    .I1(_0986_),
    .S(_0978_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3815_ (.I0(\mem[15][7] ),
    .I1(_0729_),
    .S(_0976_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3816_ (.I0(_0728_),
    .I1(_0987_),
    .S(_0978_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3817_ (.I0(\mem[15][8] ),
    .I1(_0732_),
    .S(_0950_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3818_ (.I0(_0731_),
    .I1(_0988_),
    .S(_0953_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3819_ (.I0(\mem[15][9] ),
    .I1(_0735_),
    .S(_0950_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3820_ (.I0(_0734_),
    .I1(_0989_),
    .S(_0953_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _3821_ (.A1(_2700_),
    .A2(_2714_),
    .A3(_0621_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3822_ (.I(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3823_ (.I0(\mem[1][0] ),
    .I1(_0618_),
    .S(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3824_ (.A1(_0634_),
    .A2(_0637_),
    .A3(_0872_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3825_ (.I(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3826_ (.I0(_0617_),
    .I1(_0992_),
    .S(_0994_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3827_ (.I0(\mem[1][10] ),
    .I1(_0641_),
    .S(_0991_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3828_ (.I0(_0640_),
    .I1(_0995_),
    .S(_0994_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3829_ (.I0(\mem[1][11] ),
    .I1(_0644_),
    .S(_0991_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3830_ (.I0(_0643_),
    .I1(_0996_),
    .S(_0994_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3831_ (.I0(\mem[1][12] ),
    .I1(_0647_),
    .S(_0991_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3832_ (.I0(_0646_),
    .I1(_0997_),
    .S(_0994_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3833_ (.I0(\mem[1][13] ),
    .I1(_0650_),
    .S(_0991_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3834_ (.I0(_0649_),
    .I1(_0998_),
    .S(_0994_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3835_ (.I0(\mem[1][14] ),
    .I1(_0653_),
    .S(_0991_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3836_ (.I0(_0652_),
    .I1(_0999_),
    .S(_0994_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3837_ (.I0(\mem[1][15] ),
    .I1(_0656_),
    .S(_0991_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3838_ (.I0(_0655_),
    .I1(_1000_),
    .S(_0994_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3839_ (.I0(\mem[1][16] ),
    .I1(_0659_),
    .S(_0991_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3840_ (.I0(_0658_),
    .I1(_1001_),
    .S(_0994_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3841_ (.I0(\mem[1][17] ),
    .I1(_0662_),
    .S(_0991_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3842_ (.I0(_0661_),
    .I1(_1002_),
    .S(_0994_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3843_ (.I0(\mem[1][18] ),
    .I1(_0665_),
    .S(_0991_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3844_ (.I0(_0664_),
    .I1(_1003_),
    .S(_0994_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3845_ (.I(_0990_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3846_ (.I0(\mem[1][19] ),
    .I1(_0668_),
    .S(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3847_ (.I(_0993_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3848_ (.I0(_0667_),
    .I1(_1005_),
    .S(_1006_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3849_ (.I0(\mem[1][1] ),
    .I1(_0673_),
    .S(_1004_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3850_ (.I0(_0672_),
    .I1(_1007_),
    .S(_1006_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3851_ (.I0(\mem[1][20] ),
    .I1(_0676_),
    .S(_1004_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3852_ (.I0(_0675_),
    .I1(_1008_),
    .S(_1006_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3853_ (.I0(\mem[1][21] ),
    .I1(_0679_),
    .S(_1004_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3854_ (.I0(_0678_),
    .I1(_1009_),
    .S(_1006_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3855_ (.I0(\mem[1][22] ),
    .I1(_0682_),
    .S(_1004_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3856_ (.I0(_0681_),
    .I1(_1010_),
    .S(_1006_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3857_ (.I0(\mem[1][23] ),
    .I1(_0685_),
    .S(_1004_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3858_ (.I0(_0684_),
    .I1(_1011_),
    .S(_1006_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3859_ (.I0(\mem[1][24] ),
    .I1(_0688_),
    .S(_1004_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3860_ (.I0(_0687_),
    .I1(_1012_),
    .S(_1006_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3861_ (.I0(\mem[1][25] ),
    .I1(_0691_),
    .S(_1004_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3862_ (.I0(_0690_),
    .I1(_1013_),
    .S(_1006_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3863_ (.I0(\mem[1][26] ),
    .I1(_0694_),
    .S(_1004_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3864_ (.I0(_0693_),
    .I1(_1014_),
    .S(_1006_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3865_ (.I0(\mem[1][27] ),
    .I1(_0697_),
    .S(_1004_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3866_ (.I0(_0696_),
    .I1(_1015_),
    .S(_1006_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3867_ (.I(_0990_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3868_ (.I0(\mem[1][28] ),
    .I1(_0700_),
    .S(_1016_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3869_ (.I(_0993_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3870_ (.I0(_0699_),
    .I1(_1017_),
    .S(_1018_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3871_ (.I0(\mem[1][29] ),
    .I1(_0705_),
    .S(_1016_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3872_ (.I0(_0704_),
    .I1(_1019_),
    .S(_1018_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3873_ (.I0(\mem[1][2] ),
    .I1(_0708_),
    .S(_1016_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3874_ (.I0(_0707_),
    .I1(_1020_),
    .S(_1018_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3875_ (.I0(\mem[1][30] ),
    .I1(_0711_),
    .S(_1016_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3876_ (.I0(_0710_),
    .I1(_1021_),
    .S(_1018_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3877_ (.I0(\mem[1][31] ),
    .I1(_0714_),
    .S(_1016_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3878_ (.I0(_0713_),
    .I1(_1022_),
    .S(_1018_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3879_ (.I0(\mem[1][3] ),
    .I1(_0717_),
    .S(_1016_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3880_ (.I0(_0716_),
    .I1(_1023_),
    .S(_1018_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3881_ (.I0(\mem[1][4] ),
    .I1(_0720_),
    .S(_1016_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3882_ (.I0(_0719_),
    .I1(_1024_),
    .S(_1018_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3883_ (.I0(\mem[1][5] ),
    .I1(_0723_),
    .S(_1016_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3884_ (.I0(_0722_),
    .I1(_1025_),
    .S(_1018_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3885_ (.I0(\mem[1][6] ),
    .I1(_0726_),
    .S(_1016_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3886_ (.I0(_0725_),
    .I1(_1026_),
    .S(_1018_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3887_ (.I0(\mem[1][7] ),
    .I1(_0729_),
    .S(_1016_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3888_ (.I0(_0728_),
    .I1(_1027_),
    .S(_1018_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3889_ (.I0(\mem[1][8] ),
    .I1(_0732_),
    .S(_0990_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3890_ (.I0(_0731_),
    .I1(_1028_),
    .S(_0993_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3891_ (.I0(\mem[1][9] ),
    .I1(_0735_),
    .S(_0990_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3892_ (.I0(_0734_),
    .I1(_1029_),
    .S(_0993_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _3893_ (.A1(_2698_),
    .A2(_2714_),
    .A3(_0621_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3894_ (.I(_1030_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3895_ (.I0(\mem[2][0] ),
    .I1(_0618_),
    .S(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3896_ (.A1(_0634_),
    .A2(_0637_),
    .A3(_0743_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3897_ (.I(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3898_ (.I0(_0617_),
    .I1(_1032_),
    .S(_1034_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3899_ (.I0(\mem[2][10] ),
    .I1(_0641_),
    .S(_1031_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3900_ (.I0(_0640_),
    .I1(_1035_),
    .S(_1034_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3901_ (.I0(\mem[2][11] ),
    .I1(_0644_),
    .S(_1031_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3902_ (.I0(_0643_),
    .I1(_1036_),
    .S(_1034_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3903_ (.I0(\mem[2][12] ),
    .I1(_0647_),
    .S(_1031_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3904_ (.I0(_0646_),
    .I1(_1037_),
    .S(_1034_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3905_ (.I0(\mem[2][13] ),
    .I1(_0650_),
    .S(_1031_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3906_ (.I0(_0649_),
    .I1(_1038_),
    .S(_1034_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3907_ (.I0(\mem[2][14] ),
    .I1(_0653_),
    .S(_1031_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3908_ (.I0(_0652_),
    .I1(_1039_),
    .S(_1034_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3909_ (.I0(\mem[2][15] ),
    .I1(_0656_),
    .S(_1031_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3910_ (.I0(_0655_),
    .I1(_1040_),
    .S(_1034_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3911_ (.I0(\mem[2][16] ),
    .I1(_0659_),
    .S(_1031_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3912_ (.I0(_0658_),
    .I1(_1041_),
    .S(_1034_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3913_ (.I0(\mem[2][17] ),
    .I1(_0662_),
    .S(_1031_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3914_ (.I0(_0661_),
    .I1(_1042_),
    .S(_1034_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3915_ (.I0(\mem[2][18] ),
    .I1(_0665_),
    .S(_1031_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3916_ (.I0(_0664_),
    .I1(_1043_),
    .S(_1034_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _3917_ (.I(_1030_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3918_ (.I0(\mem[2][19] ),
    .I1(_0668_),
    .S(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3919_ (.I(_1033_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3920_ (.I0(_0667_),
    .I1(_1045_),
    .S(_1046_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3921_ (.I0(\mem[2][1] ),
    .I1(_0673_),
    .S(_1044_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3922_ (.I0(_0672_),
    .I1(_1047_),
    .S(_1046_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3923_ (.I0(\mem[2][20] ),
    .I1(_0676_),
    .S(_1044_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3924_ (.I0(_0675_),
    .I1(_1048_),
    .S(_1046_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3925_ (.I0(\mem[2][21] ),
    .I1(_0679_),
    .S(_1044_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3926_ (.I0(_0678_),
    .I1(_1049_),
    .S(_1046_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3927_ (.I0(\mem[2][22] ),
    .I1(_0682_),
    .S(_1044_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3928_ (.I0(_0681_),
    .I1(_1050_),
    .S(_1046_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3929_ (.I0(\mem[2][23] ),
    .I1(_0685_),
    .S(_1044_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3930_ (.I0(_0684_),
    .I1(_1051_),
    .S(_1046_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3931_ (.I0(\mem[2][24] ),
    .I1(_0688_),
    .S(_1044_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3932_ (.I0(_0687_),
    .I1(_1052_),
    .S(_1046_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3933_ (.I0(\mem[2][25] ),
    .I1(_0691_),
    .S(_1044_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3934_ (.I0(_0690_),
    .I1(_1053_),
    .S(_1046_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3935_ (.I0(\mem[2][26] ),
    .I1(_0694_),
    .S(_1044_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3936_ (.I0(_0693_),
    .I1(_1054_),
    .S(_1046_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3937_ (.I0(\mem[2][27] ),
    .I1(_0697_),
    .S(_1044_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3938_ (.I0(_0696_),
    .I1(_1055_),
    .S(_1046_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3939_ (.I(_1030_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3940_ (.I0(\mem[2][28] ),
    .I1(_0700_),
    .S(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _3941_ (.I(_1033_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3942_ (.I0(_0699_),
    .I1(_1057_),
    .S(_1058_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3943_ (.I0(\mem[2][29] ),
    .I1(_0705_),
    .S(_1056_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3944_ (.I0(_0704_),
    .I1(_1059_),
    .S(_1058_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3945_ (.I0(\mem[2][2] ),
    .I1(_0708_),
    .S(_1056_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3946_ (.I0(_0707_),
    .I1(_1060_),
    .S(_1058_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3947_ (.I0(\mem[2][30] ),
    .I1(_0711_),
    .S(_1056_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3948_ (.I0(_0710_),
    .I1(_1061_),
    .S(_1058_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3949_ (.I0(\mem[2][31] ),
    .I1(_0714_),
    .S(_1056_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3950_ (.I0(_0713_),
    .I1(_1062_),
    .S(_1058_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3951_ (.I0(\mem[2][3] ),
    .I1(_0717_),
    .S(_1056_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3952_ (.I0(_0716_),
    .I1(_1063_),
    .S(_1058_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3953_ (.I0(\mem[2][4] ),
    .I1(_0720_),
    .S(_1056_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3954_ (.I0(_0719_),
    .I1(_1064_),
    .S(_1058_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3955_ (.I0(\mem[2][5] ),
    .I1(_0723_),
    .S(_1056_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3956_ (.I0(_0722_),
    .I1(_1065_),
    .S(_1058_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3957_ (.I0(\mem[2][6] ),
    .I1(_0726_),
    .S(_1056_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3958_ (.I0(_0725_),
    .I1(_1066_),
    .S(_1058_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3959_ (.I0(\mem[2][7] ),
    .I1(_0729_),
    .S(_1056_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3960_ (.I0(_0728_),
    .I1(_1067_),
    .S(_1058_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3961_ (.I0(\mem[2][8] ),
    .I1(_0732_),
    .S(_1030_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3962_ (.I0(_0731_),
    .I1(_1068_),
    .S(_1033_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3963_ (.I0(\mem[2][9] ),
    .I1(_0735_),
    .S(_1030_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3964_ (.I0(_0734_),
    .I1(_1069_),
    .S(_1033_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _3965_ (.A1(_0635_),
    .A2(_0621_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3966_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3967_ (.I0(\mem[3][0] ),
    .I1(_0618_),
    .S(_1071_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3968_ (.A1(_0634_),
    .A2(_0637_),
    .A3(_0787_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3969_ (.I(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3970_ (.I0(_0617_),
    .I1(_1072_),
    .S(_1074_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3971_ (.I0(\mem[3][10] ),
    .I1(_0641_),
    .S(_1071_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3972_ (.I0(_0640_),
    .I1(_1075_),
    .S(_1074_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3973_ (.I0(\mem[3][11] ),
    .I1(_0644_),
    .S(_1071_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3974_ (.I0(_0643_),
    .I1(_1076_),
    .S(_1074_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3975_ (.I0(\mem[3][12] ),
    .I1(_0647_),
    .S(_1071_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3976_ (.I0(_0646_),
    .I1(_1077_),
    .S(_1074_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3977_ (.I0(\mem[3][13] ),
    .I1(_0650_),
    .S(_1071_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3978_ (.I0(_0649_),
    .I1(_1078_),
    .S(_1074_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3979_ (.I0(\mem[3][14] ),
    .I1(_0653_),
    .S(_1071_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3980_ (.I0(_0652_),
    .I1(_1079_),
    .S(_1074_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3981_ (.I0(\mem[3][15] ),
    .I1(_0656_),
    .S(_1071_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3982_ (.I0(_0655_),
    .I1(_1080_),
    .S(_1074_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3983_ (.I0(\mem[3][16] ),
    .I1(_0659_),
    .S(_1071_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3984_ (.I0(_0658_),
    .I1(_1081_),
    .S(_1074_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3985_ (.I0(\mem[3][17] ),
    .I1(_0662_),
    .S(_1071_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3986_ (.I0(_0661_),
    .I1(_1082_),
    .S(_1074_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3987_ (.I0(\mem[3][18] ),
    .I1(_0665_),
    .S(_1071_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3988_ (.I0(_0664_),
    .I1(_1083_),
    .S(_1074_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3989_ (.I(_1070_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3990_ (.I0(\mem[3][19] ),
    .I1(_0668_),
    .S(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _3991_ (.I(_1073_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3992_ (.I0(_0667_),
    .I1(_1085_),
    .S(_1086_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3993_ (.I0(\mem[3][1] ),
    .I1(_0673_),
    .S(_1084_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3994_ (.I0(_0672_),
    .I1(_1087_),
    .S(_1086_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3995_ (.I0(\mem[3][20] ),
    .I1(_0676_),
    .S(_1084_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3996_ (.I0(_0675_),
    .I1(_1088_),
    .S(_1086_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3997_ (.I0(\mem[3][21] ),
    .I1(_0679_),
    .S(_1084_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3998_ (.I0(_0678_),
    .I1(_1089_),
    .S(_1086_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3999_ (.I0(\mem[3][22] ),
    .I1(_0682_),
    .S(_1084_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4000_ (.I0(_0681_),
    .I1(_1090_),
    .S(_1086_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4001_ (.I0(\mem[3][23] ),
    .I1(_0685_),
    .S(_1084_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4002_ (.I0(_0684_),
    .I1(_1091_),
    .S(_1086_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4003_ (.I0(\mem[3][24] ),
    .I1(_0688_),
    .S(_1084_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4004_ (.I0(_0687_),
    .I1(_1092_),
    .S(_1086_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4005_ (.I0(\mem[3][25] ),
    .I1(_0691_),
    .S(_1084_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4006_ (.I0(_0690_),
    .I1(_1093_),
    .S(_1086_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4007_ (.I0(\mem[3][26] ),
    .I1(_0694_),
    .S(_1084_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4008_ (.I0(_0693_),
    .I1(_1094_),
    .S(_1086_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4009_ (.I0(\mem[3][27] ),
    .I1(_0697_),
    .S(_1084_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4010_ (.I0(_0696_),
    .I1(_1095_),
    .S(_1086_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4011_ (.I(_1070_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4012_ (.I0(\mem[3][28] ),
    .I1(_0700_),
    .S(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4013_ (.I(_1073_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4014_ (.I0(_0699_),
    .I1(_1097_),
    .S(_1098_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4015_ (.I0(\mem[3][29] ),
    .I1(_0705_),
    .S(_1096_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4016_ (.I0(_0704_),
    .I1(_1099_),
    .S(_1098_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4017_ (.I0(\mem[3][2] ),
    .I1(_0708_),
    .S(_1096_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4018_ (.I0(_0707_),
    .I1(_1100_),
    .S(_1098_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4019_ (.I0(\mem[3][30] ),
    .I1(_0711_),
    .S(_1096_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4020_ (.I0(_0710_),
    .I1(_1101_),
    .S(_1098_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4021_ (.I0(\mem[3][31] ),
    .I1(_0714_),
    .S(_1096_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4022_ (.I0(_0713_),
    .I1(_1102_),
    .S(_1098_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4023_ (.I0(\mem[3][3] ),
    .I1(_0717_),
    .S(_1096_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4024_ (.I0(_0716_),
    .I1(_1103_),
    .S(_1098_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4025_ (.I0(\mem[3][4] ),
    .I1(_0720_),
    .S(_1096_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4026_ (.I0(_0719_),
    .I1(_1104_),
    .S(_1098_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4027_ (.I0(\mem[3][5] ),
    .I1(_0723_),
    .S(_1096_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4028_ (.I0(_0722_),
    .I1(_1105_),
    .S(_1098_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4029_ (.I0(\mem[3][6] ),
    .I1(_0726_),
    .S(_1096_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4030_ (.I0(_0725_),
    .I1(_1106_),
    .S(_1098_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4031_ (.I0(\mem[3][7] ),
    .I1(_0729_),
    .S(_1096_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4032_ (.I0(_0728_),
    .I1(_1107_),
    .S(_1098_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4033_ (.I0(\mem[3][8] ),
    .I1(_0732_),
    .S(_1070_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4034_ (.I0(_0731_),
    .I1(_1108_),
    .S(_1073_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4035_ (.I0(\mem[3][9] ),
    .I1(_0735_),
    .S(_1070_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4036_ (.I0(_0734_),
    .I1(_1109_),
    .S(_1073_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4037_ (.A1(_0619_),
    .A2(\wr_ptr[2] ),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _4038_ (.A1(_2696_),
    .A2(_2714_),
    .A3(_1110_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4039_ (.I(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4040_ (.I0(\mem[4][0] ),
    .I1(net4),
    .S(_1112_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4041_ (.A1(_0628_),
    .A2(_0634_),
    .A3(_0829_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4042_ (.I(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4043_ (.I0(net29),
    .I1(_1113_),
    .S(_1115_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4044_ (.I0(\mem[4][10] ),
    .I1(net5),
    .S(_1112_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4045_ (.I0(net40),
    .I1(_1116_),
    .S(_1115_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4046_ (.I0(\mem[4][11] ),
    .I1(net6),
    .S(_1112_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4047_ (.I0(net41),
    .I1(_1117_),
    .S(_1115_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4048_ (.I0(\mem[4][12] ),
    .I1(net7),
    .S(_1112_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4049_ (.I0(net42),
    .I1(_1118_),
    .S(_1115_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4050_ (.I0(\mem[4][13] ),
    .I1(net8),
    .S(_1112_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4051_ (.I0(net43),
    .I1(_1119_),
    .S(_1115_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4052_ (.I0(\mem[4][14] ),
    .I1(net9),
    .S(_1112_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4053_ (.I0(net44),
    .I1(_1120_),
    .S(_1115_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4054_ (.I0(\mem[4][15] ),
    .I1(net10),
    .S(_1112_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4055_ (.I0(net45),
    .I1(_1121_),
    .S(_1115_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4056_ (.I0(\mem[4][16] ),
    .I1(net11),
    .S(_1112_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4057_ (.I0(net46),
    .I1(_1122_),
    .S(_1115_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4058_ (.I0(\mem[4][17] ),
    .I1(net12),
    .S(_1112_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4059_ (.I0(net47),
    .I1(_1123_),
    .S(_1115_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4060_ (.I0(\mem[4][18] ),
    .I1(net13),
    .S(_1112_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4061_ (.I0(net49),
    .I1(_1124_),
    .S(_1115_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4062_ (.I(_1111_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4063_ (.I0(\mem[4][19] ),
    .I1(net14),
    .S(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4064_ (.I(_1114_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4065_ (.I0(net50),
    .I1(_1126_),
    .S(_1127_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4066_ (.I0(\mem[4][1] ),
    .I1(net15),
    .S(_1125_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4067_ (.I0(net30),
    .I1(_1128_),
    .S(_1127_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4068_ (.I0(\mem[4][20] ),
    .I1(net16),
    .S(_1125_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4069_ (.I0(net51),
    .I1(_1129_),
    .S(_1127_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4070_ (.I0(\mem[4][21] ),
    .I1(net17),
    .S(_1125_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4071_ (.I0(net52),
    .I1(_1130_),
    .S(_1127_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4072_ (.I0(\mem[4][22] ),
    .I1(net18),
    .S(_1125_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4073_ (.I0(net53),
    .I1(_1131_),
    .S(_1127_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4074_ (.I0(\mem[4][23] ),
    .I1(net19),
    .S(_1125_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4075_ (.I0(net54),
    .I1(_1132_),
    .S(_1127_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4076_ (.I0(\mem[4][24] ),
    .I1(net20),
    .S(_1125_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4077_ (.I0(net55),
    .I1(_1133_),
    .S(_1127_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4078_ (.I0(\mem[4][25] ),
    .I1(net21),
    .S(_1125_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4079_ (.I0(net56),
    .I1(_1134_),
    .S(_1127_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4080_ (.I0(\mem[4][26] ),
    .I1(net22),
    .S(_1125_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4081_ (.I0(net57),
    .I1(_1135_),
    .S(_1127_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4082_ (.I0(\mem[4][27] ),
    .I1(net23),
    .S(_1125_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4083_ (.I0(net58),
    .I1(_1136_),
    .S(_1127_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4084_ (.I(_1111_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4085_ (.I0(\mem[4][28] ),
    .I1(net24),
    .S(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4086_ (.I(_1114_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4087_ (.I0(net60),
    .I1(_1138_),
    .S(_1139_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4088_ (.I0(\mem[4][29] ),
    .I1(net25),
    .S(_1137_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4089_ (.I0(net61),
    .I1(_1140_),
    .S(_1139_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4090_ (.I0(\mem[4][2] ),
    .I1(net26),
    .S(_1137_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4091_ (.I0(net31),
    .I1(_1141_),
    .S(_1139_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4092_ (.I0(\mem[4][30] ),
    .I1(net27),
    .S(_1137_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4093_ (.I0(net62),
    .I1(_1142_),
    .S(_1139_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4094_ (.I0(\mem[4][31] ),
    .I1(net28),
    .S(_1137_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4095_ (.I0(net63),
    .I1(_1143_),
    .S(_1139_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4096_ (.I0(\mem[4][3] ),
    .I1(net37),
    .S(_1137_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4097_ (.I0(net32),
    .I1(_1144_),
    .S(_1139_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4098_ (.I0(\mem[4][4] ),
    .I1(net48),
    .S(_1137_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4099_ (.I0(net33),
    .I1(_1145_),
    .S(_1139_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4100_ (.I0(\mem[4][5] ),
    .I1(net59),
    .S(_1137_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4101_ (.I0(net34),
    .I1(_1146_),
    .S(_1139_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4102_ (.I0(\mem[4][6] ),
    .I1(net64),
    .S(_1137_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4103_ (.I0(net35),
    .I1(_1147_),
    .S(_1139_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4104_ (.I0(\mem[4][7] ),
    .I1(net65),
    .S(_1137_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4105_ (.I0(net36),
    .I1(_1148_),
    .S(_1139_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4106_ (.I0(\mem[4][8] ),
    .I1(net66),
    .S(_1111_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4107_ (.I0(net38),
    .I1(_1149_),
    .S(_1114_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4108_ (.I0(\mem[4][9] ),
    .I1(net67),
    .S(_1111_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4109_ (.I0(net39),
    .I1(_1150_),
    .S(_1114_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _4110_ (.A1(_2700_),
    .A2(_2714_),
    .A3(_1110_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4111_ (.I(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4112_ (.I0(\mem[5][0] ),
    .I1(net4),
    .S(_1152_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4113_ (.A1(_0634_),
    .A2(_0829_),
    .A3(_0872_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4114_ (.I(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4115_ (.I0(net29),
    .I1(_1153_),
    .S(_1155_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4116_ (.I0(\mem[5][10] ),
    .I1(net5),
    .S(_1152_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4117_ (.I0(net40),
    .I1(_1156_),
    .S(_1155_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4118_ (.I0(\mem[5][11] ),
    .I1(net6),
    .S(_1152_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4119_ (.I0(net41),
    .I1(_1157_),
    .S(_1155_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4120_ (.I0(\mem[5][12] ),
    .I1(net7),
    .S(_1152_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4121_ (.I0(net42),
    .I1(_1158_),
    .S(_1155_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4122_ (.I0(\mem[5][13] ),
    .I1(net8),
    .S(_1152_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4123_ (.I0(net43),
    .I1(_1159_),
    .S(_1155_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4124_ (.I0(\mem[5][14] ),
    .I1(net9),
    .S(_1152_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4125_ (.I0(net44),
    .I1(_1160_),
    .S(_1155_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4126_ (.I0(\mem[5][15] ),
    .I1(net10),
    .S(_1152_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4127_ (.I0(net45),
    .I1(_1161_),
    .S(_1155_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4128_ (.I0(\mem[5][16] ),
    .I1(net11),
    .S(_1152_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4129_ (.I0(net46),
    .I1(_1162_),
    .S(_1155_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4130_ (.I0(\mem[5][17] ),
    .I1(net12),
    .S(_1152_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4131_ (.I0(net47),
    .I1(_1163_),
    .S(_1155_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4132_ (.I0(\mem[5][18] ),
    .I1(net13),
    .S(_1152_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4133_ (.I0(net49),
    .I1(_1164_),
    .S(_1155_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4134_ (.I(_1151_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4135_ (.I0(\mem[5][19] ),
    .I1(net14),
    .S(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4136_ (.I(_1154_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4137_ (.I0(net50),
    .I1(_1166_),
    .S(_1167_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4138_ (.I0(\mem[5][1] ),
    .I1(net15),
    .S(_1165_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4139_ (.I0(net30),
    .I1(_1168_),
    .S(_1167_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4140_ (.I0(\mem[5][20] ),
    .I1(net16),
    .S(_1165_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4141_ (.I0(net51),
    .I1(_1169_),
    .S(_1167_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4142_ (.I0(\mem[5][21] ),
    .I1(net17),
    .S(_1165_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4143_ (.I0(net52),
    .I1(_1170_),
    .S(_1167_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4144_ (.I0(\mem[5][22] ),
    .I1(net18),
    .S(_1165_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4145_ (.I0(net53),
    .I1(_1171_),
    .S(_1167_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4146_ (.I0(\mem[5][23] ),
    .I1(net19),
    .S(_1165_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4147_ (.I0(net54),
    .I1(_1172_),
    .S(_1167_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4148_ (.I0(\mem[5][24] ),
    .I1(net20),
    .S(_1165_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4149_ (.I0(net55),
    .I1(_1173_),
    .S(_1167_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4150_ (.I0(\mem[5][25] ),
    .I1(net21),
    .S(_1165_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4151_ (.I0(net56),
    .I1(_1174_),
    .S(_1167_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4152_ (.I0(\mem[5][26] ),
    .I1(net22),
    .S(_1165_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4153_ (.I0(net57),
    .I1(_1175_),
    .S(_1167_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4154_ (.I0(\mem[5][27] ),
    .I1(net23),
    .S(_1165_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4155_ (.I0(net58),
    .I1(_1176_),
    .S(_1167_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4156_ (.I(_1151_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4157_ (.I0(\mem[5][28] ),
    .I1(net24),
    .S(_1177_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4158_ (.I(_1154_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4159_ (.I0(net60),
    .I1(_1178_),
    .S(_1179_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4160_ (.I0(\mem[5][29] ),
    .I1(net25),
    .S(_1177_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4161_ (.I0(net61),
    .I1(_1180_),
    .S(_1179_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4162_ (.I0(\mem[5][2] ),
    .I1(net26),
    .S(_1177_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4163_ (.I0(net31),
    .I1(_1181_),
    .S(_1179_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4164_ (.I0(\mem[5][30] ),
    .I1(net27),
    .S(_1177_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4165_ (.I0(net62),
    .I1(_1182_),
    .S(_1179_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4166_ (.I0(\mem[5][31] ),
    .I1(net28),
    .S(_1177_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4167_ (.I0(net63),
    .I1(_1183_),
    .S(_1179_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4168_ (.I0(\mem[5][3] ),
    .I1(net37),
    .S(_1177_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4169_ (.I0(net32),
    .I1(_1184_),
    .S(_1179_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4170_ (.I0(\mem[5][4] ),
    .I1(net48),
    .S(_1177_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4171_ (.I0(net33),
    .I1(_1185_),
    .S(_1179_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4172_ (.I0(\mem[5][5] ),
    .I1(net59),
    .S(_1177_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4173_ (.I0(net34),
    .I1(_1186_),
    .S(_1179_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4174_ (.I0(\mem[5][6] ),
    .I1(net64),
    .S(_1177_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4175_ (.I0(net35),
    .I1(_1187_),
    .S(_1179_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4176_ (.I0(\mem[5][7] ),
    .I1(net65),
    .S(_1177_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4177_ (.I0(net36),
    .I1(_1188_),
    .S(_1179_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4178_ (.I0(\mem[5][8] ),
    .I1(net66),
    .S(_1151_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4179_ (.I0(net38),
    .I1(_1189_),
    .S(_1154_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4180_ (.I0(\mem[5][9] ),
    .I1(net67),
    .S(_1151_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4181_ (.I0(net39),
    .I1(_1190_),
    .S(_1154_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _4182_ (.A1(_2698_),
    .A2(_2714_),
    .A3(_1110_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4183_ (.I(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4184_ (.I0(\mem[6][0] ),
    .I1(net4),
    .S(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4185_ (.A1(_0634_),
    .A2(_0829_),
    .A3(_0743_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4186_ (.I(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4187_ (.I0(net29),
    .I1(_1193_),
    .S(_1195_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4188_ (.I0(\mem[6][10] ),
    .I1(net5),
    .S(_1192_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4189_ (.I0(net40),
    .I1(_1196_),
    .S(_1195_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4190_ (.I0(\mem[6][11] ),
    .I1(net6),
    .S(_1192_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4191_ (.I0(net41),
    .I1(_1197_),
    .S(_1195_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4192_ (.I0(\mem[6][12] ),
    .I1(net7),
    .S(_1192_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4193_ (.I0(net42),
    .I1(_1198_),
    .S(_1195_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4194_ (.I0(\mem[6][13] ),
    .I1(net8),
    .S(_1192_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4195_ (.I0(net43),
    .I1(_1199_),
    .S(_1195_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4196_ (.I0(\mem[6][14] ),
    .I1(net9),
    .S(_1192_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4197_ (.I0(net44),
    .I1(_1200_),
    .S(_1195_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4198_ (.I0(\mem[6][15] ),
    .I1(net10),
    .S(_1192_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4199_ (.I0(net45),
    .I1(_1201_),
    .S(_1195_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4200_ (.I0(\mem[6][16] ),
    .I1(net11),
    .S(_1192_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4201_ (.I0(net46),
    .I1(_1202_),
    .S(_1195_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4202_ (.I0(\mem[6][17] ),
    .I1(net12),
    .S(_1192_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4203_ (.I0(net47),
    .I1(_1203_),
    .S(_1195_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4204_ (.I0(\mem[6][18] ),
    .I1(net13),
    .S(_1192_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4205_ (.I0(net49),
    .I1(_1204_),
    .S(_1195_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4206_ (.I(_1191_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4207_ (.I0(\mem[6][19] ),
    .I1(net14),
    .S(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4208_ (.I(_1194_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4209_ (.I0(net50),
    .I1(_1206_),
    .S(_1207_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4210_ (.I0(\mem[6][1] ),
    .I1(net15),
    .S(_1205_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4211_ (.I0(net30),
    .I1(_1208_),
    .S(_1207_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4212_ (.I0(\mem[6][20] ),
    .I1(net16),
    .S(_1205_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4213_ (.I0(net51),
    .I1(_1209_),
    .S(_1207_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4214_ (.I0(\mem[6][21] ),
    .I1(net17),
    .S(_1205_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4215_ (.I0(net52),
    .I1(_1210_),
    .S(_1207_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4216_ (.I0(\mem[6][22] ),
    .I1(net18),
    .S(_1205_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4217_ (.I0(net53),
    .I1(_1211_),
    .S(_1207_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4218_ (.I0(\mem[6][23] ),
    .I1(net19),
    .S(_1205_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4219_ (.I0(net54),
    .I1(_1212_),
    .S(_1207_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4220_ (.I0(\mem[6][24] ),
    .I1(net20),
    .S(_1205_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4221_ (.I0(net55),
    .I1(_1213_),
    .S(_1207_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4222_ (.I0(\mem[6][25] ),
    .I1(net21),
    .S(_1205_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4223_ (.I0(net56),
    .I1(_1214_),
    .S(_1207_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4224_ (.I0(\mem[6][26] ),
    .I1(net22),
    .S(_1205_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4225_ (.I0(net57),
    .I1(_1215_),
    .S(_1207_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4226_ (.I0(\mem[6][27] ),
    .I1(net23),
    .S(_1205_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4227_ (.I0(net58),
    .I1(_1216_),
    .S(_1207_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4228_ (.I(_1191_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4229_ (.I0(\mem[6][28] ),
    .I1(net24),
    .S(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4230_ (.I(_1194_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4231_ (.I0(net60),
    .I1(_1218_),
    .S(_1219_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4232_ (.I0(\mem[6][29] ),
    .I1(net25),
    .S(_1217_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4233_ (.I0(net61),
    .I1(_1220_),
    .S(_1219_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4234_ (.I0(\mem[6][2] ),
    .I1(net26),
    .S(_1217_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4235_ (.I0(net31),
    .I1(_1221_),
    .S(_1219_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4236_ (.I0(\mem[6][30] ),
    .I1(net27),
    .S(_1217_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4237_ (.I0(net62),
    .I1(_1222_),
    .S(_1219_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4238_ (.I0(\mem[6][31] ),
    .I1(net28),
    .S(_1217_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4239_ (.I0(net63),
    .I1(_1223_),
    .S(_1219_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4240_ (.I0(\mem[6][3] ),
    .I1(net37),
    .S(_1217_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4241_ (.I0(net32),
    .I1(_1224_),
    .S(_1219_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4242_ (.I0(\mem[6][4] ),
    .I1(net48),
    .S(_1217_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4243_ (.I0(net33),
    .I1(_1225_),
    .S(_1219_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4244_ (.I0(\mem[6][5] ),
    .I1(net59),
    .S(_1217_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4245_ (.I0(net34),
    .I1(_1226_),
    .S(_1219_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4246_ (.I0(\mem[6][6] ),
    .I1(net64),
    .S(_1217_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4247_ (.I0(net35),
    .I1(_1227_),
    .S(_1219_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4248_ (.I0(\mem[6][7] ),
    .I1(net65),
    .S(_1217_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4249_ (.I0(net36),
    .I1(_1228_),
    .S(_1219_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4250_ (.I0(\mem[6][8] ),
    .I1(net66),
    .S(_1191_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4251_ (.I0(net38),
    .I1(_1229_),
    .S(_1194_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4252_ (.I0(\mem[6][9] ),
    .I1(net67),
    .S(_1191_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4253_ (.I0(net39),
    .I1(_1230_),
    .S(_1194_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4254_ (.A1(_0635_),
    .A2(_1110_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4255_ (.I(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4256_ (.I0(\mem[7][0] ),
    .I1(net4),
    .S(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4257_ (.A1(_0634_),
    .A2(_0829_),
    .A3(_0787_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4258_ (.I(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4259_ (.I0(net29),
    .I1(_1233_),
    .S(_1235_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4260_ (.I0(\mem[7][10] ),
    .I1(net5),
    .S(_1232_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4261_ (.I0(net40),
    .I1(_1236_),
    .S(_1235_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4262_ (.I0(\mem[7][11] ),
    .I1(net6),
    .S(_1232_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4263_ (.I0(net41),
    .I1(_1237_),
    .S(_1235_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4264_ (.I0(\mem[7][12] ),
    .I1(net7),
    .S(_1232_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4265_ (.I0(net42),
    .I1(_1238_),
    .S(_1235_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4266_ (.I0(\mem[7][13] ),
    .I1(net8),
    .S(_1232_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4267_ (.I0(net43),
    .I1(_1239_),
    .S(_1235_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4268_ (.I0(\mem[7][14] ),
    .I1(net9),
    .S(_1232_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4269_ (.I0(net44),
    .I1(_1240_),
    .S(_1235_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4270_ (.I0(\mem[7][15] ),
    .I1(net10),
    .S(_1232_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4271_ (.I0(net45),
    .I1(_1241_),
    .S(_1235_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4272_ (.I0(\mem[7][16] ),
    .I1(net11),
    .S(_1232_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4273_ (.I0(net46),
    .I1(_1242_),
    .S(_1235_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4274_ (.I0(\mem[7][17] ),
    .I1(net12),
    .S(_1232_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4275_ (.I0(net47),
    .I1(_1243_),
    .S(_1235_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4276_ (.I0(\mem[7][18] ),
    .I1(net13),
    .S(_1232_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4277_ (.I0(net49),
    .I1(_1244_),
    .S(_1235_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4278_ (.I(_1231_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4279_ (.I0(\mem[7][19] ),
    .I1(net14),
    .S(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4280_ (.I(_1234_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4281_ (.I0(net50),
    .I1(_1246_),
    .S(_1247_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4282_ (.I0(\mem[7][1] ),
    .I1(net15),
    .S(_1245_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4283_ (.I0(net30),
    .I1(_1248_),
    .S(_1247_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4284_ (.I0(\mem[7][20] ),
    .I1(net16),
    .S(_1245_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4285_ (.I0(net51),
    .I1(_1249_),
    .S(_1247_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4286_ (.I0(\mem[7][21] ),
    .I1(net17),
    .S(_1245_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4287_ (.I0(net52),
    .I1(_1250_),
    .S(_1247_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4288_ (.I0(\mem[7][22] ),
    .I1(net18),
    .S(_1245_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4289_ (.I0(net53),
    .I1(_1251_),
    .S(_1247_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4290_ (.I0(\mem[7][23] ),
    .I1(net19),
    .S(_1245_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4291_ (.I0(net54),
    .I1(_1252_),
    .S(_1247_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4292_ (.I0(\mem[7][24] ),
    .I1(net20),
    .S(_1245_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4293_ (.I0(net55),
    .I1(_1253_),
    .S(_1247_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4294_ (.I0(\mem[7][25] ),
    .I1(net21),
    .S(_1245_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4295_ (.I0(net56),
    .I1(_1254_),
    .S(_1247_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4296_ (.I0(\mem[7][26] ),
    .I1(net22),
    .S(_1245_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4297_ (.I0(net57),
    .I1(_1255_),
    .S(_1247_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4298_ (.I0(\mem[7][27] ),
    .I1(net23),
    .S(_1245_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4299_ (.I0(net58),
    .I1(_1256_),
    .S(_1247_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4300_ (.I(_1231_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4301_ (.I0(\mem[7][28] ),
    .I1(net24),
    .S(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4302_ (.I(_1234_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4303_ (.I0(net60),
    .I1(_1258_),
    .S(_1259_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4304_ (.I0(\mem[7][29] ),
    .I1(net25),
    .S(_1257_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4305_ (.I0(net61),
    .I1(_1260_),
    .S(_1259_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4306_ (.I0(\mem[7][2] ),
    .I1(net26),
    .S(_1257_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4307_ (.I0(net31),
    .I1(_1261_),
    .S(_1259_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4308_ (.I0(\mem[7][30] ),
    .I1(net27),
    .S(_1257_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4309_ (.I0(net62),
    .I1(_1262_),
    .S(_1259_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4310_ (.I0(\mem[7][31] ),
    .I1(net28),
    .S(_1257_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4311_ (.I0(net63),
    .I1(_1263_),
    .S(_1259_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4312_ (.I0(\mem[7][3] ),
    .I1(net37),
    .S(_1257_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4313_ (.I0(net32),
    .I1(_1264_),
    .S(_1259_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4314_ (.I0(\mem[7][4] ),
    .I1(net48),
    .S(_1257_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4315_ (.I0(net33),
    .I1(_1265_),
    .S(_1259_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4316_ (.I0(\mem[7][5] ),
    .I1(net59),
    .S(_1257_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4317_ (.I0(net34),
    .I1(_1266_),
    .S(_1259_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4318_ (.I0(\mem[7][6] ),
    .I1(net64),
    .S(_1257_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4319_ (.I0(net35),
    .I1(_1267_),
    .S(_1259_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4320_ (.I0(\mem[7][7] ),
    .I1(net65),
    .S(_1257_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4321_ (.I0(net36),
    .I1(_1268_),
    .S(_1259_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4322_ (.I0(\mem[7][8] ),
    .I1(net66),
    .S(_1231_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4323_ (.I0(net38),
    .I1(_1269_),
    .S(_1234_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4324_ (.I0(\mem[7][9] ),
    .I1(net67),
    .S(_1231_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4325_ (.I0(net39),
    .I1(_1270_),
    .S(_1234_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _4326_ (.A1(_2696_),
    .A2(_2714_),
    .A3(_0737_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4327_ (.I(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4328_ (.I0(\mem[8][0] ),
    .I1(net4),
    .S(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4329_ (.A1(_0628_),
    .A2(_0637_),
    .A3(_0745_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4330_ (.I(_1274_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4331_ (.I0(net29),
    .I1(_1273_),
    .S(_1275_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4332_ (.I0(\mem[8][10] ),
    .I1(net5),
    .S(_1272_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4333_ (.I0(net40),
    .I1(_1276_),
    .S(_1275_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4334_ (.I0(\mem[8][11] ),
    .I1(net6),
    .S(_1272_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4335_ (.I0(net41),
    .I1(_1277_),
    .S(_1275_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4336_ (.I0(\mem[8][12] ),
    .I1(net7),
    .S(_1272_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4337_ (.I0(net42),
    .I1(_1278_),
    .S(_1275_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4338_ (.I0(\mem[8][13] ),
    .I1(net8),
    .S(_1272_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4339_ (.I0(net43),
    .I1(_1279_),
    .S(_1275_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4340_ (.I0(\mem[8][14] ),
    .I1(net9),
    .S(_1272_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4341_ (.I0(net44),
    .I1(_1280_),
    .S(_1275_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4342_ (.I0(\mem[8][15] ),
    .I1(net10),
    .S(_1272_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4343_ (.I0(net45),
    .I1(_1281_),
    .S(_1275_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4344_ (.I0(\mem[8][16] ),
    .I1(net11),
    .S(_1272_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4345_ (.I0(net46),
    .I1(_1282_),
    .S(_1275_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4346_ (.I0(\mem[8][17] ),
    .I1(net12),
    .S(_1272_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4347_ (.I0(net47),
    .I1(_1283_),
    .S(_1275_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4348_ (.I0(\mem[8][18] ),
    .I1(net13),
    .S(_1272_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4349_ (.I0(net49),
    .I1(_1284_),
    .S(_1275_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4350_ (.I(_1271_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4351_ (.I0(\mem[8][19] ),
    .I1(net14),
    .S(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4352_ (.I(_1274_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4353_ (.I0(net50),
    .I1(_1286_),
    .S(_1287_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4354_ (.I0(\mem[8][1] ),
    .I1(net15),
    .S(_1285_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4355_ (.I0(net30),
    .I1(_1288_),
    .S(_1287_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4356_ (.I0(\mem[8][20] ),
    .I1(net16),
    .S(_1285_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4357_ (.I0(net51),
    .I1(_1289_),
    .S(_1287_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4358_ (.I0(\mem[8][21] ),
    .I1(net17),
    .S(_1285_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4359_ (.I0(net52),
    .I1(_1290_),
    .S(_1287_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4360_ (.I0(\mem[8][22] ),
    .I1(net18),
    .S(_1285_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4361_ (.I0(net53),
    .I1(_1291_),
    .S(_1287_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4362_ (.I0(\mem[8][23] ),
    .I1(net19),
    .S(_1285_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4363_ (.I0(net54),
    .I1(_1292_),
    .S(_1287_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4364_ (.I0(\mem[8][24] ),
    .I1(net20),
    .S(_1285_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4365_ (.I0(net55),
    .I1(_1293_),
    .S(_1287_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4366_ (.I0(\mem[8][25] ),
    .I1(net21),
    .S(_1285_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4367_ (.I0(net56),
    .I1(_1294_),
    .S(_1287_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4368_ (.I0(\mem[8][26] ),
    .I1(net22),
    .S(_1285_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4369_ (.I0(net57),
    .I1(_1295_),
    .S(_1287_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4370_ (.I0(\mem[8][27] ),
    .I1(net23),
    .S(_1285_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4371_ (.I0(net58),
    .I1(_1296_),
    .S(_1287_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4372_ (.I(_1271_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4373_ (.I0(\mem[8][28] ),
    .I1(net24),
    .S(_1297_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4374_ (.I(_1274_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4375_ (.I0(net60),
    .I1(_1298_),
    .S(_1299_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4376_ (.I0(\mem[8][29] ),
    .I1(net25),
    .S(_1297_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4377_ (.I0(net61),
    .I1(_1300_),
    .S(_1299_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4378_ (.I0(\mem[8][2] ),
    .I1(net26),
    .S(_1297_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4379_ (.I0(net31),
    .I1(_1301_),
    .S(_1299_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4380_ (.I0(\mem[8][30] ),
    .I1(net27),
    .S(_1297_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4381_ (.I0(net62),
    .I1(_1302_),
    .S(_1299_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4382_ (.I0(\mem[8][31] ),
    .I1(net28),
    .S(_1297_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4383_ (.I0(net63),
    .I1(_1303_),
    .S(_1299_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4384_ (.I0(\mem[8][3] ),
    .I1(net37),
    .S(_1297_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4385_ (.I0(net32),
    .I1(_1304_),
    .S(_1299_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4386_ (.I0(\mem[8][4] ),
    .I1(net48),
    .S(_1297_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4387_ (.I0(net33),
    .I1(_1305_),
    .S(_1299_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4388_ (.I0(\mem[8][5] ),
    .I1(net59),
    .S(_1297_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4389_ (.I0(net34),
    .I1(_1306_),
    .S(_1299_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4390_ (.I0(\mem[8][6] ),
    .I1(net64),
    .S(_1297_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4391_ (.I0(net35),
    .I1(_1307_),
    .S(_1299_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4392_ (.I0(\mem[8][7] ),
    .I1(net65),
    .S(_1297_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4393_ (.I0(net36),
    .I1(_1308_),
    .S(_1299_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4394_ (.I0(\mem[8][8] ),
    .I1(net66),
    .S(_1271_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4395_ (.I0(net38),
    .I1(_1309_),
    .S(_1274_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4396_ (.I0(\mem[8][9] ),
    .I1(net67),
    .S(_1271_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4397_ (.I0(net39),
    .I1(_1310_),
    .S(_1274_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _4398_ (.A1(_2700_),
    .A2(_0596_),
    .A3(_0737_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4399_ (.I(_1311_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4400_ (.I0(\mem[9][0] ),
    .I1(net4),
    .S(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4401_ (.A1(_0637_),
    .A2(_0745_),
    .A3(_0872_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4402_ (.I(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4403_ (.I0(net29),
    .I1(_1313_),
    .S(_1315_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4404_ (.I0(\mem[9][10] ),
    .I1(net5),
    .S(_1312_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4405_ (.I0(net40),
    .I1(_1316_),
    .S(_1315_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4406_ (.I0(\mem[9][11] ),
    .I1(net6),
    .S(_1312_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4407_ (.I0(net41),
    .I1(_1317_),
    .S(_1315_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4408_ (.I0(\mem[9][12] ),
    .I1(net7),
    .S(_1312_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4409_ (.I0(net42),
    .I1(_1318_),
    .S(_1315_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4410_ (.I0(\mem[9][13] ),
    .I1(net8),
    .S(_1312_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4411_ (.I0(net43),
    .I1(_1319_),
    .S(_1315_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4412_ (.I0(\mem[9][14] ),
    .I1(net9),
    .S(_1312_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4413_ (.I0(net44),
    .I1(_1320_),
    .S(_1315_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4414_ (.I0(\mem[9][15] ),
    .I1(net10),
    .S(_1312_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4415_ (.I0(net45),
    .I1(_1321_),
    .S(_1315_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4416_ (.I0(\mem[9][16] ),
    .I1(net11),
    .S(_1312_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4417_ (.I0(net46),
    .I1(_1322_),
    .S(_1315_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4418_ (.I0(\mem[9][17] ),
    .I1(net12),
    .S(_1312_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4419_ (.I0(net47),
    .I1(_1323_),
    .S(_1315_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4420_ (.I0(\mem[9][18] ),
    .I1(net13),
    .S(_1312_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4421_ (.I0(net49),
    .I1(_1324_),
    .S(_1315_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4422_ (.I(_1311_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4423_ (.I0(\mem[9][19] ),
    .I1(net14),
    .S(_1325_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4424_ (.I(_1314_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4425_ (.I0(net50),
    .I1(_1326_),
    .S(_1327_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4426_ (.I0(\mem[9][1] ),
    .I1(net15),
    .S(_1325_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4427_ (.I0(net30),
    .I1(_1328_),
    .S(_1327_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4428_ (.I0(\mem[9][20] ),
    .I1(net16),
    .S(_1325_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4429_ (.I0(net51),
    .I1(_1329_),
    .S(_1327_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4430_ (.I0(\mem[9][21] ),
    .I1(net17),
    .S(_1325_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4431_ (.I0(net52),
    .I1(_1330_),
    .S(_1327_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4432_ (.I0(\mem[9][22] ),
    .I1(net18),
    .S(_1325_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4433_ (.I0(net53),
    .I1(_1331_),
    .S(_1327_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4434_ (.I0(\mem[9][23] ),
    .I1(net19),
    .S(_1325_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4435_ (.I0(net54),
    .I1(_1332_),
    .S(_1327_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4436_ (.I0(\mem[9][24] ),
    .I1(net20),
    .S(_1325_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4437_ (.I0(net55),
    .I1(_1333_),
    .S(_1327_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4438_ (.I0(\mem[9][25] ),
    .I1(net21),
    .S(_1325_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4439_ (.I0(net56),
    .I1(_1334_),
    .S(_1327_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4440_ (.I0(\mem[9][26] ),
    .I1(net22),
    .S(_1325_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4441_ (.I0(net57),
    .I1(_1335_),
    .S(_1327_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4442_ (.I0(\mem[9][27] ),
    .I1(net23),
    .S(_1325_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4443_ (.I0(net58),
    .I1(_1336_),
    .S(_1327_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4444_ (.I(_1311_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4445_ (.I0(\mem[9][28] ),
    .I1(net24),
    .S(_1337_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4446_ (.I(_1314_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4447_ (.I0(net60),
    .I1(_1338_),
    .S(_1339_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4448_ (.I0(\mem[9][29] ),
    .I1(net25),
    .S(_1337_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4449_ (.I0(net61),
    .I1(_1340_),
    .S(_1339_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4450_ (.I0(\mem[9][2] ),
    .I1(net26),
    .S(_1337_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4451_ (.I0(net31),
    .I1(_1341_),
    .S(_1339_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4452_ (.I0(\mem[9][30] ),
    .I1(net27),
    .S(_1337_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4453_ (.I0(net62),
    .I1(_1342_),
    .S(_1339_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4454_ (.I0(\mem[9][31] ),
    .I1(net28),
    .S(_1337_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4455_ (.I0(net63),
    .I1(_1343_),
    .S(_1339_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4456_ (.I0(\mem[9][3] ),
    .I1(net37),
    .S(_1337_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4457_ (.I0(net32),
    .I1(_1344_),
    .S(_1339_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4458_ (.I0(\mem[9][4] ),
    .I1(net48),
    .S(_1337_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4459_ (.I0(net33),
    .I1(_1345_),
    .S(_1339_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4460_ (.I0(\mem[9][5] ),
    .I1(net59),
    .S(_1337_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4461_ (.I0(net34),
    .I1(_1346_),
    .S(_1339_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4462_ (.I0(\mem[9][6] ),
    .I1(net64),
    .S(_1337_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4463_ (.I0(net35),
    .I1(_1347_),
    .S(_1339_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4464_ (.I0(\mem[9][7] ),
    .I1(net65),
    .S(_1337_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4465_ (.I0(net36),
    .I1(_1348_),
    .S(_1339_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4466_ (.I0(\mem[9][8] ),
    .I1(net66),
    .S(_1311_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4467_ (.I0(net38),
    .I1(_1349_),
    .S(_1314_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4468_ (.I0(\mem[9][9] ),
    .I1(net67),
    .S(_1311_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4469_ (.I0(net39),
    .I1(_1350_),
    .S(_1314_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4470_ (.I(_0612_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4471_ (.I0(\mem[4][0] ),
    .I1(\mem[6][0] ),
    .S(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4472_ (.I(_0613_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4473_ (.I0(\mem[5][0] ),
    .I1(\mem[7][0] ),
    .S(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4474_ (.I(\rd_ptr[1] ),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4475_ (.I(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4476_ (.I0(\mem[12][0] ),
    .I1(\mem[14][0] ),
    .S(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4477_ (.I(_0612_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4478_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4479_ (.I0(\mem[13][0] ),
    .I1(\mem[15][0] ),
    .S(_1359_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4480_ (.I(\rd_ptr[0] ),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4481_ (.I(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4482_ (.I(\rd_ptr[3] ),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4483_ (.I(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4484_ (.I0(_1352_),
    .I1(_1354_),
    .I2(_1357_),
    .I3(_1360_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4485_ (.I0(\mem[0][0] ),
    .I1(\mem[2][0] ),
    .S(_1355_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4486_ (.I(_0612_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4487_ (.I0(\mem[1][0] ),
    .I1(\mem[3][0] ),
    .S(_1367_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4488_ (.I0(\mem[8][0] ),
    .I1(\mem[10][0] ),
    .S(_1353_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4489_ (.I(_1358_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4490_ (.I0(\mem[9][0] ),
    .I1(\mem[11][0] ),
    .S(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4491_ (.I(_1361_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4492_ (.I(_1363_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4493_ (.I0(_1366_),
    .I1(_1368_),
    .I2(_1369_),
    .I3(_1371_),
    .S0(_1372_),
    .S1(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _4494_ (.I(\rd_ptr[2] ),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4495_ (.I(_1375_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4496_ (.I(_1376_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4497_ (.I(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4498_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4499_ (.I0(_1365_),
    .I1(_1374_),
    .S(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4500_ (.I0(net79),
    .I1(_1380_),
    .S(_0001_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4501_ (.I(\rd_ptr[1] ),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4502_ (.I(_1381_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4503_ (.I0(\mem[4][10] ),
    .I1(\mem[6][10] ),
    .S(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4504_ (.I0(\mem[5][10] ),
    .I1(\mem[7][10] ),
    .S(_1353_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4505_ (.I0(\mem[12][10] ),
    .I1(\mem[14][10] ),
    .S(_1381_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4506_ (.I(_0613_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4507_ (.I0(\mem[13][10] ),
    .I1(\mem[15][10] ),
    .S(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4508_ (.I0(_1383_),
    .I1(_1384_),
    .I2(_1385_),
    .I3(_1387_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4509_ (.I(_0613_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4510_ (.I0(\mem[1][10] ),
    .I1(\mem[3][10] ),
    .S(_1389_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4511_ (.I(_0613_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4512_ (.I0(\mem[0][10] ),
    .I1(\mem[2][10] ),
    .S(_1391_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4513_ (.I0(\mem[9][10] ),
    .I1(\mem[11][10] ),
    .S(_1367_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4514_ (.I0(\mem[8][10] ),
    .I1(\mem[10][10] ),
    .S(_1358_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _4515_ (.I(_1361_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4516_ (.I(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4517_ (.I0(_1390_),
    .I1(_1392_),
    .I2(_1393_),
    .I3(_1394_),
    .S0(_1396_),
    .S1(_1373_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4518_ (.I0(_1388_),
    .I1(_1397_),
    .S(_1379_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4519_ (.I0(net80),
    .I1(_1398_),
    .S(_0001_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4520_ (.I0(\mem[4][11] ),
    .I1(\mem[6][11] ),
    .S(_1382_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4521_ (.I(_0613_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4522_ (.I0(\mem[5][11] ),
    .I1(\mem[7][11] ),
    .S(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4523_ (.I0(\mem[12][11] ),
    .I1(\mem[14][11] ),
    .S(_1381_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4524_ (.I0(\mem[13][11] ),
    .I1(\mem[15][11] ),
    .S(_1386_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4525_ (.I0(_1399_),
    .I1(_1401_),
    .I2(_1402_),
    .I3(_1403_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4526_ (.I(_1381_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4527_ (.I0(\mem[1][11] ),
    .I1(\mem[3][11] ),
    .S(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4528_ (.I0(\mem[0][11] ),
    .I1(\mem[2][11] ),
    .S(_1391_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4529_ (.I0(\mem[9][11] ),
    .I1(\mem[11][11] ),
    .S(_1367_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4530_ (.I0(\mem[8][11] ),
    .I1(\mem[10][11] ),
    .S(_1358_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4531_ (.I0(_1406_),
    .I1(_1407_),
    .I2(_1408_),
    .I3(_1409_),
    .S0(_1396_),
    .S1(_1373_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4532_ (.I0(_1404_),
    .I1(_1410_),
    .S(_1379_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4533_ (.I0(net81),
    .I1(_1411_),
    .S(_0001_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4534_ (.I0(\mem[4][12] ),
    .I1(\mem[6][12] ),
    .S(_1382_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4535_ (.I0(\mem[5][12] ),
    .I1(\mem[7][12] ),
    .S(_1400_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4536_ (.I0(\mem[12][12] ),
    .I1(\mem[14][12] ),
    .S(_1381_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4537_ (.I0(\mem[13][12] ),
    .I1(\mem[15][12] ),
    .S(_1386_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4538_ (.I0(_1412_),
    .I1(_1413_),
    .I2(_1414_),
    .I3(_1415_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4539_ (.I0(\mem[1][12] ),
    .I1(\mem[3][12] ),
    .S(_1405_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4540_ (.I0(\mem[0][12] ),
    .I1(\mem[2][12] ),
    .S(_1391_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4541_ (.I0(\mem[9][12] ),
    .I1(\mem[11][12] ),
    .S(_1367_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4542_ (.I0(\mem[8][12] ),
    .I1(\mem[10][12] ),
    .S(_1358_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4543_ (.I0(_1417_),
    .I1(_1418_),
    .I2(_1419_),
    .I3(_1420_),
    .S0(_1396_),
    .S1(_1373_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4544_ (.I0(_1416_),
    .I1(_1421_),
    .S(_1379_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4545_ (.I0(net82),
    .I1(_1422_),
    .S(_0001_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4546_ (.I0(\mem[4][13] ),
    .I1(\mem[6][13] ),
    .S(_1382_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4547_ (.I0(\mem[5][13] ),
    .I1(\mem[7][13] ),
    .S(_1400_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4548_ (.I0(\mem[12][13] ),
    .I1(\mem[14][13] ),
    .S(_1381_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4549_ (.I0(\mem[13][13] ),
    .I1(\mem[15][13] ),
    .S(_1386_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4550_ (.I0(_1423_),
    .I1(_1424_),
    .I2(_1425_),
    .I3(_1426_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4551_ (.I0(\mem[1][13] ),
    .I1(\mem[3][13] ),
    .S(_1405_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4552_ (.I0(\mem[0][13] ),
    .I1(\mem[2][13] ),
    .S(_1391_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4553_ (.I0(\mem[9][13] ),
    .I1(\mem[11][13] ),
    .S(_1367_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4554_ (.I0(\mem[8][13] ),
    .I1(\mem[10][13] ),
    .S(_1358_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4555_ (.I0(_1428_),
    .I1(_1429_),
    .I2(_1430_),
    .I3(_1431_),
    .S0(_1396_),
    .S1(_1373_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4556_ (.I0(_1427_),
    .I1(_1432_),
    .S(_1379_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4557_ (.I0(net83),
    .I1(_1433_),
    .S(_0001_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4558_ (.I0(\mem[4][14] ),
    .I1(\mem[6][14] ),
    .S(_1382_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4559_ (.I0(\mem[5][14] ),
    .I1(\mem[7][14] ),
    .S(_1400_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4560_ (.I0(\mem[12][14] ),
    .I1(\mem[14][14] ),
    .S(_1381_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4561_ (.I0(\mem[13][14] ),
    .I1(\mem[15][14] ),
    .S(_1386_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4562_ (.I0(_1434_),
    .I1(_1435_),
    .I2(_1436_),
    .I3(_1437_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4563_ (.I0(\mem[1][14] ),
    .I1(\mem[3][14] ),
    .S(_1405_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4564_ (.I(_0613_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4565_ (.I0(\mem[0][14] ),
    .I1(\mem[2][14] ),
    .S(_1440_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4566_ (.I0(\mem[9][14] ),
    .I1(\mem[11][14] ),
    .S(_1367_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4567_ (.I0(\mem[8][14] ),
    .I1(\mem[10][14] ),
    .S(_1358_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4568_ (.I(_1395_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4569_ (.I0(_1439_),
    .I1(_1441_),
    .I2(_1442_),
    .I3(_1443_),
    .S0(_1444_),
    .S1(_1373_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4570_ (.I0(_1438_),
    .I1(_1445_),
    .S(_1379_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4571_ (.I0(net84),
    .I1(_1446_),
    .S(_0001_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4572_ (.I0(\mem[4][15] ),
    .I1(\mem[6][15] ),
    .S(_1382_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4573_ (.I0(\mem[5][15] ),
    .I1(\mem[7][15] ),
    .S(_1400_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4574_ (.I0(\mem[12][15] ),
    .I1(\mem[14][15] ),
    .S(_1381_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4575_ (.I0(\mem[13][15] ),
    .I1(\mem[15][15] ),
    .S(_1386_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4576_ (.I0(_1447_),
    .I1(_1448_),
    .I2(_1449_),
    .I3(_1450_),
    .S0(_1362_),
    .S1(_1364_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4577_ (.I0(\mem[1][15] ),
    .I1(\mem[3][15] ),
    .S(_1405_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4578_ (.I0(\mem[0][15] ),
    .I1(\mem[2][15] ),
    .S(_1440_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4579_ (.I(_0612_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4580_ (.I0(\mem[9][15] ),
    .I1(\mem[11][15] ),
    .S(_1454_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4581_ (.I0(\mem[8][15] ),
    .I1(\mem[10][15] ),
    .S(_1358_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4582_ (.I0(_1452_),
    .I1(_1453_),
    .I2(_1455_),
    .I3(_1456_),
    .S0(_1444_),
    .S1(_1373_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4583_ (.I0(_1451_),
    .I1(_1457_),
    .S(_1379_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4584_ (.I0(net85),
    .I1(_1458_),
    .S(_0001_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4585_ (.I(_1381_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4586_ (.I0(\mem[4][16] ),
    .I1(\mem[6][16] ),
    .S(_1459_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4587_ (.I0(\mem[5][16] ),
    .I1(\mem[7][16] ),
    .S(_1400_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4588_ (.I(_0612_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4589_ (.I0(\mem[12][16] ),
    .I1(\mem[14][16] ),
    .S(_1462_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4590_ (.I(_0613_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4591_ (.I0(\mem[13][16] ),
    .I1(\mem[15][16] ),
    .S(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4592_ (.I(_1361_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4593_ (.I0(_1460_),
    .I1(_1461_),
    .I2(_1463_),
    .I3(_1465_),
    .S0(_1466_),
    .S1(_1364_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4594_ (.I0(\mem[1][16] ),
    .I1(\mem[3][16] ),
    .S(_1405_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4595_ (.I0(\mem[0][16] ),
    .I1(\mem[2][16] ),
    .S(_1440_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4596_ (.I0(\mem[9][16] ),
    .I1(\mem[11][16] ),
    .S(_1454_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4597_ (.I0(\mem[8][16] ),
    .I1(\mem[10][16] ),
    .S(_1358_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4598_ (.I(_1363_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4599_ (.I0(_1468_),
    .I1(_1469_),
    .I2(_1470_),
    .I3(_1471_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4600_ (.I0(_1467_),
    .I1(_1473_),
    .S(_1379_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4601_ (.I0(net86),
    .I1(_1474_),
    .S(_0001_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4602_ (.I0(\mem[4][17] ),
    .I1(\mem[6][17] ),
    .S(_1459_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4603_ (.I0(\mem[5][17] ),
    .I1(\mem[7][17] ),
    .S(_1400_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4604_ (.I0(\mem[12][17] ),
    .I1(\mem[14][17] ),
    .S(_1462_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4605_ (.I0(\mem[13][17] ),
    .I1(\mem[15][17] ),
    .S(_1464_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4606_ (.I0(_1475_),
    .I1(_1476_),
    .I2(_1477_),
    .I3(_1478_),
    .S0(_1466_),
    .S1(_1364_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4607_ (.I0(\mem[1][17] ),
    .I1(\mem[3][17] ),
    .S(_1405_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4608_ (.I0(\mem[0][17] ),
    .I1(\mem[2][17] ),
    .S(_1440_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4609_ (.I0(\mem[9][17] ),
    .I1(\mem[11][17] ),
    .S(_1454_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4610_ (.I0(\mem[8][17] ),
    .I1(\mem[10][17] ),
    .S(_1358_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4611_ (.I0(_1480_),
    .I1(_1481_),
    .I2(_1482_),
    .I3(_1483_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4612_ (.I0(_1479_),
    .I1(_1484_),
    .S(_1379_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4613_ (.I0(net87),
    .I1(_1485_),
    .S(_0001_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4614_ (.I0(\mem[4][18] ),
    .I1(\mem[6][18] ),
    .S(_1459_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4615_ (.I0(\mem[5][18] ),
    .I1(\mem[7][18] ),
    .S(_1400_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4616_ (.I0(\mem[12][18] ),
    .I1(\mem[14][18] ),
    .S(_1462_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4617_ (.I0(\mem[13][18] ),
    .I1(\mem[15][18] ),
    .S(_1464_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4618_ (.I(_1363_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4619_ (.I0(_1486_),
    .I1(_1487_),
    .I2(_1488_),
    .I3(_1489_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4620_ (.I0(\mem[1][18] ),
    .I1(\mem[3][18] ),
    .S(_1405_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4621_ (.I0(\mem[0][18] ),
    .I1(\mem[2][18] ),
    .S(_1440_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4622_ (.I0(\mem[9][18] ),
    .I1(\mem[11][18] ),
    .S(_1454_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4623_ (.I(_0612_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4624_ (.I0(\mem[8][18] ),
    .I1(\mem[10][18] ),
    .S(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4625_ (.I0(_1492_),
    .I1(_1493_),
    .I2(_1494_),
    .I3(_1496_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4626_ (.I(_1378_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4627_ (.I0(_1491_),
    .I1(_1497_),
    .S(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4628_ (.I(_0604_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4629_ (.I0(net88),
    .I1(_1499_),
    .S(_1500_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4630_ (.I0(\mem[4][19] ),
    .I1(\mem[6][19] ),
    .S(_1459_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4631_ (.I0(\mem[5][19] ),
    .I1(\mem[7][19] ),
    .S(_1400_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4632_ (.I0(\mem[12][19] ),
    .I1(\mem[14][19] ),
    .S(_1462_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4633_ (.I0(\mem[13][19] ),
    .I1(\mem[15][19] ),
    .S(_1464_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4634_ (.I0(_1501_),
    .I1(_1502_),
    .I2(_1503_),
    .I3(_1504_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4635_ (.I0(\mem[1][19] ),
    .I1(\mem[3][19] ),
    .S(_1405_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4636_ (.I0(\mem[0][19] ),
    .I1(\mem[2][19] ),
    .S(_1440_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4637_ (.I0(\mem[9][19] ),
    .I1(\mem[11][19] ),
    .S(_1454_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4638_ (.I0(\mem[8][19] ),
    .I1(\mem[10][19] ),
    .S(_1495_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4639_ (.I0(_1506_),
    .I1(_1507_),
    .I2(_1508_),
    .I3(_1509_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4640_ (.I0(_1505_),
    .I1(_1510_),
    .S(_1498_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4641_ (.I0(net89),
    .I1(_1511_),
    .S(_1500_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4642_ (.I0(\mem[4][1] ),
    .I1(\mem[6][1] ),
    .S(_1459_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4643_ (.I0(\mem[5][1] ),
    .I1(\mem[7][1] ),
    .S(_1400_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4644_ (.I0(\mem[12][1] ),
    .I1(\mem[14][1] ),
    .S(_1462_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4645_ (.I0(\mem[13][1] ),
    .I1(\mem[15][1] ),
    .S(_1464_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4646_ (.I0(_1512_),
    .I1(_1513_),
    .I2(_1514_),
    .I3(_1515_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4647_ (.I0(\mem[1][1] ),
    .I1(\mem[3][1] ),
    .S(_1405_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4648_ (.I0(\mem[0][1] ),
    .I1(\mem[2][1] ),
    .S(_1440_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4649_ (.I0(\mem[9][1] ),
    .I1(\mem[11][1] ),
    .S(_1454_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4650_ (.I0(\mem[8][1] ),
    .I1(\mem[10][1] ),
    .S(_1495_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4651_ (.I0(_1517_),
    .I1(_1518_),
    .I2(_1519_),
    .I3(_1520_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4652_ (.I0(_1516_),
    .I1(_1521_),
    .S(_1498_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4653_ (.I0(net90),
    .I1(_1522_),
    .S(_1500_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4654_ (.I(_1355_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4655_ (.I0(\mem[5][20] ),
    .I1(\mem[7][20] ),
    .S(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4656_ (.I(_0612_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4657_ (.I0(\mem[4][20] ),
    .I1(\mem[6][20] ),
    .S(_1525_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4658_ (.I0(\mem[13][20] ),
    .I1(\mem[15][20] ),
    .S(_1356_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4659_ (.I0(\mem[12][20] ),
    .I1(\mem[14][20] ),
    .S(_1359_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4660_ (.I0(_1524_),
    .I1(_1526_),
    .I2(_1527_),
    .I3(_1528_),
    .S0(_1396_),
    .S1(_1490_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4661_ (.I0(\mem[0][20] ),
    .I1(\mem[2][20] ),
    .S(_1525_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4662_ (.I0(\mem[1][20] ),
    .I1(\mem[3][20] ),
    .S(_1523_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4663_ (.I0(\mem[8][20] ),
    .I1(\mem[10][20] ),
    .S(_1353_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4664_ (.I0(\mem[9][20] ),
    .I1(\mem[11][20] ),
    .S(_1359_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4665_ (.I(_1361_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4666_ (.I0(_1530_),
    .I1(_1531_),
    .I2(_1532_),
    .I3(_1533_),
    .S0(_1534_),
    .S1(_1472_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4667_ (.I0(_1529_),
    .I1(_1535_),
    .S(_1498_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4668_ (.I0(net91),
    .I1(_1536_),
    .S(_1500_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4669_ (.I0(\mem[4][21] ),
    .I1(\mem[6][21] ),
    .S(_1459_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4670_ (.I(_0613_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4671_ (.I0(\mem[5][21] ),
    .I1(\mem[7][21] ),
    .S(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4672_ (.I0(\mem[12][21] ),
    .I1(\mem[14][21] ),
    .S(_1462_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4673_ (.I0(\mem[13][21] ),
    .I1(\mem[15][21] ),
    .S(_1464_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4674_ (.I0(_1537_),
    .I1(_1539_),
    .I2(_1540_),
    .I3(_1541_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4675_ (.I(_1381_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4676_ (.I0(\mem[1][21] ),
    .I1(\mem[3][21] ),
    .S(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4677_ (.I0(\mem[0][21] ),
    .I1(\mem[2][21] ),
    .S(_1440_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4678_ (.I0(\mem[9][21] ),
    .I1(\mem[11][21] ),
    .S(_1454_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4679_ (.I0(\mem[8][21] ),
    .I1(\mem[10][21] ),
    .S(_1495_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4680_ (.I0(_1544_),
    .I1(_1545_),
    .I2(_1546_),
    .I3(_1547_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4681_ (.I0(_1542_),
    .I1(_1548_),
    .S(_1498_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4682_ (.I0(net92),
    .I1(_1549_),
    .S(_1500_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4683_ (.I0(\mem[5][22] ),
    .I1(\mem[7][22] ),
    .S(_1523_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4684_ (.I0(\mem[4][22] ),
    .I1(\mem[6][22] ),
    .S(_1525_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4685_ (.I0(\mem[13][22] ),
    .I1(\mem[15][22] ),
    .S(_1356_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4686_ (.I0(\mem[12][22] ),
    .I1(\mem[14][22] ),
    .S(_1359_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4687_ (.I0(_1550_),
    .I1(_1551_),
    .I2(_1552_),
    .I3(_1553_),
    .S0(_1396_),
    .S1(_1490_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4688_ (.I0(\mem[0][22] ),
    .I1(\mem[2][22] ),
    .S(_1525_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4689_ (.I0(\mem[1][22] ),
    .I1(\mem[3][22] ),
    .S(_1523_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4690_ (.I0(\mem[8][22] ),
    .I1(\mem[10][22] ),
    .S(_1353_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4691_ (.I0(\mem[9][22] ),
    .I1(\mem[11][22] ),
    .S(_1359_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4692_ (.I0(_1555_),
    .I1(_1556_),
    .I2(_1557_),
    .I3(_1558_),
    .S0(_1534_),
    .S1(_1472_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4693_ (.I0(_1554_),
    .I1(_1559_),
    .S(_1498_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4694_ (.I0(net93),
    .I1(_1560_),
    .S(_1500_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4695_ (.I0(\mem[4][23] ),
    .I1(\mem[6][23] ),
    .S(_1459_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4696_ (.I0(\mem[5][23] ),
    .I1(\mem[7][23] ),
    .S(_1538_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4697_ (.I0(\mem[12][23] ),
    .I1(\mem[14][23] ),
    .S(_1462_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4698_ (.I0(\mem[13][23] ),
    .I1(\mem[15][23] ),
    .S(_1464_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4699_ (.I0(_1561_),
    .I1(_1562_),
    .I2(_1563_),
    .I3(_1564_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4700_ (.I0(\mem[1][23] ),
    .I1(\mem[3][23] ),
    .S(_1543_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4701_ (.I0(\mem[0][23] ),
    .I1(\mem[2][23] ),
    .S(_1440_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4702_ (.I0(\mem[9][23] ),
    .I1(\mem[11][23] ),
    .S(_1454_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4703_ (.I0(\mem[8][23] ),
    .I1(\mem[10][23] ),
    .S(_1495_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4704_ (.I0(_1566_),
    .I1(_1567_),
    .I2(_1568_),
    .I3(_1569_),
    .S0(_1444_),
    .S1(_1472_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4705_ (.I0(_1565_),
    .I1(_1570_),
    .S(_1498_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4706_ (.I0(net94),
    .I1(_1571_),
    .S(_1500_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4707_ (.I0(\mem[5][24] ),
    .I1(\mem[7][24] ),
    .S(_1523_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4708_ (.I0(\mem[4][24] ),
    .I1(\mem[6][24] ),
    .S(_1525_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4709_ (.I0(\mem[13][24] ),
    .I1(\mem[15][24] ),
    .S(_1356_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4710_ (.I0(\mem[12][24] ),
    .I1(\mem[14][24] ),
    .S(_1359_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4711_ (.I0(_1572_),
    .I1(_1573_),
    .I2(_1574_),
    .I3(_1575_),
    .S0(_1396_),
    .S1(_1490_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4712_ (.I0(\mem[0][24] ),
    .I1(\mem[2][24] ),
    .S(_1367_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4713_ (.I0(\mem[1][24] ),
    .I1(\mem[3][24] ),
    .S(_1523_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4714_ (.I0(\mem[8][24] ),
    .I1(\mem[10][24] ),
    .S(_1353_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4715_ (.I0(\mem[9][24] ),
    .I1(\mem[11][24] ),
    .S(_1359_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4716_ (.I0(_1577_),
    .I1(_1578_),
    .I2(_1579_),
    .I3(_1580_),
    .S0(_1534_),
    .S1(_1472_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4717_ (.I0(_1576_),
    .I1(_1581_),
    .S(_1498_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4718_ (.I0(net95),
    .I1(_1582_),
    .S(_1500_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4719_ (.I0(\mem[4][25] ),
    .I1(\mem[6][25] ),
    .S(_1459_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4720_ (.I0(\mem[5][25] ),
    .I1(\mem[7][25] ),
    .S(_1538_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4721_ (.I0(\mem[12][25] ),
    .I1(\mem[14][25] ),
    .S(_1462_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4722_ (.I0(\mem[13][25] ),
    .I1(\mem[15][25] ),
    .S(_1464_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4723_ (.I0(_1583_),
    .I1(_1584_),
    .I2(_1585_),
    .I3(_1586_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4724_ (.I0(\mem[1][25] ),
    .I1(\mem[3][25] ),
    .S(_1543_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4725_ (.I0(\mem[0][25] ),
    .I1(\mem[2][25] ),
    .S(_1440_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4726_ (.I0(\mem[9][25] ),
    .I1(\mem[11][25] ),
    .S(_1454_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4727_ (.I0(\mem[8][25] ),
    .I1(\mem[10][25] ),
    .S(_1495_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4728_ (.I(\rd_ptr[3] ),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4729_ (.I0(_1588_),
    .I1(_1589_),
    .I2(_1590_),
    .I3(_1591_),
    .S0(_1444_),
    .S1(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4730_ (.I0(_1587_),
    .I1(_1593_),
    .S(_1498_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4731_ (.I0(net96),
    .I1(_1594_),
    .S(_1500_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4732_ (.I0(\mem[4][26] ),
    .I1(\mem[6][26] ),
    .S(_1459_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4733_ (.I0(\mem[5][26] ),
    .I1(\mem[7][26] ),
    .S(_1538_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4734_ (.I0(\mem[12][26] ),
    .I1(\mem[14][26] ),
    .S(_1462_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4735_ (.I0(\mem[13][26] ),
    .I1(\mem[15][26] ),
    .S(_1464_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4736_ (.I0(_1595_),
    .I1(_1596_),
    .I2(_1597_),
    .I3(_1598_),
    .S0(_1466_),
    .S1(_1490_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4737_ (.I0(\mem[1][26] ),
    .I1(\mem[3][26] ),
    .S(_1543_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4738_ (.I(_0613_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4739_ (.I0(\mem[0][26] ),
    .I1(\mem[2][26] ),
    .S(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4740_ (.I0(\mem[9][26] ),
    .I1(\mem[11][26] ),
    .S(_1454_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4741_ (.I0(\mem[8][26] ),
    .I1(\mem[10][26] ),
    .S(_1495_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4742_ (.I(_1395_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4743_ (.I0(_1600_),
    .I1(_1602_),
    .I2(_1603_),
    .I3(_1604_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4744_ (.I0(_1599_),
    .I1(_1606_),
    .S(_1498_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4745_ (.I0(net97),
    .I1(_1607_),
    .S(_1500_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4746_ (.I0(\mem[4][27] ),
    .I1(\mem[6][27] ),
    .S(_1459_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4747_ (.I0(\mem[5][27] ),
    .I1(\mem[7][27] ),
    .S(_1538_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4748_ (.I0(\mem[12][27] ),
    .I1(\mem[14][27] ),
    .S(_1462_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4749_ (.I0(\mem[13][27] ),
    .I1(\mem[15][27] ),
    .S(_1464_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4750_ (.I(_1363_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4751_ (.I0(_1608_),
    .I1(_1609_),
    .I2(_1610_),
    .I3(_1611_),
    .S0(_1466_),
    .S1(_1612_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4752_ (.I0(\mem[1][27] ),
    .I1(\mem[3][27] ),
    .S(_1543_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4753_ (.I0(\mem[0][27] ),
    .I1(\mem[2][27] ),
    .S(_1601_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4754_ (.I(_0612_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4755_ (.I0(\mem[9][27] ),
    .I1(\mem[11][27] ),
    .S(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4756_ (.I0(\mem[8][27] ),
    .I1(\mem[10][27] ),
    .S(_1495_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4757_ (.I0(_1614_),
    .I1(_1615_),
    .I2(_1617_),
    .I3(_1618_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4758_ (.I(_1378_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4759_ (.I0(_1613_),
    .I1(_1619_),
    .S(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4760_ (.I(_0604_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4761_ (.I0(net98),
    .I1(_1621_),
    .S(_1622_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4762_ (.I0(\mem[4][28] ),
    .I1(\mem[6][28] ),
    .S(_1370_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4763_ (.I0(\mem[5][28] ),
    .I1(\mem[7][28] ),
    .S(_1538_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4764_ (.I0(\mem[12][28] ),
    .I1(\mem[14][28] ),
    .S(_1351_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4765_ (.I0(\mem[13][28] ),
    .I1(\mem[15][28] ),
    .S(_1389_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4766_ (.I0(_1623_),
    .I1(_1624_),
    .I2(_1625_),
    .I3(_1626_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4767_ (.I0(\mem[1][28] ),
    .I1(\mem[3][28] ),
    .S(_1543_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4768_ (.I0(\mem[0][28] ),
    .I1(\mem[2][28] ),
    .S(_1601_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4769_ (.I0(\mem[9][28] ),
    .I1(\mem[11][28] ),
    .S(_1616_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4770_ (.I0(\mem[8][28] ),
    .I1(\mem[10][28] ),
    .S(_1495_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4771_ (.I0(_1628_),
    .I1(_1629_),
    .I2(_1630_),
    .I3(_1631_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4772_ (.I0(_1627_),
    .I1(_1632_),
    .S(_1620_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4773_ (.I0(net99),
    .I1(_1633_),
    .S(_1622_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4774_ (.I0(\mem[4][29] ),
    .I1(\mem[6][29] ),
    .S(_1370_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4775_ (.I0(\mem[5][29] ),
    .I1(\mem[7][29] ),
    .S(_1538_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4776_ (.I0(\mem[12][29] ),
    .I1(\mem[14][29] ),
    .S(_1351_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4777_ (.I0(\mem[13][29] ),
    .I1(\mem[15][29] ),
    .S(_1389_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4778_ (.I0(_1634_),
    .I1(_1635_),
    .I2(_1636_),
    .I3(_1637_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4779_ (.I0(\mem[1][29] ),
    .I1(\mem[3][29] ),
    .S(_1543_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4780_ (.I0(\mem[0][29] ),
    .I1(\mem[2][29] ),
    .S(_1601_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4781_ (.I0(\mem[9][29] ),
    .I1(\mem[11][29] ),
    .S(_1616_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4782_ (.I0(\mem[8][29] ),
    .I1(\mem[10][29] ),
    .S(_1495_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4783_ (.I0(_1639_),
    .I1(_1640_),
    .I2(_1641_),
    .I3(_1642_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4784_ (.I0(_1638_),
    .I1(_1643_),
    .S(_1620_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4785_ (.I0(net100),
    .I1(_1644_),
    .S(_1622_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4786_ (.I0(\mem[4][2] ),
    .I1(\mem[6][2] ),
    .S(_1370_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4787_ (.I0(\mem[5][2] ),
    .I1(\mem[7][2] ),
    .S(_1538_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4788_ (.I0(\mem[12][2] ),
    .I1(\mem[14][2] ),
    .S(_1351_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4789_ (.I0(\mem[13][2] ),
    .I1(\mem[15][2] ),
    .S(_1389_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4790_ (.I0(_1645_),
    .I1(_1646_),
    .I2(_1647_),
    .I3(_1648_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4791_ (.I0(\mem[1][2] ),
    .I1(\mem[3][2] ),
    .S(_1543_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4792_ (.I0(\mem[0][2] ),
    .I1(\mem[2][2] ),
    .S(_1601_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4793_ (.I0(\mem[9][2] ),
    .I1(\mem[11][2] ),
    .S(_1616_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4794_ (.I0(\mem[8][2] ),
    .I1(\mem[10][2] ),
    .S(_1355_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4795_ (.I0(_1650_),
    .I1(_1651_),
    .I2(_1652_),
    .I3(_1653_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4796_ (.I0(_1649_),
    .I1(_1654_),
    .S(_1620_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4797_ (.I0(net101),
    .I1(_1655_),
    .S(_1622_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4798_ (.I0(\mem[4][30] ),
    .I1(\mem[6][30] ),
    .S(_1370_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4799_ (.I0(\mem[5][30] ),
    .I1(\mem[7][30] ),
    .S(_1538_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4800_ (.I0(\mem[12][30] ),
    .I1(\mem[14][30] ),
    .S(_1351_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4801_ (.I0(\mem[13][30] ),
    .I1(\mem[15][30] ),
    .S(_1389_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4802_ (.I0(_1656_),
    .I1(_1657_),
    .I2(_1658_),
    .I3(_1659_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4803_ (.I0(\mem[1][30] ),
    .I1(\mem[3][30] ),
    .S(_1543_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4804_ (.I0(\mem[0][30] ),
    .I1(\mem[2][30] ),
    .S(_1601_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4805_ (.I0(\mem[9][30] ),
    .I1(\mem[11][30] ),
    .S(_1616_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4806_ (.I0(\mem[8][30] ),
    .I1(\mem[10][30] ),
    .S(_1355_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4807_ (.I0(_1661_),
    .I1(_1662_),
    .I2(_1663_),
    .I3(_1664_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4808_ (.I0(_1660_),
    .I1(_1665_),
    .S(_1620_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4809_ (.I0(net102),
    .I1(_1666_),
    .S(_1622_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4810_ (.I0(\mem[4][31] ),
    .I1(\mem[6][31] ),
    .S(_1370_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4811_ (.I0(\mem[5][31] ),
    .I1(\mem[7][31] ),
    .S(_1538_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4812_ (.I0(\mem[12][31] ),
    .I1(\mem[14][31] ),
    .S(_1351_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4813_ (.I0(\mem[13][31] ),
    .I1(\mem[15][31] ),
    .S(_1389_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4814_ (.I0(_1667_),
    .I1(_1668_),
    .I2(_1669_),
    .I3(_1670_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4815_ (.I0(\mem[1][31] ),
    .I1(\mem[3][31] ),
    .S(_1543_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4816_ (.I0(\mem[0][31] ),
    .I1(\mem[2][31] ),
    .S(_1601_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4817_ (.I0(\mem[9][31] ),
    .I1(\mem[11][31] ),
    .S(_1616_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4818_ (.I0(\mem[8][31] ),
    .I1(\mem[10][31] ),
    .S(_1355_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4819_ (.I0(_1672_),
    .I1(_1673_),
    .I2(_1674_),
    .I3(_1675_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4820_ (.I0(_1671_),
    .I1(_1676_),
    .S(_1620_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4821_ (.I0(net103),
    .I1(_1677_),
    .S(_1622_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4822_ (.I0(\mem[4][3] ),
    .I1(\mem[6][3] ),
    .S(_1370_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4823_ (.I0(\mem[5][3] ),
    .I1(\mem[7][3] ),
    .S(_1386_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4824_ (.I0(\mem[12][3] ),
    .I1(\mem[14][3] ),
    .S(_1351_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4825_ (.I0(\mem[13][3] ),
    .I1(\mem[15][3] ),
    .S(_1389_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4826_ (.I0(_1678_),
    .I1(_1679_),
    .I2(_1680_),
    .I3(_1681_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4827_ (.I0(\mem[1][3] ),
    .I1(\mem[3][3] ),
    .S(_1382_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4828_ (.I0(\mem[0][3] ),
    .I1(\mem[2][3] ),
    .S(_1601_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4829_ (.I0(\mem[9][3] ),
    .I1(\mem[11][3] ),
    .S(_1616_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4830_ (.I0(\mem[8][3] ),
    .I1(\mem[10][3] ),
    .S(_1355_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4831_ (.I0(_1683_),
    .I1(_1684_),
    .I2(_1685_),
    .I3(_1686_),
    .S0(_1605_),
    .S1(_1592_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4832_ (.I0(_1682_),
    .I1(_1687_),
    .S(_1620_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4833_ (.I0(net112),
    .I1(_1688_),
    .S(_1622_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4834_ (.I0(\mem[5][4] ),
    .I1(\mem[7][4] ),
    .S(_1523_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4835_ (.I0(\mem[4][4] ),
    .I1(\mem[6][4] ),
    .S(_1525_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4836_ (.I0(\mem[13][4] ),
    .I1(\mem[15][4] ),
    .S(_1356_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4837_ (.I0(\mem[12][4] ),
    .I1(\mem[14][4] ),
    .S(_1356_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4838_ (.I0(_1689_),
    .I1(_1690_),
    .I2(_1691_),
    .I3(_1692_),
    .S0(_1396_),
    .S1(_1612_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4839_ (.I0(\mem[0][4] ),
    .I1(\mem[2][4] ),
    .S(_1367_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4840_ (.I0(\mem[1][4] ),
    .I1(\mem[3][4] ),
    .S(_1523_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4841_ (.I0(\mem[8][4] ),
    .I1(\mem[10][4] ),
    .S(_1353_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4842_ (.I0(\mem[9][4] ),
    .I1(\mem[11][4] ),
    .S(_1359_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4843_ (.I0(_1694_),
    .I1(_1695_),
    .I2(_1696_),
    .I3(_1697_),
    .S0(_1534_),
    .S1(_1592_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4844_ (.I0(_1693_),
    .I1(_1698_),
    .S(_1620_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4845_ (.I0(net123),
    .I1(_1699_),
    .S(_1622_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4846_ (.I0(\mem[4][5] ),
    .I1(\mem[6][5] ),
    .S(_1370_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4847_ (.I0(\mem[5][5] ),
    .I1(\mem[7][5] ),
    .S(_1386_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4848_ (.I0(\mem[12][5] ),
    .I1(\mem[14][5] ),
    .S(_1351_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4849_ (.I0(\mem[13][5] ),
    .I1(\mem[15][5] ),
    .S(_1389_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4850_ (.I0(_1700_),
    .I1(_1701_),
    .I2(_1702_),
    .I3(_1703_),
    .S0(_1372_),
    .S1(_1612_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4851_ (.I0(\mem[1][5] ),
    .I1(\mem[3][5] ),
    .S(_1382_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4852_ (.I0(\mem[0][5] ),
    .I1(\mem[2][5] ),
    .S(_1601_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4853_ (.I0(\mem[9][5] ),
    .I1(\mem[11][5] ),
    .S(_1616_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4854_ (.I0(\mem[8][5] ),
    .I1(\mem[10][5] ),
    .S(_1355_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4855_ (.I0(_1705_),
    .I1(_1706_),
    .I2(_1707_),
    .I3(_1708_),
    .S0(_1605_),
    .S1(_1363_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4856_ (.I0(_1704_),
    .I1(_1709_),
    .S(_1620_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4857_ (.I0(net134),
    .I1(_1710_),
    .S(_1622_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4858_ (.I0(\mem[5][6] ),
    .I1(\mem[7][6] ),
    .S(_1523_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4859_ (.I0(\mem[4][6] ),
    .I1(\mem[6][6] ),
    .S(_1525_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4860_ (.I0(\mem[13][6] ),
    .I1(\mem[15][6] ),
    .S(_1356_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4861_ (.I0(\mem[12][6] ),
    .I1(\mem[14][6] ),
    .S(_1356_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4862_ (.I0(_1711_),
    .I1(_1712_),
    .I2(_1713_),
    .I3(_1714_),
    .S0(_1396_),
    .S1(_1612_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4863_ (.I0(\mem[0][6] ),
    .I1(\mem[2][6] ),
    .S(_1367_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4864_ (.I0(\mem[1][6] ),
    .I1(\mem[3][6] ),
    .S(_1525_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4865_ (.I0(\mem[8][6] ),
    .I1(\mem[10][6] ),
    .S(_1353_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4866_ (.I0(\mem[9][6] ),
    .I1(\mem[11][6] ),
    .S(_1359_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4867_ (.I0(_1716_),
    .I1(_1717_),
    .I2(_1718_),
    .I3(_1719_),
    .S0(_1534_),
    .S1(_1363_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4868_ (.I0(_1715_),
    .I1(_1720_),
    .S(_1620_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4869_ (.I0(net139),
    .I1(_1721_),
    .S(_1622_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4870_ (.I0(\mem[4][7] ),
    .I1(\mem[6][7] ),
    .S(_1370_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4871_ (.I0(\mem[5][7] ),
    .I1(\mem[7][7] ),
    .S(_1386_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4872_ (.I0(\mem[12][7] ),
    .I1(\mem[14][7] ),
    .S(_1351_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4873_ (.I0(\mem[13][7] ),
    .I1(\mem[15][7] ),
    .S(_1389_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4874_ (.I0(_1722_),
    .I1(_1723_),
    .I2(_1724_),
    .I3(_1725_),
    .S0(_1372_),
    .S1(_1373_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4875_ (.I0(\mem[1][7] ),
    .I1(\mem[3][7] ),
    .S(_1382_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4876_ (.I0(\mem[0][7] ),
    .I1(\mem[2][7] ),
    .S(_1601_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4877_ (.I0(\mem[9][7] ),
    .I1(\mem[11][7] ),
    .S(_1616_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4878_ (.I0(\mem[8][7] ),
    .I1(\mem[10][7] ),
    .S(_1355_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4879_ (.I0(_1727_),
    .I1(_1728_),
    .I2(_1729_),
    .I3(_1730_),
    .S0(_1605_),
    .S1(_1363_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4880_ (.I(_1376_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4881_ (.I(_1732_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4882_ (.I0(_1726_),
    .I1(_1731_),
    .S(_1733_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4883_ (.I(_0602_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4884_ (.I(_1735_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4885_ (.I0(net140),
    .I1(_1734_),
    .S(_1736_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4886_ (.I0(\mem[5][8] ),
    .I1(\mem[7][8] ),
    .S(_1523_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4887_ (.I0(\mem[4][8] ),
    .I1(\mem[6][8] ),
    .S(_1525_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4888_ (.I0(\mem[13][8] ),
    .I1(\mem[15][8] ),
    .S(_1356_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4889_ (.I0(\mem[12][8] ),
    .I1(\mem[14][8] ),
    .S(_1356_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4890_ (.I0(_1737_),
    .I1(_1738_),
    .I2(_1739_),
    .I3(_1740_),
    .S0(_1396_),
    .S1(_1373_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4891_ (.I0(\mem[0][8] ),
    .I1(\mem[2][8] ),
    .S(_1367_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4892_ (.I0(\mem[1][8] ),
    .I1(\mem[3][8] ),
    .S(_1525_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4893_ (.I0(\mem[8][8] ),
    .I1(\mem[10][8] ),
    .S(_1353_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4894_ (.I0(\mem[9][8] ),
    .I1(\mem[11][8] ),
    .S(_1359_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4895_ (.I0(_1742_),
    .I1(_1743_),
    .I2(_1744_),
    .I3(_1745_),
    .S0(_1534_),
    .S1(_1363_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4896_ (.I0(_1741_),
    .I1(_1746_),
    .S(_1733_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4897_ (.I0(net141),
    .I1(_1747_),
    .S(_1736_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4898_ (.I0(\mem[4][9] ),
    .I1(\mem[6][9] ),
    .S(_1370_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4899_ (.I0(\mem[5][9] ),
    .I1(\mem[7][9] ),
    .S(_1386_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4900_ (.I0(\mem[12][9] ),
    .I1(\mem[14][9] ),
    .S(_1351_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4901_ (.I0(\mem[13][9] ),
    .I1(\mem[15][9] ),
    .S(_1389_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4902_ (.I0(_1748_),
    .I1(_1749_),
    .I2(_1750_),
    .I3(_1751_),
    .S0(_1372_),
    .S1(_1373_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4903_ (.I0(\mem[1][9] ),
    .I1(\mem[3][9] ),
    .S(_1382_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4904_ (.I0(\mem[0][9] ),
    .I1(\mem[2][9] ),
    .S(_1353_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4905_ (.I0(\mem[9][9] ),
    .I1(\mem[11][9] ),
    .S(_1616_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4906_ (.I0(\mem[8][9] ),
    .I1(\mem[10][9] ),
    .S(_1355_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4907_ (.I0(_1753_),
    .I1(_1754_),
    .I2(_1755_),
    .I3(_1756_),
    .S0(_1395_),
    .S1(_1363_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4908_ (.I0(_1752_),
    .I1(_1757_),
    .S(_1733_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4909_ (.I0(net142),
    .I1(_1758_),
    .S(_1736_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _4910_ (.A1(net104),
    .A2(_2731_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4911_ (.I(_1362_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4912_ (.I(_2712_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _4913_ (.A1(_0600_),
    .A2(_0593_),
    .B(net2),
    .C(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4914_ (.I(_1762_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _4915_ (.A1(_2686_),
    .A2(\mem[10][0] ),
    .A3(_1735_),
    .B1(_1763_),
    .B2(\mem[11][0] ),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _4916_ (.A1(net73),
    .A2(net72),
    .A3(net74),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _4917_ (.A1(net2),
    .A2(_2711_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _4918_ (.A1(_2751_),
    .A2(_1765_),
    .B(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _4919_ (.A1(_1376_),
    .A2(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4920_ (.I(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4921_ (.I(_1391_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4922_ (.I(_0602_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _4923_ (.I(_2712_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _4924_ (.A1(_0600_),
    .A2(_0593_),
    .B(net2),
    .C(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4925_ (.I(_1773_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _4926_ (.A1(_1770_),
    .A2(\mem[8][0] ),
    .A3(_1771_),
    .B1(_1774_),
    .B2(\mem[9][0] ),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _4927_ (.A1(_1760_),
    .A2(_1764_),
    .A3(_1769_),
    .A4(_1775_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4928_ (.A1(_1395_),
    .A2(\rd_ptr[2] ),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4929_ (.A1(_1395_),
    .A2(_1375_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4930_ (.I0(_1777_),
    .I1(_1778_),
    .S(_1767_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4931_ (.I(_1779_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4932_ (.I(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4933_ (.I(_2712_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4934_ (.I(_1782_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4935_ (.I0(\mem[13][0] ),
    .I1(\mem[15][0] ),
    .S(_1783_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4936_ (.I0(_1357_),
    .I1(_1784_),
    .S(_1735_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4937_ (.A1(_1361_),
    .A2(\rd_ptr[2] ),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4938_ (.A1(_1361_),
    .A2(_1376_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4939_ (.I0(_1786_),
    .I1(_1787_),
    .S(_1767_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4940_ (.I(_1788_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4941_ (.I(_1789_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4942_ (.I(_1761_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4943_ (.I0(\mem[12][0] ),
    .I1(\mem[14][0] ),
    .S(_1791_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4944_ (.I(_0603_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4945_ (.I0(_1360_),
    .I1(_1792_),
    .S(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _4946_ (.A1(_1781_),
    .A2(_1785_),
    .B1(_1790_),
    .B2(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _4947_ (.A1(net2),
    .A2(_1361_),
    .A3(\rd_ptr[2] ),
    .A4(_0612_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _4948_ (.A1(_2751_),
    .A2(_1765_),
    .B(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _4949_ (.A1(\rd_ptr[3] ),
    .A2(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4950_ (.A1(_0611_),
    .A2(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4951_ (.I(_1761_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4952_ (.I(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4953_ (.I0(\mem[8][0] ),
    .I1(\mem[10][0] ),
    .S(_1801_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _4954_ (.A1(\rd_ptr[2] ),
    .A2(_2711_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _4955_ (.I(net2),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _4956_ (.A1(_2751_),
    .A2(_1765_),
    .B(_1803_),
    .C(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4957_ (.I(_1805_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4958_ (.A1(_1802_),
    .A2(_1806_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4959_ (.I(_0601_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _4960_ (.A1(_1733_),
    .A2(_1808_),
    .A3(_1371_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4961_ (.I(_1534_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4962_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _4963_ (.A1(_1807_),
    .A2(_1809_),
    .B(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _4964_ (.A1(_1776_),
    .A2(_1795_),
    .A3(_1799_),
    .A4(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _4965_ (.A1(\rd_ptr[3] ),
    .A2(_1797_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _4966_ (.A1(_0611_),
    .A2(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4967_ (.I(_1782_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4968_ (.I0(\mem[4][0] ),
    .I1(\mem[6][0] ),
    .S(_1816_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4969_ (.A1(_1361_),
    .A2(_1803_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _4970_ (.A1(_0604_),
    .A2(_1817_),
    .A3(_1818_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4971_ (.I(_1786_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _4972_ (.A1(_2729_),
    .A2(_1354_),
    .A3(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4973_ (.I(_1761_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4974_ (.I(_1803_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4975_ (.I0(\mem[1][0] ),
    .I1(\mem[3][0] ),
    .I2(\mem[5][0] ),
    .I3(\mem[7][0] ),
    .S0(_1822_),
    .S1(_1823_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4976_ (.I0(_1352_),
    .I1(_1366_),
    .S(_1377_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _4977_ (.A1(\rd_ptr[2] ),
    .A2(_2711_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4978_ (.I(_1826_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4979_ (.I0(\mem[0][0] ),
    .I1(\mem[2][0] ),
    .S(_1782_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4980_ (.A1(_1827_),
    .A2(_1828_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4981_ (.A1(_1732_),
    .A2(_1368_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4982_ (.I(_0601_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _4983_ (.I0(_1824_),
    .I1(_1825_),
    .I2(_1829_),
    .I3(_1830_),
    .S0(_1831_),
    .S1(_1810_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _4984_ (.A1(_1815_),
    .A2(_1819_),
    .A3(_1821_),
    .A4(_1832_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _4985_ (.A1(_1759_),
    .A2(_1813_),
    .A3(_1833_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _4986_ (.A1(net115),
    .A2(_2731_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4987_ (.A1(_0611_),
    .A2(_1814_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4988_ (.I(_1835_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4989_ (.I(_1362_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4990_ (.I(_1768_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _4991_ (.A1(_1770_),
    .A2(\mem[0][10] ),
    .A3(_1771_),
    .B1(_1774_),
    .B2(\mem[1][10] ),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4992_ (.I(_0602_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _4993_ (.A1(_2686_),
    .A2(\mem[2][10] ),
    .A3(_1840_),
    .B1(_1763_),
    .B2(\mem[3][10] ),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _4994_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_1839_),
    .A4(_1841_),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4995_ (.I(_1789_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4996_ (.I0(\mem[4][10] ),
    .I1(\mem[6][10] ),
    .S(_1783_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4997_ (.I0(_1384_),
    .I1(_1844_),
    .S(_1735_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4998_ (.I0(\mem[5][10] ),
    .I1(\mem[7][10] ),
    .S(_1791_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4999_ (.I0(_1383_),
    .I1(_1846_),
    .S(_1793_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5000_ (.A1(_1843_),
    .A2(_1845_),
    .B1(_1847_),
    .B2(_1781_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5001_ (.I(_1806_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5002_ (.I0(\mem[0][10] ),
    .I1(\mem[2][10] ),
    .S(_1801_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5003_ (.A1(_1849_),
    .A2(_1850_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5004_ (.A1(_1733_),
    .A2(_1808_),
    .A3(_1390_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5005_ (.A1(_1851_),
    .A2(_1852_),
    .B(_1811_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5006_ (.A1(_1836_),
    .A2(_1842_),
    .A3(_1848_),
    .A4(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _5007_ (.A1(_0610_),
    .A2(_1798_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5008_ (.I(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5009_ (.I(_1818_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5010_ (.I0(\mem[12][10] ),
    .I1(\mem[14][10] ),
    .S(_1816_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5011_ (.A1(_0604_),
    .A2(_1857_),
    .A3(_1858_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5012_ (.A1(_2729_),
    .A2(_1387_),
    .A3(_1820_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5013_ (.I0(\mem[9][10] ),
    .I1(\mem[11][10] ),
    .I2(\mem[13][10] ),
    .I3(\mem[15][10] ),
    .S0(_1822_),
    .S1(_1823_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5014_ (.I0(_1385_),
    .I1(_1394_),
    .S(_1377_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5015_ (.I0(\mem[8][10] ),
    .I1(\mem[10][10] ),
    .S(_1782_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5016_ (.A1(_1827_),
    .A2(_1863_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5017_ (.A1(_1732_),
    .A2(_1393_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5018_ (.I0(_1861_),
    .I1(_1862_),
    .I2(_1864_),
    .I3(_1865_),
    .S0(_1831_),
    .S1(_1810_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5019_ (.A1(_1856_),
    .A2(_1859_),
    .A3(_1860_),
    .A4(_1866_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5020_ (.A1(_1834_),
    .A2(_1854_),
    .A3(_1867_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5021_ (.I(_0611_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5022_ (.A1(net116),
    .A2(_1868_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5023_ (.I(_0602_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5024_ (.A1(_1770_),
    .A2(\mem[0][11] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][11] ),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5025_ (.A1(_2686_),
    .A2(\mem[2][11] ),
    .A3(_1840_),
    .B1(_1763_),
    .B2(\mem[3][11] ),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5026_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_1871_),
    .A4(_1872_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5027_ (.I0(\mem[4][11] ),
    .I1(\mem[6][11] ),
    .S(_1783_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5028_ (.I0(_1401_),
    .I1(_1874_),
    .S(_1735_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5029_ (.I0(\mem[5][11] ),
    .I1(\mem[7][11] ),
    .S(_1791_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5030_ (.I0(_1399_),
    .I1(_1876_),
    .S(_1793_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5031_ (.A1(_1843_),
    .A2(_1875_),
    .B1(_1877_),
    .B2(_1781_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5032_ (.I(_1800_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5033_ (.I0(\mem[0][11] ),
    .I1(\mem[2][11] ),
    .S(_1879_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5034_ (.A1(_1849_),
    .A2(_1880_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5035_ (.A1(_1733_),
    .A2(_1808_),
    .A3(_1406_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5036_ (.A1(_1881_),
    .A2(_1882_),
    .B(_1811_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5037_ (.A1(_1836_),
    .A2(_1873_),
    .A3(_1878_),
    .A4(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5038_ (.I(_0603_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5039_ (.I0(\mem[12][11] ),
    .I1(\mem[14][11] ),
    .S(_1816_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5040_ (.A1(_1885_),
    .A2(_1857_),
    .A3(_1886_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5041_ (.A1(_2729_),
    .A2(_1403_),
    .A3(_1820_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5042_ (.I0(\mem[9][11] ),
    .I1(\mem[11][11] ),
    .I2(\mem[13][11] ),
    .I3(\mem[15][11] ),
    .S0(_1822_),
    .S1(_1823_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5043_ (.I0(_1402_),
    .I1(_1409_),
    .S(_1377_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5044_ (.I0(\mem[8][11] ),
    .I1(\mem[10][11] ),
    .S(_1782_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5045_ (.A1(_1827_),
    .A2(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5046_ (.A1(_1732_),
    .A2(_1408_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5047_ (.I0(_1889_),
    .I1(_1890_),
    .I2(_1892_),
    .I3(_1893_),
    .S0(_1831_),
    .S1(_1810_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5048_ (.A1(_1856_),
    .A2(_1887_),
    .A3(_1888_),
    .A4(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5049_ (.A1(_1869_),
    .A2(_1884_),
    .A3(_1895_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5050_ (.A1(net117),
    .A2(_1868_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5051_ (.A1(_1770_),
    .A2(\mem[0][12] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][12] ),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5052_ (.A1(_2686_),
    .A2(\mem[2][12] ),
    .A3(_1840_),
    .B1(_1763_),
    .B2(\mem[3][12] ),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5053_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_1897_),
    .A4(_1898_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5054_ (.I0(\mem[4][12] ),
    .I1(\mem[6][12] ),
    .S(_1783_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5055_ (.I0(_1413_),
    .I1(_1900_),
    .S(_1735_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5056_ (.I0(\mem[5][12] ),
    .I1(\mem[7][12] ),
    .S(_1791_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5057_ (.I0(_1412_),
    .I1(_1902_),
    .S(_1793_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5058_ (.A1(_1843_),
    .A2(_1901_),
    .B1(_1903_),
    .B2(_1781_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5059_ (.I0(\mem[0][12] ),
    .I1(\mem[2][12] ),
    .S(_1879_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5060_ (.A1(_1849_),
    .A2(_1905_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5061_ (.A1(_1733_),
    .A2(_1808_),
    .A3(_1417_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5062_ (.I(_1810_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5063_ (.A1(_1906_),
    .A2(_1907_),
    .B(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5064_ (.A1(_1836_),
    .A2(_1899_),
    .A3(_1904_),
    .A4(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5065_ (.I0(\mem[12][12] ),
    .I1(\mem[14][12] ),
    .S(_1816_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5066_ (.A1(_1885_),
    .A2(_1857_),
    .A3(_1911_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5067_ (.I(_0601_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5068_ (.I(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5069_ (.A1(_1914_),
    .A2(_1415_),
    .A3(_1820_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5070_ (.I0(\mem[9][12] ),
    .I1(\mem[11][12] ),
    .I2(\mem[13][12] ),
    .I3(\mem[15][12] ),
    .S0(_1822_),
    .S1(_1823_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5071_ (.I0(_1414_),
    .I1(_1420_),
    .S(_1377_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5072_ (.I0(\mem[8][12] ),
    .I1(\mem[10][12] ),
    .S(_1782_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5073_ (.A1(_1827_),
    .A2(_1918_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5074_ (.A1(_1732_),
    .A2(_1419_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5075_ (.I0(_1916_),
    .I1(_1917_),
    .I2(_1919_),
    .I3(_1920_),
    .S0(_1831_),
    .S1(_1810_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5076_ (.A1(_1856_),
    .A2(_1912_),
    .A3(_1915_),
    .A4(_1921_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5077_ (.A1(_1896_),
    .A2(_1910_),
    .A3(_1922_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5078_ (.A1(net118),
    .A2(_1868_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5079_ (.A1(_1770_),
    .A2(\mem[0][13] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][13] ),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5080_ (.A1(_2686_),
    .A2(\mem[2][13] ),
    .A3(_1840_),
    .B1(_1763_),
    .B2(\mem[3][13] ),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5081_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_1924_),
    .A4(_1925_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5082_ (.I(_1782_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5083_ (.I0(\mem[4][13] ),
    .I1(\mem[6][13] ),
    .S(_1927_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5084_ (.I(_0603_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5085_ (.I0(_1424_),
    .I1(_1928_),
    .S(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5086_ (.I0(\mem[5][13] ),
    .I1(\mem[7][13] ),
    .S(_1791_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5087_ (.I0(_1423_),
    .I1(_1931_),
    .S(_1793_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5088_ (.A1(_1843_),
    .A2(_1930_),
    .B1(_1932_),
    .B2(_1781_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5089_ (.I0(\mem[0][13] ),
    .I1(\mem[2][13] ),
    .S(_1879_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5090_ (.A1(_1849_),
    .A2(_1934_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5091_ (.A1(_1733_),
    .A2(_1808_),
    .A3(_1428_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5092_ (.A1(_1935_),
    .A2(_1936_),
    .B(_1908_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5093_ (.A1(_1836_),
    .A2(_1926_),
    .A3(_1933_),
    .A4(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5094_ (.I0(\mem[12][13] ),
    .I1(\mem[14][13] ),
    .S(_1816_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5095_ (.A1(_1885_),
    .A2(_1857_),
    .A3(_1939_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5096_ (.I(_1786_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5097_ (.A1(_1914_),
    .A2(_1426_),
    .A3(_1941_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5098_ (.I(_1803_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5099_ (.I0(\mem[9][13] ),
    .I1(\mem[11][13] ),
    .I2(\mem[13][13] ),
    .I3(\mem[15][13] ),
    .S0(_1822_),
    .S1(_1943_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5100_ (.I(_1376_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5101_ (.I0(_1425_),
    .I1(_1431_),
    .S(_1945_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5102_ (.I(_2712_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5103_ (.I0(\mem[8][13] ),
    .I1(\mem[10][13] ),
    .S(_1947_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5104_ (.A1(_1827_),
    .A2(_1948_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5105_ (.A1(_1732_),
    .A2(_1430_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5106_ (.I0(_1944_),
    .I1(_1946_),
    .I2(_1949_),
    .I3(_1950_),
    .S0(_1831_),
    .S1(_1810_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5107_ (.A1(_1856_),
    .A2(_1940_),
    .A3(_1942_),
    .A4(_1951_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5108_ (.A1(_1923_),
    .A2(_1938_),
    .A3(_1952_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5109_ (.A1(net119),
    .A2(_1868_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5110_ (.A1(_1770_),
    .A2(\mem[0][14] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][14] ),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5111_ (.A1(_2686_),
    .A2(\mem[2][14] ),
    .A3(_1840_),
    .B1(_1763_),
    .B2(\mem[3][14] ),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5112_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_1954_),
    .A4(_1955_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5113_ (.I0(\mem[4][14] ),
    .I1(\mem[6][14] ),
    .S(_1927_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5114_ (.I0(_1435_),
    .I1(_1957_),
    .S(_1929_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5115_ (.I0(\mem[5][14] ),
    .I1(\mem[7][14] ),
    .S(_1791_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5116_ (.I0(_1434_),
    .I1(_1959_),
    .S(_1793_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5117_ (.A1(_1843_),
    .A2(_1958_),
    .B1(_1960_),
    .B2(_1781_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5118_ (.I(_1806_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5119_ (.I0(\mem[0][14] ),
    .I1(\mem[2][14] ),
    .S(_1879_),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5120_ (.A1(_1962_),
    .A2(_1963_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5121_ (.A1(_1733_),
    .A2(_1808_),
    .A3(_1439_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5122_ (.A1(_1964_),
    .A2(_1965_),
    .B(_1908_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5123_ (.A1(_1836_),
    .A2(_1956_),
    .A3(_1961_),
    .A4(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5124_ (.I(_1818_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5125_ (.I0(\mem[12][14] ),
    .I1(\mem[14][14] ),
    .S(_1816_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5126_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_1969_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5127_ (.A1(_1914_),
    .A2(_1437_),
    .A3(_1941_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5128_ (.I0(\mem[9][14] ),
    .I1(\mem[11][14] ),
    .I2(\mem[13][14] ),
    .I3(\mem[15][14] ),
    .S0(_1822_),
    .S1(_1943_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5129_ (.I0(_1436_),
    .I1(_1443_),
    .S(_1945_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5130_ (.I0(\mem[8][14] ),
    .I1(\mem[10][14] ),
    .S(_1947_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5131_ (.A1(_1827_),
    .A2(_1974_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5132_ (.A1(_1732_),
    .A2(_1442_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5133_ (.I0(_1972_),
    .I1(_1973_),
    .I2(_1975_),
    .I3(_1976_),
    .S0(_1831_),
    .S1(_1810_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5134_ (.A1(_1856_),
    .A2(_1970_),
    .A3(_1971_),
    .A4(_1977_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5135_ (.A1(_1953_),
    .A2(_1967_),
    .A3(_1978_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5136_ (.A1(net120),
    .A2(_1868_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5137_ (.A1(_1770_),
    .A2(\mem[0][15] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][15] ),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5138_ (.A1(_2686_),
    .A2(\mem[2][15] ),
    .A3(_1840_),
    .B1(_1763_),
    .B2(\mem[3][15] ),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5139_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_1980_),
    .A4(_1981_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5140_ (.I0(\mem[4][15] ),
    .I1(\mem[6][15] ),
    .S(_1927_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5141_ (.I0(_1448_),
    .I1(_1983_),
    .S(_1929_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5142_ (.I0(\mem[5][15] ),
    .I1(\mem[7][15] ),
    .S(_1791_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5143_ (.I0(_1447_),
    .I1(_1985_),
    .S(_1793_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5144_ (.A1(_1843_),
    .A2(_1984_),
    .B1(_1986_),
    .B2(_1781_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5145_ (.I0(\mem[0][15] ),
    .I1(\mem[2][15] ),
    .S(_1879_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5146_ (.A1(_1962_),
    .A2(_1988_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5147_ (.I(_1732_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5148_ (.A1(_1990_),
    .A2(_1808_),
    .A3(_1452_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5149_ (.A1(_1989_),
    .A2(_1991_),
    .B(_1908_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5150_ (.A1(_1836_),
    .A2(_1982_),
    .A3(_1987_),
    .A4(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5151_ (.I(_1782_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5152_ (.I0(\mem[12][15] ),
    .I1(\mem[14][15] ),
    .S(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5153_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_1995_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5154_ (.A1(_1914_),
    .A2(_1450_),
    .A3(_1941_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5155_ (.I0(\mem[9][15] ),
    .I1(\mem[11][15] ),
    .I2(\mem[13][15] ),
    .I3(\mem[15][15] ),
    .S0(_1822_),
    .S1(_1943_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5156_ (.I0(_1449_),
    .I1(_1456_),
    .S(_1945_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5157_ (.I0(\mem[8][15] ),
    .I1(\mem[10][15] ),
    .S(_1947_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5158_ (.A1(_1827_),
    .A2(_2000_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5159_ (.A1(_1732_),
    .A2(_1455_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5160_ (.I(_1534_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5161_ (.I0(_1998_),
    .I1(_1999_),
    .I2(_2001_),
    .I3(_2002_),
    .S0(_1831_),
    .S1(_2003_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5162_ (.A1(_1856_),
    .A2(_1996_),
    .A3(_1997_),
    .A4(_2004_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5163_ (.A1(_1979_),
    .A2(_1993_),
    .A3(_2005_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5164_ (.A1(net121),
    .A2(_1868_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5165_ (.A1(_1770_),
    .A2(\mem[0][16] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][16] ),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5166_ (.I(_0602_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5167_ (.A1(_2686_),
    .A2(\mem[2][16] ),
    .A3(_2008_),
    .B1(_1763_),
    .B2(\mem[3][16] ),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5168_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_2007_),
    .A4(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5169_ (.I0(\mem[4][16] ),
    .I1(\mem[6][16] ),
    .S(_1927_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5170_ (.I0(_1461_),
    .I1(_2011_),
    .S(_1929_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5171_ (.I(_1761_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5172_ (.I0(\mem[5][16] ),
    .I1(\mem[7][16] ),
    .S(_2013_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5173_ (.I0(_1460_),
    .I1(_2014_),
    .S(_1793_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5174_ (.A1(_1843_),
    .A2(_2012_),
    .B1(_2015_),
    .B2(_1781_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5175_ (.I0(\mem[0][16] ),
    .I1(\mem[2][16] ),
    .S(_1879_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5176_ (.A1(_1962_),
    .A2(_2017_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5177_ (.I(_0601_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5178_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1468_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5179_ (.A1(_2018_),
    .A2(_2020_),
    .B(_1908_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5180_ (.A1(_1836_),
    .A2(_2010_),
    .A3(_2016_),
    .A4(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5181_ (.I0(\mem[12][16] ),
    .I1(\mem[14][16] ),
    .S(_1994_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5182_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_2023_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5183_ (.A1(_1914_),
    .A2(_1465_),
    .A3(_1941_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5184_ (.I0(\mem[9][16] ),
    .I1(\mem[11][16] ),
    .I2(\mem[13][16] ),
    .I3(\mem[15][16] ),
    .S0(_1822_),
    .S1(_1943_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5185_ (.I0(_1463_),
    .I1(_1471_),
    .S(_1945_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5186_ (.I0(\mem[8][16] ),
    .I1(\mem[10][16] ),
    .S(_1947_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5187_ (.A1(_1827_),
    .A2(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5188_ (.I(_1376_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5189_ (.A1(_2030_),
    .A2(_1470_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5190_ (.I0(_2026_),
    .I1(_2027_),
    .I2(_2029_),
    .I3(_2031_),
    .S0(_1831_),
    .S1(_2003_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5191_ (.A1(_1856_),
    .A2(_2024_),
    .A3(_2025_),
    .A4(_2032_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5192_ (.A1(_2006_),
    .A2(_2022_),
    .A3(_2033_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5193_ (.A1(net122),
    .A2(_1868_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5194_ (.A1(_1770_),
    .A2(\mem[0][17] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][17] ),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5195_ (.A1(_2686_),
    .A2(\mem[2][17] ),
    .A3(_2008_),
    .B1(_1763_),
    .B2(\mem[3][17] ),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5196_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_2035_),
    .A4(_2036_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5197_ (.I0(\mem[4][17] ),
    .I1(\mem[6][17] ),
    .S(_1927_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5198_ (.I0(_1476_),
    .I1(_2038_),
    .S(_1929_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5199_ (.I0(\mem[5][17] ),
    .I1(\mem[7][17] ),
    .S(_2013_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5200_ (.I(_0603_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5201_ (.I0(_1475_),
    .I1(_2040_),
    .S(_2041_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5202_ (.A1(_1843_),
    .A2(_2039_),
    .B1(_2042_),
    .B2(_1781_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5203_ (.I0(\mem[0][17] ),
    .I1(\mem[2][17] ),
    .S(_1879_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5204_ (.A1(_1962_),
    .A2(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5205_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1480_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5206_ (.A1(_2045_),
    .A2(_2046_),
    .B(_1908_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5207_ (.A1(_1836_),
    .A2(_2037_),
    .A3(_2043_),
    .A4(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5208_ (.I0(\mem[12][17] ),
    .I1(\mem[14][17] ),
    .S(_1994_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5209_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_2049_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5210_ (.A1(_1914_),
    .A2(_1478_),
    .A3(_1941_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5211_ (.I0(\mem[9][17] ),
    .I1(\mem[11][17] ),
    .I2(\mem[13][17] ),
    .I3(\mem[15][17] ),
    .S0(_1822_),
    .S1(_1943_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5212_ (.I0(_1477_),
    .I1(_1483_),
    .S(_1945_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5213_ (.I0(\mem[8][17] ),
    .I1(\mem[10][17] ),
    .S(_1947_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5214_ (.A1(_1827_),
    .A2(_2054_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5215_ (.A1(_2030_),
    .A2(_1482_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5216_ (.I(_0601_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5217_ (.I0(_2052_),
    .I1(_2053_),
    .I2(_2055_),
    .I3(_2056_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5218_ (.A1(_1856_),
    .A2(_2050_),
    .A3(_2051_),
    .A4(_2058_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5219_ (.A1(_2034_),
    .A2(_2048_),
    .A3(_2059_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5220_ (.A1(net124),
    .A2(_1868_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5221_ (.I(_1391_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5222_ (.A1(_2061_),
    .A2(\mem[0][18] ),
    .A3(_1870_),
    .B1(_1774_),
    .B2(\mem[1][18] ),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5223_ (.I(_0614_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5224_ (.A1(_2063_),
    .A2(\mem[2][18] ),
    .A3(_2008_),
    .B1(_1763_),
    .B2(\mem[3][18] ),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5225_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_2062_),
    .A4(_2064_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5226_ (.I0(\mem[4][18] ),
    .I1(\mem[6][18] ),
    .S(_1927_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5227_ (.I0(_1487_),
    .I1(_2066_),
    .S(_1929_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5228_ (.I0(\mem[5][18] ),
    .I1(\mem[7][18] ),
    .S(_2013_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5229_ (.I0(_1486_),
    .I1(_2068_),
    .S(_2041_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5230_ (.A1(_1843_),
    .A2(_2067_),
    .B1(_2069_),
    .B2(_1781_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5231_ (.I0(\mem[0][18] ),
    .I1(\mem[2][18] ),
    .S(_1879_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5232_ (.A1(_1962_),
    .A2(_2071_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5233_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1492_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5234_ (.A1(_2072_),
    .A2(_2073_),
    .B(_1908_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5235_ (.A1(_1836_),
    .A2(_2065_),
    .A3(_2070_),
    .A4(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5236_ (.I0(\mem[12][18] ),
    .I1(\mem[14][18] ),
    .S(_1994_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5237_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_2076_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5238_ (.A1(_1914_),
    .A2(_1489_),
    .A3(_1941_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5239_ (.I(_1761_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5240_ (.I0(\mem[9][18] ),
    .I1(\mem[11][18] ),
    .I2(\mem[13][18] ),
    .I3(\mem[15][18] ),
    .S0(_2079_),
    .S1(_1943_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5241_ (.I0(_1488_),
    .I1(_1496_),
    .S(_1945_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5242_ (.I0(\mem[8][18] ),
    .I1(\mem[10][18] ),
    .S(_1947_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5243_ (.A1(_1827_),
    .A2(_2082_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5244_ (.A1(_2030_),
    .A2(_1494_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5245_ (.I0(_2080_),
    .I1(_2081_),
    .I2(_2083_),
    .I3(_2084_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5246_ (.A1(_1856_),
    .A2(_2077_),
    .A3(_2078_),
    .A4(_2085_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5247_ (.A1(_2060_),
    .A2(_2075_),
    .A3(_2086_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5248_ (.A1(net125),
    .A2(_1868_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5249_ (.I(_1773_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5250_ (.A1(_2061_),
    .A2(\mem[0][19] ),
    .A3(_1870_),
    .B1(_2088_),
    .B2(\mem[1][19] ),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5251_ (.I(_1762_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5252_ (.A1(_2063_),
    .A2(\mem[2][19] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][19] ),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5253_ (.A1(_1837_),
    .A2(_1838_),
    .A3(_2089_),
    .A4(_2091_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5254_ (.I0(\mem[4][19] ),
    .I1(\mem[6][19] ),
    .S(_1927_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5255_ (.I0(_1502_),
    .I1(_2093_),
    .S(_1929_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5256_ (.I0(\mem[5][19] ),
    .I1(\mem[7][19] ),
    .S(_2013_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5257_ (.I0(_1501_),
    .I1(_2095_),
    .S(_2041_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5258_ (.I(_1780_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5259_ (.A1(_1843_),
    .A2(_2094_),
    .B1(_2096_),
    .B2(_2097_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5260_ (.I0(\mem[0][19] ),
    .I1(\mem[2][19] ),
    .S(_1879_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5261_ (.A1(_1962_),
    .A2(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5262_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1506_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5263_ (.A1(_2100_),
    .A2(_2101_),
    .B(_1908_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5264_ (.A1(_1836_),
    .A2(_2092_),
    .A3(_2098_),
    .A4(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5265_ (.I0(\mem[12][19] ),
    .I1(\mem[14][19] ),
    .S(_1994_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5266_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5267_ (.A1(_1914_),
    .A2(_1504_),
    .A3(_1941_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5268_ (.I0(\mem[9][19] ),
    .I1(\mem[11][19] ),
    .I2(\mem[13][19] ),
    .I3(\mem[15][19] ),
    .S0(_2079_),
    .S1(_1943_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5269_ (.I0(_1503_),
    .I1(_1509_),
    .S(_1945_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5270_ (.I(_1826_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5271_ (.I0(\mem[8][19] ),
    .I1(\mem[10][19] ),
    .S(_1947_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5272_ (.A1(_2109_),
    .A2(_2110_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5273_ (.A1(_2030_),
    .A2(_1508_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5274_ (.I0(_2107_),
    .I1(_2108_),
    .I2(_2111_),
    .I3(_2112_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5275_ (.A1(_1856_),
    .A2(_2105_),
    .A3(_2106_),
    .A4(_2113_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5276_ (.A1(_2087_),
    .A2(_2103_),
    .A3(_2114_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5277_ (.A1(net105),
    .A2(_1868_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5278_ (.I(_1835_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5279_ (.I(_1362_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5280_ (.I(_1768_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5281_ (.A1(_2061_),
    .A2(\mem[0][1] ),
    .A3(_1870_),
    .B1(_2088_),
    .B2(\mem[1][1] ),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5282_ (.A1(_2063_),
    .A2(\mem[2][1] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][1] ),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5283_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2119_),
    .A4(_2120_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5284_ (.I(_1789_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5285_ (.I0(\mem[4][1] ),
    .I1(\mem[6][1] ),
    .S(_1927_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5286_ (.I0(_1513_),
    .I1(_2123_),
    .S(_1929_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5287_ (.I0(\mem[5][1] ),
    .I1(\mem[7][1] ),
    .S(_2013_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5288_ (.I0(_1512_),
    .I1(_2125_),
    .S(_2041_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5289_ (.A1(_2122_),
    .A2(_2124_),
    .B1(_2126_),
    .B2(_2097_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5290_ (.I0(\mem[0][1] ),
    .I1(\mem[2][1] ),
    .S(_1879_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5291_ (.A1(_1962_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5292_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1517_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5293_ (.A1(_2129_),
    .A2(_2130_),
    .B(_1908_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5294_ (.A1(_2116_),
    .A2(_2121_),
    .A3(_2127_),
    .A4(_2131_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5295_ (.I(_1855_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5296_ (.I0(\mem[12][1] ),
    .I1(\mem[14][1] ),
    .S(_1994_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5297_ (.A1(_1885_),
    .A2(_1968_),
    .A3(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5298_ (.A1(_1914_),
    .A2(_1515_),
    .A3(_1941_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5299_ (.I0(\mem[9][1] ),
    .I1(\mem[11][1] ),
    .I2(\mem[13][1] ),
    .I3(\mem[15][1] ),
    .S0(_2079_),
    .S1(_1943_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5300_ (.I0(_1514_),
    .I1(_1520_),
    .S(_1945_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5301_ (.I0(\mem[8][1] ),
    .I1(\mem[10][1] ),
    .S(_1947_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5302_ (.A1(_2109_),
    .A2(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5303_ (.A1(_2030_),
    .A2(_1519_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5304_ (.I0(_2137_),
    .I1(_2138_),
    .I2(_2140_),
    .I3(_2141_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5305_ (.A1(_2133_),
    .A2(_2135_),
    .A3(_2136_),
    .A4(_2142_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5306_ (.A1(_2115_),
    .A2(_2132_),
    .A3(_2143_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5307_ (.I(_1835_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5308_ (.I(_1791_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5309_ (.I0(\mem[4][20] ),
    .I1(\mem[6][20] ),
    .S(_2145_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5310_ (.A1(_1736_),
    .A2(_1857_),
    .A3(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5311_ (.A1(_2729_),
    .A2(_1524_),
    .A3(_1820_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5312_ (.A1(_2144_),
    .A2(_2147_),
    .A3(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5313_ (.I0(\mem[1][20] ),
    .I1(\mem[3][20] ),
    .I2(\mem[5][20] ),
    .I3(\mem[7][20] ),
    .S0(_1801_),
    .S1(_1823_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5314_ (.I(_0601_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5315_ (.I(_1376_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5316_ (.I0(_1526_),
    .I1(_1530_),
    .S(_2152_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5317_ (.A1(_2151_),
    .A2(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5318_ (.A1(_1736_),
    .A2(_2150_),
    .B(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5319_ (.A1(_1378_),
    .A2(_1831_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5320_ (.I0(\mem[0][20] ),
    .I1(\mem[2][20] ),
    .S(_2145_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5321_ (.A1(_1531_),
    .A2(_2156_),
    .B1(_2157_),
    .B2(_1849_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5322_ (.I0(_2155_),
    .I1(_2158_),
    .S(_1811_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5323_ (.A1(net126),
    .A2(_2731_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5324_ (.I(_1534_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5325_ (.I(_1391_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5326_ (.I(_0602_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5327_ (.I(_1773_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5328_ (.A1(_2162_),
    .A2(\mem[8][20] ),
    .A3(_2163_),
    .B1(_2164_),
    .B2(\mem[9][20] ),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5329_ (.I(_0614_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5330_ (.I(_1762_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5331_ (.A1(_2166_),
    .A2(\mem[10][20] ),
    .A3(_2163_),
    .B1(_2167_),
    .B2(\mem[11][20] ),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5332_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2165_),
    .A4(_2168_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5333_ (.I(_1761_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5334_ (.I0(\mem[12][20] ),
    .I1(\mem[14][20] ),
    .S(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5335_ (.I(_0602_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5336_ (.I0(_1527_),
    .I1(_2171_),
    .S(_2172_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5337_ (.I(_1761_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5338_ (.I0(\mem[13][20] ),
    .I1(\mem[15][20] ),
    .S(_2174_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5339_ (.I(_0602_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5340_ (.I0(_1528_),
    .I1(_2175_),
    .S(_2176_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5341_ (.I(_1780_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5342_ (.A1(_1790_),
    .A2(_2173_),
    .B1(_2177_),
    .B2(_2178_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5343_ (.I0(\mem[8][20] ),
    .I1(\mem[10][20] ),
    .S(_1783_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5344_ (.A1(_1806_),
    .A2(_2180_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5345_ (.I(_0601_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5346_ (.A1(_1378_),
    .A2(_2182_),
    .A3(_1533_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5347_ (.A1(_2181_),
    .A2(_2183_),
    .B(_1760_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _5348_ (.A1(_1799_),
    .A2(_2169_),
    .A3(_2179_),
    .A4(_2184_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _5349_ (.A1(_2149_),
    .A2(_2159_),
    .B(_2160_),
    .C(_2185_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5350_ (.I(_0611_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5351_ (.A1(net127),
    .A2(_2186_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5352_ (.I(_0602_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5353_ (.A1(_2061_),
    .A2(\mem[0][21] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][21] ),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5354_ (.A1(_2063_),
    .A2(\mem[2][21] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][21] ),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5355_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2189_),
    .A4(_2190_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5356_ (.I0(\mem[4][21] ),
    .I1(\mem[6][21] ),
    .S(_1927_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5357_ (.I0(_1539_),
    .I1(_2192_),
    .S(_1929_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5358_ (.I0(\mem[5][21] ),
    .I1(\mem[7][21] ),
    .S(_2013_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5359_ (.I0(_1537_),
    .I1(_2194_),
    .S(_2041_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5360_ (.A1(_2122_),
    .A2(_2193_),
    .B1(_2195_),
    .B2(_2097_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5361_ (.I(_1800_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5362_ (.I0(\mem[0][21] ),
    .I1(\mem[2][21] ),
    .S(_2197_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5363_ (.A1(_1962_),
    .A2(_2198_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5364_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1544_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5365_ (.A1(_2199_),
    .A2(_2200_),
    .B(_1908_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5366_ (.A1(_2116_),
    .A2(_2191_),
    .A3(_2196_),
    .A4(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5367_ (.I(_0603_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5368_ (.I0(\mem[12][21] ),
    .I1(\mem[14][21] ),
    .S(_1994_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5369_ (.A1(_2203_),
    .A2(_1968_),
    .A3(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5370_ (.A1(_1914_),
    .A2(_1541_),
    .A3(_1941_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5371_ (.I0(\mem[9][21] ),
    .I1(\mem[11][21] ),
    .I2(\mem[13][21] ),
    .I3(\mem[15][21] ),
    .S0(_2079_),
    .S1(_1943_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5372_ (.I0(_1540_),
    .I1(_1547_),
    .S(_1945_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5373_ (.I0(\mem[8][21] ),
    .I1(\mem[10][21] ),
    .S(_1947_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5374_ (.A1(_2109_),
    .A2(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5375_ (.A1(_2030_),
    .A2(_1546_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5376_ (.I0(_2207_),
    .I1(_2208_),
    .I2(_2210_),
    .I3(_2211_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5377_ (.A1(_2133_),
    .A2(_2205_),
    .A3(_2206_),
    .A4(_2212_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5378_ (.A1(_2187_),
    .A2(_2202_),
    .A3(_2213_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5379_ (.I0(\mem[4][22] ),
    .I1(\mem[6][22] ),
    .S(_2145_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5380_ (.A1(_1736_),
    .A2(_1857_),
    .A3(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5381_ (.A1(_2729_),
    .A2(_1550_),
    .A3(_1820_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5382_ (.A1(_2144_),
    .A2(_2215_),
    .A3(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5383_ (.I0(\mem[1][22] ),
    .I1(\mem[3][22] ),
    .I2(\mem[5][22] ),
    .I3(\mem[7][22] ),
    .S0(_1801_),
    .S1(_1823_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5384_ (.I0(_1551_),
    .I1(_1555_),
    .S(_1377_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5385_ (.A1(_2182_),
    .A2(_2219_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5386_ (.A1(_0604_),
    .A2(_2218_),
    .B(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5387_ (.I0(\mem[0][22] ),
    .I1(\mem[2][22] ),
    .S(_2145_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5388_ (.A1(_1556_),
    .A2(_2156_),
    .B1(_2222_),
    .B2(_1849_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5389_ (.I0(_2221_),
    .I1(_2223_),
    .S(_1811_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5390_ (.A1(net128),
    .A2(_2731_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5391_ (.A1(_2162_),
    .A2(\mem[8][22] ),
    .A3(_2163_),
    .B1(_2164_),
    .B2(\mem[9][22] ),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5392_ (.A1(_2166_),
    .A2(\mem[10][22] ),
    .A3(_2163_),
    .B1(_2167_),
    .B2(\mem[11][22] ),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5393_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2226_),
    .A4(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5394_ (.I0(\mem[12][22] ),
    .I1(\mem[14][22] ),
    .S(_2174_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5395_ (.I0(_1552_),
    .I1(_2229_),
    .S(_2176_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5396_ (.I0(\mem[13][22] ),
    .I1(\mem[15][22] ),
    .S(_2174_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5397_ (.I0(_1553_),
    .I1(_2231_),
    .S(_2176_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5398_ (.A1(_1790_),
    .A2(_2230_),
    .B1(_2232_),
    .B2(_2178_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5399_ (.I0(\mem[8][22] ),
    .I1(\mem[10][22] ),
    .S(_1783_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5400_ (.A1(_1806_),
    .A2(_2234_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5401_ (.A1(_1378_),
    .A2(_2182_),
    .A3(_1558_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5402_ (.A1(_2235_),
    .A2(_2236_),
    .B(_1760_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _5403_ (.A1(_1799_),
    .A2(_2228_),
    .A3(_2233_),
    .A4(_2237_),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _5404_ (.A1(_2217_),
    .A2(_2224_),
    .B(_2225_),
    .C(_2238_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5405_ (.A1(net129),
    .A2(_2186_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5406_ (.A1(_2061_),
    .A2(\mem[0][23] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][23] ),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5407_ (.A1(_2063_),
    .A2(\mem[2][23] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][23] ),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5408_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2240_),
    .A4(_2241_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5409_ (.I0(\mem[4][23] ),
    .I1(\mem[6][23] ),
    .S(_1927_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5410_ (.I0(_1562_),
    .I1(_2243_),
    .S(_1929_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5411_ (.I0(\mem[5][23] ),
    .I1(\mem[7][23] ),
    .S(_2013_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5412_ (.I0(_1561_),
    .I1(_2245_),
    .S(_2041_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5413_ (.A1(_2122_),
    .A2(_2244_),
    .B1(_2246_),
    .B2(_2097_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5414_ (.I0(\mem[0][23] ),
    .I1(\mem[2][23] ),
    .S(_2197_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5415_ (.A1(_1962_),
    .A2(_2248_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5416_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1566_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5417_ (.I(_1810_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5418_ (.A1(_2249_),
    .A2(_2250_),
    .B(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5419_ (.A1(_2116_),
    .A2(_2242_),
    .A3(_2247_),
    .A4(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5420_ (.I0(\mem[12][23] ),
    .I1(\mem[14][23] ),
    .S(_1994_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5421_ (.A1(_2203_),
    .A2(_1968_),
    .A3(_2254_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _5422_ (.I(_1913_),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5423_ (.A1(_2256_),
    .A2(_1564_),
    .A3(_1941_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5424_ (.I0(\mem[9][23] ),
    .I1(\mem[11][23] ),
    .I2(\mem[13][23] ),
    .I3(\mem[15][23] ),
    .S0(_2079_),
    .S1(_1943_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5425_ (.I0(_1563_),
    .I1(_1569_),
    .S(_1945_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5426_ (.I0(\mem[8][23] ),
    .I1(\mem[10][23] ),
    .S(_1947_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5427_ (.A1(_2109_),
    .A2(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5428_ (.A1(_2030_),
    .A2(_1568_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5429_ (.I0(_2258_),
    .I1(_2259_),
    .I2(_2261_),
    .I3(_2262_),
    .S0(_2057_),
    .S1(_2003_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5430_ (.A1(_2133_),
    .A2(_2255_),
    .A3(_2257_),
    .A4(_2263_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5431_ (.A1(_2239_),
    .A2(_2253_),
    .A3(_2264_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5432_ (.I0(\mem[4][24] ),
    .I1(\mem[6][24] ),
    .S(_2145_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5433_ (.A1(_1736_),
    .A2(_1857_),
    .A3(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5434_ (.A1(_2729_),
    .A2(_1572_),
    .A3(_1820_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5435_ (.A1(_2144_),
    .A2(_2266_),
    .A3(_2267_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5436_ (.I0(\mem[1][24] ),
    .I1(\mem[3][24] ),
    .I2(\mem[5][24] ),
    .I3(\mem[7][24] ),
    .S0(_1801_),
    .S1(_1823_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5437_ (.I0(_1573_),
    .I1(_1577_),
    .S(_1377_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5438_ (.A1(_2182_),
    .A2(_2270_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5439_ (.A1(_0604_),
    .A2(_2269_),
    .B(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5440_ (.I0(\mem[0][24] ),
    .I1(\mem[2][24] ),
    .S(_2145_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5441_ (.A1(_1578_),
    .A2(_2156_),
    .B1(_2273_),
    .B2(_1849_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5442_ (.I0(_2272_),
    .I1(_2274_),
    .S(_1811_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5443_ (.A1(net130),
    .A2(_2731_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5444_ (.A1(_2162_),
    .A2(\mem[8][24] ),
    .A3(_2163_),
    .B1(_2164_),
    .B2(\mem[9][24] ),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5445_ (.A1(_2166_),
    .A2(\mem[10][24] ),
    .A3(_2163_),
    .B1(_2167_),
    .B2(\mem[11][24] ),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5446_ (.A1(_2161_),
    .A2(_1769_),
    .A3(_2277_),
    .A4(_2278_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5447_ (.I0(\mem[12][24] ),
    .I1(\mem[14][24] ),
    .S(_2174_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5448_ (.I0(_1574_),
    .I1(_2280_),
    .S(_2176_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5449_ (.I0(\mem[13][24] ),
    .I1(\mem[15][24] ),
    .S(_2174_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5450_ (.I0(_1575_),
    .I1(_2282_),
    .S(_2176_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5451_ (.A1(_1790_),
    .A2(_2281_),
    .B1(_2283_),
    .B2(_2178_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5452_ (.I0(\mem[8][24] ),
    .I1(\mem[10][24] ),
    .S(_1783_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5453_ (.A1(_1806_),
    .A2(_2285_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5454_ (.A1(_1378_),
    .A2(_2182_),
    .A3(_1580_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5455_ (.A1(_2286_),
    .A2(_2287_),
    .B(_1760_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _5456_ (.A1(_1799_),
    .A2(_2279_),
    .A3(_2284_),
    .A4(_2288_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _5457_ (.A1(_2268_),
    .A2(_2275_),
    .B(_2276_),
    .C(_2289_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5458_ (.A1(net131),
    .A2(_2186_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5459_ (.A1(_2061_),
    .A2(\mem[0][25] ),
    .A3(_2188_),
    .B1(_2088_),
    .B2(\mem[1][25] ),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _5460_ (.A1(_2063_),
    .A2(\mem[2][25] ),
    .A3(_2008_),
    .B1(_2090_),
    .B2(\mem[3][25] ),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5461_ (.A1(_2117_),
    .A2(_2118_),
    .A3(_2291_),
    .A4(_2292_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5462_ (.I(_1782_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5463_ (.I0(\mem[4][25] ),
    .I1(\mem[6][25] ),
    .S(_2294_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5464_ (.I(_0603_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5465_ (.I0(_1584_),
    .I1(_2295_),
    .S(_2296_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5466_ (.I0(\mem[5][25] ),
    .I1(\mem[7][25] ),
    .S(_2013_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5467_ (.I0(_1583_),
    .I1(_2298_),
    .S(_2041_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5468_ (.A1(_2122_),
    .A2(_2297_),
    .B1(_2299_),
    .B2(_2097_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5469_ (.I0(\mem[0][25] ),
    .I1(\mem[2][25] ),
    .S(_2197_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _5470_ (.A1(_1962_),
    .A2(_2301_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _5471_ (.A1(_1990_),
    .A2(_2019_),
    .A3(_1588_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5472_ (.A1(_2302_),
    .A2(_2303_),
    .B(_2251_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _5473_ (.A(_2686_),
    .B(_2687_),
    .CI(_2688_),
    .CO(_2689_),
    .S(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _5474_ (.A(_2690_),
    .B(_2691_),
    .CI(_2692_),
    .CO(_2693_),
    .S(\next_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5475_ (.A(_2694_),
    .B(_2695_),
    .CO(_2696_),
    .S(_2697_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5476_ (.A(_2694_),
    .B(\wr_ptr[1] ),
    .CO(_2698_),
    .S(_2699_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5477_ (.A(\wr_ptr[0] ),
    .B(_2695_),
    .CO(_2700_),
    .S(_2701_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5478_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_2702_),
    .S(_2703_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5479_ (.A(_2704_),
    .B(_2705_),
    .CO(_2706_),
    .S(_2707_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5480_ (.A(_2708_),
    .B(_0001_),
    .CO(_2709_),
    .S(_2710_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _5481_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .CO(_2711_),
    .S(_2712_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5482_ (.A(_2713_),
    .B(_2714_),
    .CO(_2715_),
    .S(_2716_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5483_ (.A(_2713_),
    .B(_2714_),
    .CO(_2717_),
    .S(_2718_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5484_ (.A(_2719_),
    .B(_2720_),
    .CO(_0002_),
    .S(_2721_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5485_ (.A(_2722_),
    .B(_2723_),
    .CO(_2724_),
    .S(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5486_ (.A(\wr_ptr[0] ),
    .B(_2716_),
    .CO(_2722_),
    .S(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5487_ (.A(\rd_ptr[1] ),
    .B(_2725_),
    .CO(_2726_),
    .S(_2727_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5488_ (.A(_2728_),
    .B(_2729_),
    .CO(_0000_),
    .S(_2730_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5489_ (.A(_2731_),
    .B(_0001_),
    .CO(_2725_),
    .S(_2732_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5490_ (.A(\rd_ptr[0] ),
    .B(_2730_),
    .CO(_2733_),
    .S(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5491_ (.A(_2734_),
    .B(_2688_),
    .CO(_2735_),
    .S(_2692_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5492_ (.A(_2691_),
    .B(_2692_),
    .CO(_2736_),
    .S(_2737_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5493_ (.A(_2708_),
    .B(_2730_),
    .CO(_2738_),
    .S(_2739_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5494_ (.A(_2740_),
    .B(_2741_),
    .CO(_2742_),
    .S(_2743_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5495_ (.A(net74),
    .B(_2741_),
    .CO(_2744_),
    .S(_2745_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5496_ (.A(net74),
    .B(net75),
    .CO(_2746_),
    .S(_2747_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _5497_ (.A(_2740_),
    .B(_2748_),
    .CO(_2749_),
    .S(_2750_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _5498_ (.A(_2741_),
    .B(_2704_),
    .CO(_2751_),
    .S(_2752_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5499_ (.A(_2741_),
    .B(_2704_),
    .CO(_2753_),
    .S(_2754_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5500_ (.A(_2741_),
    .B(net76),
    .CO(_2755_),
    .S(_2756_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5501_ (.A(net75),
    .B(_2704_),
    .CO(_2757_),
    .S(_2758_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5502_ (.A(net75),
    .B(net76),
    .CO(_2759_),
    .S(_2760_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _5503_ (.A(_2761_),
    .B(_2716_),
    .CO(_2690_),
    .S(\next_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \fifo_count[0]$_DFF_PN0_  (.D(\next_count[0] ),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \fifo_count[1]$_DFF_PN0_  (.D(\next_count[1] ),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \fifo_count[2]$_DFF_PN0_  (.D(\next_count[2] ),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \fifo_count[3]$_DFF_PN0_  (.D(\next_count[3] ),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \fifo_count[4]$_DFF_PN0_  (.D(\next_count[4] ),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net76));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][0]$_DFFE_PP_  (.D(_0007_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][10]$_DFFE_PP_  (.D(_0008_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][11]$_DFFE_PP_  (.D(_0009_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][12]$_DFFE_PP_  (.D(_0010_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][13]$_DFFE_PP_  (.D(_0011_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][14]$_DFFE_PP_  (.D(_0012_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][15]$_DFFE_PP_  (.D(_0013_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][16]$_DFFE_PP_  (.D(_0014_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][17]$_DFFE_PP_  (.D(_0015_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][18]$_DFFE_PP_  (.D(_0016_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][19]$_DFFE_PP_  (.D(_0017_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][1]$_DFFE_PP_  (.D(_0018_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][20]$_DFFE_PP_  (.D(_0019_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][21]$_DFFE_PP_  (.D(_0020_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][22]$_DFFE_PP_  (.D(_0021_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][23]$_DFFE_PP_  (.D(_0022_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][24]$_DFFE_PP_  (.D(_0023_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][25]$_DFFE_PP_  (.D(_0024_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][26]$_DFFE_PP_  (.D(_0025_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][27]$_DFFE_PP_  (.D(_0026_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][28]$_DFFE_PP_  (.D(_0027_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][29]$_DFFE_PP_  (.D(_0028_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][2]$_DFFE_PP_  (.D(_0029_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][30]$_DFFE_PP_  (.D(_0030_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][31]$_DFFE_PP_  (.D(_0031_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][3]$_DFFE_PP_  (.D(_0032_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][4]$_DFFE_PP_  (.D(_0033_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][5]$_DFFE_PP_  (.D(_0034_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][6]$_DFFE_PP_  (.D(_0035_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][7]$_DFFE_PP_  (.D(_0036_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][8]$_DFFE_PP_  (.D(_0037_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][9]$_DFFE_PP_  (.D(_0038_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][0]$_DFFE_PP_  (.D(_0039_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[10][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][10]$_DFFE_PP_  (.D(_0040_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[10][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][11]$_DFFE_PP_  (.D(_0041_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[10][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][12]$_DFFE_PP_  (.D(_0042_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[10][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][13]$_DFFE_PP_  (.D(_0043_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[10][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][14]$_DFFE_PP_  (.D(_0044_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[10][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][15]$_DFFE_PP_  (.D(_0045_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[10][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][16]$_DFFE_PP_  (.D(_0046_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[10][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][17]$_DFFE_PP_  (.D(_0047_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[10][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][18]$_DFFE_PP_  (.D(_0048_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[10][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][19]$_DFFE_PP_  (.D(_0049_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[10][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][1]$_DFFE_PP_  (.D(_0050_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[10][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][20]$_DFFE_PP_  (.D(_0051_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[10][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][21]$_DFFE_PP_  (.D(_0052_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[10][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][22]$_DFFE_PP_  (.D(_0053_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[10][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][23]$_DFFE_PP_  (.D(_0054_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[10][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][24]$_DFFE_PP_  (.D(_0055_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[10][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][25]$_DFFE_PP_  (.D(_0056_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[10][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][26]$_DFFE_PP_  (.D(_0057_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[10][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][27]$_DFFE_PP_  (.D(_0058_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[10][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][28]$_DFFE_PP_  (.D(_0059_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[10][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][29]$_DFFE_PP_  (.D(_0060_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[10][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][2]$_DFFE_PP_  (.D(_0061_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[10][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][30]$_DFFE_PP_  (.D(_0062_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[10][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][31]$_DFFE_PP_  (.D(_0063_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[10][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][3]$_DFFE_PP_  (.D(_0064_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[10][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][4]$_DFFE_PP_  (.D(_0065_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[10][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][5]$_DFFE_PP_  (.D(_0066_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[10][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][6]$_DFFE_PP_  (.D(_0067_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[10][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][7]$_DFFE_PP_  (.D(_0068_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[10][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][8]$_DFFE_PP_  (.D(_0069_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[10][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][9]$_DFFE_PP_  (.D(_0070_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[10][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][0]$_DFFE_PP_  (.D(_0071_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[11][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][10]$_DFFE_PP_  (.D(_0072_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[11][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][11]$_DFFE_PP_  (.D(_0073_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[11][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][12]$_DFFE_PP_  (.D(_0074_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[11][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][13]$_DFFE_PP_  (.D(_0075_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[11][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][14]$_DFFE_PP_  (.D(_0076_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[11][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][15]$_DFFE_PP_  (.D(_0077_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[11][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][16]$_DFFE_PP_  (.D(_0078_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[11][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][17]$_DFFE_PP_  (.D(_0079_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[11][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][18]$_DFFE_PP_  (.D(_0080_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[11][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][19]$_DFFE_PP_  (.D(_0081_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[11][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][1]$_DFFE_PP_  (.D(_0082_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[11][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][20]$_DFFE_PP_  (.D(_0083_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[11][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][21]$_DFFE_PP_  (.D(_0084_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[11][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][22]$_DFFE_PP_  (.D(_0085_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[11][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][23]$_DFFE_PP_  (.D(_0086_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[11][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][24]$_DFFE_PP_  (.D(_0087_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[11][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][25]$_DFFE_PP_  (.D(_0088_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[11][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][26]$_DFFE_PP_  (.D(_0089_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[11][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][27]$_DFFE_PP_  (.D(_0090_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[11][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][28]$_DFFE_PP_  (.D(_0091_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[11][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][29]$_DFFE_PP_  (.D(_0092_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[11][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][2]$_DFFE_PP_  (.D(_0093_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[11][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][30]$_DFFE_PP_  (.D(_0094_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[11][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][31]$_DFFE_PP_  (.D(_0095_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[11][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][3]$_DFFE_PP_  (.D(_0096_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[11][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][4]$_DFFE_PP_  (.D(_0097_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[11][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][5]$_DFFE_PP_  (.D(_0098_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[11][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][6]$_DFFE_PP_  (.D(_0099_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[11][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][7]$_DFFE_PP_  (.D(_0100_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[11][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][8]$_DFFE_PP_  (.D(_0101_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[11][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][9]$_DFFE_PP_  (.D(_0102_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[11][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][0]$_DFFE_PP_  (.D(_0103_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[12][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][10]$_DFFE_PP_  (.D(_0104_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[12][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][11]$_DFFE_PP_  (.D(_0105_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[12][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][12]$_DFFE_PP_  (.D(_0106_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[12][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][13]$_DFFE_PP_  (.D(_0107_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[12][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][14]$_DFFE_PP_  (.D(_0108_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[12][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][15]$_DFFE_PP_  (.D(_0109_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[12][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][16]$_DFFE_PP_  (.D(_0110_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[12][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][17]$_DFFE_PP_  (.D(_0111_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[12][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][18]$_DFFE_PP_  (.D(_0112_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[12][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][19]$_DFFE_PP_  (.D(_0113_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[12][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][1]$_DFFE_PP_  (.D(_0114_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[12][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][20]$_DFFE_PP_  (.D(_0115_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[12][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][21]$_DFFE_PP_  (.D(_0116_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[12][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][22]$_DFFE_PP_  (.D(_0117_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[12][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][23]$_DFFE_PP_  (.D(_0118_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[12][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][24]$_DFFE_PP_  (.D(_0119_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[12][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][25]$_DFFE_PP_  (.D(_0120_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[12][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][26]$_DFFE_PP_  (.D(_0121_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[12][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][27]$_DFFE_PP_  (.D(_0122_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[12][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][28]$_DFFE_PP_  (.D(_0123_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[12][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][29]$_DFFE_PP_  (.D(_0124_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[12][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][2]$_DFFE_PP_  (.D(_0125_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[12][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][30]$_DFFE_PP_  (.D(_0126_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[12][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][31]$_DFFE_PP_  (.D(_0127_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[12][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][3]$_DFFE_PP_  (.D(_0128_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[12][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][4]$_DFFE_PP_  (.D(_0129_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[12][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][5]$_DFFE_PP_  (.D(_0130_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[12][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][6]$_DFFE_PP_  (.D(_0131_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[12][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][7]$_DFFE_PP_  (.D(_0132_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[12][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][8]$_DFFE_PP_  (.D(_0133_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[12][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][9]$_DFFE_PP_  (.D(_0134_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[12][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][0]$_DFFE_PP_  (.D(_0135_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[13][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][10]$_DFFE_PP_  (.D(_0136_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[13][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][11]$_DFFE_PP_  (.D(_0137_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[13][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][12]$_DFFE_PP_  (.D(_0138_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[13][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][13]$_DFFE_PP_  (.D(_0139_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[13][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][14]$_DFFE_PP_  (.D(_0140_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[13][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][15]$_DFFE_PP_  (.D(_0141_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[13][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][16]$_DFFE_PP_  (.D(_0142_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[13][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][17]$_DFFE_PP_  (.D(_0143_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[13][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][18]$_DFFE_PP_  (.D(_0144_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[13][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][19]$_DFFE_PP_  (.D(_0145_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[13][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][1]$_DFFE_PP_  (.D(_0146_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[13][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][20]$_DFFE_PP_  (.D(_0147_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[13][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][21]$_DFFE_PP_  (.D(_0148_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[13][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][22]$_DFFE_PP_  (.D(_0149_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[13][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][23]$_DFFE_PP_  (.D(_0150_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[13][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][24]$_DFFE_PP_  (.D(_0151_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[13][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][25]$_DFFE_PP_  (.D(_0152_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[13][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][26]$_DFFE_PP_  (.D(_0153_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[13][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][27]$_DFFE_PP_  (.D(_0154_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[13][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][28]$_DFFE_PP_  (.D(_0155_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[13][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][29]$_DFFE_PP_  (.D(_0156_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[13][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][2]$_DFFE_PP_  (.D(_0157_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[13][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][30]$_DFFE_PP_  (.D(_0158_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[13][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][31]$_DFFE_PP_  (.D(_0159_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[13][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][3]$_DFFE_PP_  (.D(_0160_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[13][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][4]$_DFFE_PP_  (.D(_0161_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[13][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][5]$_DFFE_PP_  (.D(_0162_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[13][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][6]$_DFFE_PP_  (.D(_0163_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[13][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][7]$_DFFE_PP_  (.D(_0164_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[13][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][8]$_DFFE_PP_  (.D(_0165_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[13][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][9]$_DFFE_PP_  (.D(_0166_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[13][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][0]$_DFFE_PP_  (.D(_0167_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[14][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][10]$_DFFE_PP_  (.D(_0168_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[14][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][11]$_DFFE_PP_  (.D(_0169_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[14][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][12]$_DFFE_PP_  (.D(_0170_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[14][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][13]$_DFFE_PP_  (.D(_0171_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[14][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][14]$_DFFE_PP_  (.D(_0172_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[14][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][15]$_DFFE_PP_  (.D(_0173_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[14][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][16]$_DFFE_PP_  (.D(_0174_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[14][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][17]$_DFFE_PP_  (.D(_0175_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[14][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][18]$_DFFE_PP_  (.D(_0176_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[14][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][19]$_DFFE_PP_  (.D(_0177_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[14][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][1]$_DFFE_PP_  (.D(_0178_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[14][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][20]$_DFFE_PP_  (.D(_0179_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[14][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][21]$_DFFE_PP_  (.D(_0180_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[14][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][22]$_DFFE_PP_  (.D(_0181_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[14][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][23]$_DFFE_PP_  (.D(_0182_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[14][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][24]$_DFFE_PP_  (.D(_0183_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[14][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][25]$_DFFE_PP_  (.D(_0184_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[14][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][26]$_DFFE_PP_  (.D(_0185_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[14][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][27]$_DFFE_PP_  (.D(_0186_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[14][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][28]$_DFFE_PP_  (.D(_0187_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[14][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][29]$_DFFE_PP_  (.D(_0188_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[14][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][2]$_DFFE_PP_  (.D(_0189_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[14][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][30]$_DFFE_PP_  (.D(_0190_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[14][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][31]$_DFFE_PP_  (.D(_0191_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[14][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][3]$_DFFE_PP_  (.D(_0192_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[14][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][4]$_DFFE_PP_  (.D(_0193_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[14][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][5]$_DFFE_PP_  (.D(_0194_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[14][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][6]$_DFFE_PP_  (.D(_0195_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[14][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][7]$_DFFE_PP_  (.D(_0196_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[14][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][8]$_DFFE_PP_  (.D(_0197_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[14][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][9]$_DFFE_PP_  (.D(_0198_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[14][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][0]$_DFFE_PP_  (.D(_0199_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[15][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][10]$_DFFE_PP_  (.D(_0200_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[15][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][11]$_DFFE_PP_  (.D(_0201_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[15][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][12]$_DFFE_PP_  (.D(_0202_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[15][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][13]$_DFFE_PP_  (.D(_0203_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[15][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][14]$_DFFE_PP_  (.D(_0204_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[15][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][15]$_DFFE_PP_  (.D(_0205_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[15][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][16]$_DFFE_PP_  (.D(_0206_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[15][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][17]$_DFFE_PP_  (.D(_0207_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[15][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][18]$_DFFE_PP_  (.D(_0208_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[15][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][19]$_DFFE_PP_  (.D(_0209_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[15][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][1]$_DFFE_PP_  (.D(_0210_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[15][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][20]$_DFFE_PP_  (.D(_0211_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[15][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][21]$_DFFE_PP_  (.D(_0212_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[15][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][22]$_DFFE_PP_  (.D(_0213_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[15][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][23]$_DFFE_PP_  (.D(_0214_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[15][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][24]$_DFFE_PP_  (.D(_0215_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[15][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][25]$_DFFE_PP_  (.D(_0216_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[15][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][26]$_DFFE_PP_  (.D(_0217_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[15][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][27]$_DFFE_PP_  (.D(_0218_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[15][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][28]$_DFFE_PP_  (.D(_0219_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[15][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][29]$_DFFE_PP_  (.D(_0220_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[15][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][2]$_DFFE_PP_  (.D(_0221_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[15][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][30]$_DFFE_PP_  (.D(_0222_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[15][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][31]$_DFFE_PP_  (.D(_0223_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[15][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][3]$_DFFE_PP_  (.D(_0224_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[15][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][4]$_DFFE_PP_  (.D(_0225_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[15][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][5]$_DFFE_PP_  (.D(_0226_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[15][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][6]$_DFFE_PP_  (.D(_0227_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[15][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][7]$_DFFE_PP_  (.D(_0228_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[15][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][8]$_DFFE_PP_  (.D(_0229_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[15][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][9]$_DFFE_PP_  (.D(_0230_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[15][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][0]$_DFFE_PP_  (.D(_0231_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][10]$_DFFE_PP_  (.D(_0232_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][11]$_DFFE_PP_  (.D(_0233_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][12]$_DFFE_PP_  (.D(_0234_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][13]$_DFFE_PP_  (.D(_0235_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][14]$_DFFE_PP_  (.D(_0236_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][15]$_DFFE_PP_  (.D(_0237_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][16]$_DFFE_PP_  (.D(_0238_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][17]$_DFFE_PP_  (.D(_0239_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][18]$_DFFE_PP_  (.D(_0240_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][19]$_DFFE_PP_  (.D(_0241_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][1]$_DFFE_PP_  (.D(_0242_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][20]$_DFFE_PP_  (.D(_0243_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][21]$_DFFE_PP_  (.D(_0244_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][22]$_DFFE_PP_  (.D(_0245_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][23]$_DFFE_PP_  (.D(_0246_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][24]$_DFFE_PP_  (.D(_0247_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][25]$_DFFE_PP_  (.D(_0248_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][26]$_DFFE_PP_  (.D(_0249_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][27]$_DFFE_PP_  (.D(_0250_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][28]$_DFFE_PP_  (.D(_0251_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][29]$_DFFE_PP_  (.D(_0252_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][2]$_DFFE_PP_  (.D(_0253_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][30]$_DFFE_PP_  (.D(_0254_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][31]$_DFFE_PP_  (.D(_0255_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][3]$_DFFE_PP_  (.D(_0256_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][4]$_DFFE_PP_  (.D(_0257_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][5]$_DFFE_PP_  (.D(_0258_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][6]$_DFFE_PP_  (.D(_0259_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][7]$_DFFE_PP_  (.D(_0260_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][8]$_DFFE_PP_  (.D(_0261_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][9]$_DFFE_PP_  (.D(_0262_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][0]$_DFFE_PP_  (.D(_0263_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][10]$_DFFE_PP_  (.D(_0264_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][11]$_DFFE_PP_  (.D(_0265_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][12]$_DFFE_PP_  (.D(_0266_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][13]$_DFFE_PP_  (.D(_0267_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][14]$_DFFE_PP_  (.D(_0268_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][15]$_DFFE_PP_  (.D(_0269_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][16]$_DFFE_PP_  (.D(_0270_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][17]$_DFFE_PP_  (.D(_0271_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][18]$_DFFE_PP_  (.D(_0272_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][19]$_DFFE_PP_  (.D(_0273_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][1]$_DFFE_PP_  (.D(_0274_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][20]$_DFFE_PP_  (.D(_0275_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][21]$_DFFE_PP_  (.D(_0276_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][22]$_DFFE_PP_  (.D(_0277_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][23]$_DFFE_PP_  (.D(_0278_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][24]$_DFFE_PP_  (.D(_0279_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][25]$_DFFE_PP_  (.D(_0280_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][26]$_DFFE_PP_  (.D(_0281_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][27]$_DFFE_PP_  (.D(_0282_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][28]$_DFFE_PP_  (.D(_0283_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][29]$_DFFE_PP_  (.D(_0284_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][2]$_DFFE_PP_  (.D(_0285_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][30]$_DFFE_PP_  (.D(_0286_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][31]$_DFFE_PP_  (.D(_0287_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][3]$_DFFE_PP_  (.D(_0288_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][4]$_DFFE_PP_  (.D(_0289_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][5]$_DFFE_PP_  (.D(_0290_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][6]$_DFFE_PP_  (.D(_0291_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][7]$_DFFE_PP_  (.D(_0292_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][8]$_DFFE_PP_  (.D(_0293_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][9]$_DFFE_PP_  (.D(_0294_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][0]$_DFFE_PP_  (.D(_0295_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][10]$_DFFE_PP_  (.D(_0296_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][11]$_DFFE_PP_  (.D(_0297_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][12]$_DFFE_PP_  (.D(_0298_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][13]$_DFFE_PP_  (.D(_0299_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][14]$_DFFE_PP_  (.D(_0300_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][15]$_DFFE_PP_  (.D(_0301_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][16]$_DFFE_PP_  (.D(_0302_),
    .CLK(clknet_leaf_20_clk),
    .Q(\mem[3][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][17]$_DFFE_PP_  (.D(_0303_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[3][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][18]$_DFFE_PP_  (.D(_0304_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[3][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][19]$_DFFE_PP_  (.D(_0305_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[3][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][1]$_DFFE_PP_  (.D(_0306_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][20]$_DFFE_PP_  (.D(_0307_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[3][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][21]$_DFFE_PP_  (.D(_0308_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[3][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][22]$_DFFE_PP_  (.D(_0309_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[3][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][23]$_DFFE_PP_  (.D(_0310_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[3][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][24]$_DFFE_PP_  (.D(_0311_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[3][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][25]$_DFFE_PP_  (.D(_0312_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[3][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][26]$_DFFE_PP_  (.D(_0313_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[3][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][27]$_DFFE_PP_  (.D(_0314_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[3][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][28]$_DFFE_PP_  (.D(_0315_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[3][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][29]$_DFFE_PP_  (.D(_0316_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[3][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][2]$_DFFE_PP_  (.D(_0317_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][30]$_DFFE_PP_  (.D(_0318_),
    .CLK(clknet_leaf_6_clk),
    .Q(\mem[3][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][31]$_DFFE_PP_  (.D(_0319_),
    .CLK(clknet_leaf_7_clk),
    .Q(\mem[3][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][3]$_DFFE_PP_  (.D(_0320_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][4]$_DFFE_PP_  (.D(_0321_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][5]$_DFFE_PP_  (.D(_0322_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][6]$_DFFE_PP_  (.D(_0323_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][7]$_DFFE_PP_  (.D(_0324_),
    .CLK(clknet_leaf_1_clk),
    .Q(\mem[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][8]$_DFFE_PP_  (.D(_0325_),
    .CLK(clknet_leaf_21_clk),
    .Q(\mem[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][9]$_DFFE_PP_  (.D(_0326_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][0]$_DFFE_PP_  (.D(_0327_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][10]$_DFFE_PP_  (.D(_0328_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][11]$_DFFE_PP_  (.D(_0329_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][12]$_DFFE_PP_  (.D(_0330_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][13]$_DFFE_PP_  (.D(net203),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][14]$_DFFE_PP_  (.D(net209),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][15]$_DFFE_PP_  (.D(_0333_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][16]$_DFFE_PP_  (.D(net215),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[4][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][17]$_DFFE_PP_  (.D(_0335_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[4][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][18]$_DFFE_PP_  (.D(_0336_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[4][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][19]$_DFFE_PP_  (.D(_0337_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[4][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][1]$_DFFE_PP_  (.D(_0338_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][20]$_DFFE_PP_  (.D(_0339_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[4][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][21]$_DFFE_PP_  (.D(_0340_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[4][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][22]$_DFFE_PP_  (.D(_0341_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[4][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][23]$_DFFE_PP_  (.D(_0342_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[4][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][24]$_DFFE_PP_  (.D(_0343_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[4][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][25]$_DFFE_PP_  (.D(_0344_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[4][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][26]$_DFFE_PP_  (.D(_0345_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[4][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][27]$_DFFE_PP_  (.D(_0346_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[4][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][28]$_DFFE_PP_  (.D(_0347_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[4][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][29]$_DFFE_PP_  (.D(_0348_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[4][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][2]$_DFFE_PP_  (.D(_0349_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][30]$_DFFE_PP_  (.D(_0350_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[4][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][31]$_DFFE_PP_  (.D(net158),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[4][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][3]$_DFFE_PP_  (.D(_0352_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][4]$_DFFE_PP_  (.D(net184),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][5]$_DFFE_PP_  (.D(_0354_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][6]$_DFFE_PP_  (.D(_0355_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][7]$_DFFE_PP_  (.D(_0356_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][8]$_DFFE_PP_  (.D(_0357_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][9]$_DFFE_PP_  (.D(_0358_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][0]$_DFFE_PP_  (.D(net226),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][10]$_DFFE_PP_  (.D(_0360_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][11]$_DFFE_PP_  (.D(net206),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][12]$_DFFE_PP_  (.D(net200),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][13]$_DFFE_PP_  (.D(_0363_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][14]$_DFFE_PP_  (.D(_0364_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][15]$_DFFE_PP_  (.D(_0365_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][16]$_DFFE_PP_  (.D(_0366_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[5][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][17]$_DFFE_PP_  (.D(_0367_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[5][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][18]$_DFFE_PP_  (.D(_0368_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[5][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][19]$_DFFE_PP_  (.D(_0369_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[5][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][1]$_DFFE_PP_  (.D(net160),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][20]$_DFFE_PP_  (.D(_0371_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[5][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][21]$_DFFE_PP_  (.D(_0372_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[5][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][22]$_DFFE_PP_  (.D(net212),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[5][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][23]$_DFFE_PP_  (.D(_0374_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[5][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][24]$_DFFE_PP_  (.D(net239),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[5][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][25]$_DFFE_PP_  (.D(_0376_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[5][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][26]$_DFFE_PP_  (.D(_0377_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[5][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][27]$_DFFE_PP_  (.D(net164),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[5][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][28]$_DFFE_PP_  (.D(_0379_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[5][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][29]$_DFFE_PP_  (.D(_0380_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[5][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][2]$_DFFE_PP_  (.D(_0381_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][30]$_DFFE_PP_  (.D(_0382_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[5][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][31]$_DFFE_PP_  (.D(_0383_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[5][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][3]$_DFFE_PP_  (.D(_0384_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][4]$_DFFE_PP_  (.D(_0385_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][5]$_DFFE_PP_  (.D(_0386_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][6]$_DFFE_PP_  (.D(net186),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][7]$_DFFE_PP_  (.D(_0388_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][8]$_DFFE_PP_  (.D(_0389_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][9]$_DFFE_PP_  (.D(_0390_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][0]$_DFFE_PP_  (.D(_0391_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][10]$_DFFE_PP_  (.D(net218),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][11]$_DFFE_PP_  (.D(_0393_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][12]$_DFFE_PP_  (.D(_0394_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][13]$_DFFE_PP_  (.D(_0395_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][14]$_DFFE_PP_  (.D(_0396_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][15]$_DFFE_PP_  (.D(net224),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][16]$_DFFE_PP_  (.D(_0398_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[6][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][17]$_DFFE_PP_  (.D(_0399_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[6][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][18]$_DFFE_PP_  (.D(_0400_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[6][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][19]$_DFFE_PP_  (.D(_0401_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[6][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][1]$_DFFE_PP_  (.D(_0402_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][20]$_DFFE_PP_  (.D(_0403_),
    .CLK(clknet_leaf_9_clk),
    .Q(\mem[6][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][21]$_DFFE_PP_  (.D(net155),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[6][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][22]$_DFFE_PP_  (.D(_0405_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[6][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][23]$_DFFE_PP_  (.D(_0406_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[6][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][24]$_DFFE_PP_  (.D(_0407_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[6][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][25]$_DFFE_PP_  (.D(net181),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[6][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][26]$_DFFE_PP_  (.D(_0409_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[6][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][27]$_DFFE_PP_  (.D(_0410_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[6][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][28]$_DFFE_PP_  (.D(net194),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[6][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][29]$_DFFE_PP_  (.D(net176),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[6][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][2]$_DFFE_PP_  (.D(net196),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][30]$_DFFE_PP_  (.D(_0414_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[6][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][31]$_DFFE_PP_  (.D(_0415_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[6][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][3]$_DFFE_PP_  (.D(_0416_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][4]$_DFFE_PP_  (.D(_0417_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][5]$_DFFE_PP_  (.D(_0418_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][6]$_DFFE_PP_  (.D(_0419_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][7]$_DFFE_PP_  (.D(_0420_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][8]$_DFFE_PP_  (.D(_0421_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][9]$_DFFE_PP_  (.D(net236),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][0]$_DFFE_PP_  (.D(_0423_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][10]$_DFFE_PP_  (.D(_0424_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][11]$_DFFE_PP_  (.D(_0425_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][12]$_DFFE_PP_  (.D(_0426_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][13]$_DFFE_PP_  (.D(_0427_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][14]$_DFFE_PP_  (.D(_0428_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][15]$_DFFE_PP_  (.D(_0429_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][16]$_DFFE_PP_  (.D(_0430_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[7][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][17]$_DFFE_PP_  (.D(_0431_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[7][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][18]$_DFFE_PP_  (.D(_0432_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[7][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][19]$_DFFE_PP_  (.D(_0433_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[7][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][1]$_DFFE_PP_  (.D(_0434_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][20]$_DFFE_PP_  (.D(net190),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[7][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][21]$_DFFE_PP_  (.D(_0436_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[7][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][22]$_DFFE_PP_  (.D(_0437_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[7][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][23]$_DFFE_PP_  (.D(net152),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[7][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][24]$_DFFE_PP_  (.D(_0439_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[7][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][25]$_DFFE_PP_  (.D(_0440_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[7][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][26]$_DFFE_PP_  (.D(_0441_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[7][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][27]$_DFFE_PP_  (.D(_0442_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[7][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][28]$_DFFE_PP_  (.D(_0443_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[7][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][29]$_DFFE_PP_  (.D(_0444_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[7][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][2]$_DFFE_PP_  (.D(_0445_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][30]$_DFFE_PP_  (.D(net168),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[7][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][31]$_DFFE_PP_  (.D(_0447_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[7][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][3]$_DFFE_PP_  (.D(_0448_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][4]$_DFFE_PP_  (.D(_0449_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][5]$_DFFE_PP_  (.D(_0450_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][6]$_DFFE_PP_  (.D(_0451_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][7]$_DFFE_PP_  (.D(_0452_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][8]$_DFFE_PP_  (.D(_0453_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][9]$_DFFE_PP_  (.D(_0454_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][0]$_DFFE_PP_  (.D(_0455_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[8][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][10]$_DFFE_PP_  (.D(_0456_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[8][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][11]$_DFFE_PP_  (.D(_0457_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[8][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][12]$_DFFE_PP_  (.D(_0458_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[8][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][13]$_DFFE_PP_  (.D(_0459_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[8][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][14]$_DFFE_PP_  (.D(_0460_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[8][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][15]$_DFFE_PP_  (.D(_0461_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[8][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][16]$_DFFE_PP_  (.D(_0462_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[8][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][17]$_DFFE_PP_  (.D(net232),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[8][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][18]$_DFFE_PP_  (.D(net221),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[8][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][19]$_DFFE_PP_  (.D(net172),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[8][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][1]$_DFFE_PP_  (.D(_0466_),
    .CLK(clknet_leaf_13_clk),
    .Q(\mem[8][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][20]$_DFFE_PP_  (.D(_0467_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[8][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][21]$_DFFE_PP_  (.D(_0468_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[8][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][22]$_DFFE_PP_  (.D(_0469_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[8][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][23]$_DFFE_PP_  (.D(_0470_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[8][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][24]$_DFFE_PP_  (.D(_0471_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[8][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][25]$_DFFE_PP_  (.D(_0472_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[8][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][26]$_DFFE_PP_  (.D(net149),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[8][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][27]$_DFFE_PP_  (.D(_0474_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[8][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][28]$_DFFE_PP_  (.D(_0475_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[8][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][29]$_DFFE_PP_  (.D(_0476_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[8][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][2]$_DFFE_PP_  (.D(_0477_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[8][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][30]$_DFFE_PP_  (.D(_0478_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[8][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][31]$_DFFE_PP_  (.D(_0479_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[8][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][3]$_DFFE_PP_  (.D(_0480_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[8][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][4]$_DFFE_PP_  (.D(_0481_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[8][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][5]$_DFFE_PP_  (.D(_0482_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[8][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][6]$_DFFE_PP_  (.D(_0483_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[8][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][7]$_DFFE_PP_  (.D(_0484_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[8][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][8]$_DFFE_PP_  (.D(net242),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[8][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][9]$_DFFE_PP_  (.D(_0486_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[8][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][0]$_DFFE_PP_  (.D(_0487_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[9][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][10]$_DFFE_PP_  (.D(_0488_),
    .CLK(clknet_leaf_23_clk),
    .Q(\mem[9][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][11]$_DFFE_PP_  (.D(_0489_),
    .CLK(clknet_leaf_22_clk),
    .Q(\mem[9][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][12]$_DFFE_PP_  (.D(_0490_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[9][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][13]$_DFFE_PP_  (.D(_0491_),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem[9][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][14]$_DFFE_PP_  (.D(_0492_),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem[9][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][15]$_DFFE_PP_  (.D(_0493_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[9][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][16]$_DFFE_PP_  (.D(_0494_),
    .CLK(clknet_leaf_17_clk),
    .Q(\mem[9][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][17]$_DFFE_PP_  (.D(_0495_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[9][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][18]$_DFFE_PP_  (.D(_0496_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[9][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][19]$_DFFE_PP_  (.D(_0497_),
    .CLK(clknet_leaf_16_clk),
    .Q(\mem[9][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][1]$_DFFE_PP_  (.D(_0498_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[9][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][20]$_DFFE_PP_  (.D(_0499_),
    .CLK(clknet_leaf_8_clk),
    .Q(\mem[9][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][21]$_DFFE_PP_  (.D(_0500_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[9][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][22]$_DFFE_PP_  (.D(_0501_),
    .CLK(clknet_leaf_14_clk),
    .Q(\mem[9][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][23]$_DFFE_PP_  (.D(_0502_),
    .CLK(clknet_leaf_12_clk),
    .Q(\mem[9][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][24]$_DFFE_PP_  (.D(_0503_),
    .CLK(clknet_leaf_15_clk),
    .Q(\mem[9][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][25]$_DFFE_PP_  (.D(_0504_),
    .CLK(clknet_leaf_11_clk),
    .Q(\mem[9][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][26]$_DFFE_PP_  (.D(_0505_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[9][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][27]$_DFFE_PP_  (.D(_0506_),
    .CLK(clknet_leaf_10_clk),
    .Q(\mem[9][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][28]$_DFFE_PP_  (.D(_0507_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[9][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][29]$_DFFE_PP_  (.D(_0508_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[9][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][2]$_DFFE_PP_  (.D(_0509_),
    .CLK(clknet_leaf_5_clk),
    .Q(\mem[9][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][30]$_DFFE_PP_  (.D(_0510_),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[9][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][31]$_DFFE_PP_  (.D(_0511_),
    .CLK(clknet_leaf_3_clk),
    .Q(\mem[9][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][3]$_DFFE_PP_  (.D(net162),
    .CLK(clknet_leaf_4_clk),
    .Q(\mem[9][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][4]$_DFFE_PP_  (.D(_0513_),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[9][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][5]$_DFFE_PP_  (.D(net179),
    .CLK(clknet_leaf_2_clk),
    .Q(\mem[9][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][6]$_DFFE_PP_  (.D(_0515_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[9][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][7]$_DFFE_PP_  (.D(net229),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[9][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][8]$_DFFE_PP_  (.D(_0517_),
    .CLK(clknet_leaf_0_clk),
    .Q(\mem[9][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][9]$_DFFE_PP_  (.D(_0518_),
    .CLK(clknet_leaf_24_clk),
    .Q(\mem[9][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][0]$_DFFE_PN0P_  (.D(_0519_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net79));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][10]$_DFFE_PN0P_  (.D(_0520_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net80));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][11]$_DFFE_PN0P_  (.D(_0521_),
    .RN(net1),
    .CLK(clknet_leaf_19_clk),
    .Q(net81));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][12]$_DFFE_PN0P_  (.D(_0522_),
    .RN(net1),
    .CLK(clknet_leaf_19_clk),
    .Q(net82));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][13]$_DFFE_PN0P_  (.D(_0523_),
    .RN(net1),
    .CLK(clknet_leaf_19_clk),
    .Q(net83));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][14]$_DFFE_PN0P_  (.D(_0524_),
    .RN(net1),
    .CLK(clknet_leaf_18_clk),
    .Q(net84));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][15]$_DFFE_PN0P_  (.D(_0525_),
    .RN(net1),
    .CLK(clknet_leaf_17_clk),
    .Q(net85));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][16]$_DFFE_PN0P_  (.D(_0526_),
    .RN(net1),
    .CLK(clknet_leaf_17_clk),
    .Q(net86));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][17]$_DFFE_PN0P_  (.D(_0527_),
    .RN(net1),
    .CLK(clknet_leaf_17_clk),
    .Q(net87));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][18]$_DFFE_PN0P_  (.D(_0528_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net88));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][19]$_DFFE_PN0P_  (.D(_0529_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net89));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][1]$_DFFE_PN0P_  (.D(_0530_),
    .RN(net1),
    .CLK(clknet_leaf_13_clk),
    .Q(net90));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][20]$_DFFE_PN0P_  (.D(_0531_),
    .RN(net1),
    .CLK(clknet_leaf_10_clk),
    .Q(net91));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][21]$_DFFE_PN0P_  (.D(_0532_),
    .RN(net1),
    .CLK(clknet_leaf_12_clk),
    .Q(net92));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][22]$_DFFE_PN0P_  (.D(_0533_),
    .RN(net1),
    .CLK(clknet_leaf_10_clk),
    .Q(net93));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][23]$_DFFE_PN0P_  (.D(_0534_),
    .RN(net1),
    .CLK(clknet_leaf_11_clk),
    .Q(net94));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][24]$_DFFE_PN0P_  (.D(_0535_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net95));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][25]$_DFFE_PN0P_  (.D(_0536_),
    .RN(net1),
    .CLK(clknet_leaf_10_clk),
    .Q(net96));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][26]$_DFFE_PN0P_  (.D(_0537_),
    .RN(net1),
    .CLK(clknet_leaf_10_clk),
    .Q(net97));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][27]$_DFFE_PN0P_  (.D(_0538_),
    .RN(net1),
    .CLK(clknet_leaf_7_clk),
    .Q(net98));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][28]$_DFFE_PN0P_  (.D(_0539_),
    .RN(net1),
    .CLK(clknet_leaf_6_clk),
    .Q(net99));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][29]$_DFFE_PN0P_  (.D(_0540_),
    .RN(net1),
    .CLK(clknet_leaf_4_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][2]$_DFFE_PN0P_  (.D(_0541_),
    .RN(net1),
    .CLK(clknet_leaf_4_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][30]$_DFFE_PN0P_  (.D(_0542_),
    .RN(net1),
    .CLK(clknet_leaf_4_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][31]$_DFFE_PN0P_  (.D(_0543_),
    .RN(net1),
    .CLK(clknet_leaf_3_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][3]$_DFFE_PN0P_  (.D(_0544_),
    .RN(net1),
    .CLK(clknet_leaf_3_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][4]$_DFFE_PN0P_  (.D(_0545_),
    .RN(net1),
    .CLK(clknet_leaf_6_clk),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][5]$_DFFE_PN0P_  (.D(_0546_),
    .RN(net1),
    .CLK(clknet_leaf_3_clk),
    .Q(net134));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][6]$_DFFE_PN0P_  (.D(_0547_),
    .RN(net1),
    .CLK(clknet_leaf_6_clk),
    .Q(net139));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][7]$_DFFE_PN0P_  (.D(_0548_),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(net140));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][8]$_DFFE_PN0P_  (.D(_0549_),
    .RN(net1),
    .CLK(clknet_leaf_21_clk),
    .Q(net141));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[0][9]$_DFFE_PN0P_  (.D(_0550_),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(net142));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][0]$_DFFE_PN0P_  (.D(_0551_),
    .RN(net1),
    .CLK(clknet_leaf_22_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][10]$_DFFE_PN0P_  (.D(_0552_),
    .RN(net1),
    .CLK(clknet_leaf_22_clk),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][11]$_DFFE_PN0P_  (.D(_0553_),
    .RN(net1),
    .CLK(clknet_leaf_20_clk),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][12]$_DFFE_PN0P_  (.D(_0554_),
    .RN(net1),
    .CLK(clknet_leaf_20_clk),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][13]$_DFFE_PN0P_  (.D(_0555_),
    .RN(net1),
    .CLK(clknet_leaf_18_clk),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][14]$_DFFE_PN0P_  (.D(_0556_),
    .RN(net1),
    .CLK(clknet_leaf_18_clk),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][15]$_DFFE_PN0P_  (.D(_0557_),
    .RN(net1),
    .CLK(clknet_leaf_17_clk),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][16]$_DFFE_PN0P_  (.D(_0558_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][17]$_DFFE_PN0P_  (.D(_0559_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][18]$_DFFE_PN0P_  (.D(_0560_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][19]$_DFFE_PN0P_  (.D(_0561_),
    .RN(net1),
    .CLK(clknet_leaf_16_clk),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][1]$_DFFE_PN0P_  (.D(_0562_),
    .RN(net1),
    .CLK(clknet_leaf_13_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][20]$_DFFE_PN0P_  (.D(_0563_),
    .RN(net1),
    .CLK(clknet_leaf_8_clk),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][21]$_DFFE_PN0P_  (.D(_0564_),
    .RN(net1),
    .CLK(clknet_leaf_12_clk),
    .Q(net127));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][22]$_DFFE_PN0P_  (.D(_0565_),
    .RN(net1),
    .CLK(clknet_leaf_14_clk),
    .Q(net128));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][23]$_DFFE_PN0P_  (.D(_0566_),
    .RN(net1),
    .CLK(clknet_leaf_12_clk),
    .Q(net129));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][24]$_DFFE_PN0P_  (.D(_0567_),
    .RN(net1),
    .CLK(clknet_leaf_15_clk),
    .Q(net130));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][25]$_DFFE_PN0P_  (.D(_0568_),
    .RN(net1),
    .CLK(clknet_leaf_11_clk),
    .Q(net131));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][26]$_DFFE_PN0P_  (.D(_0569_),
    .RN(net1),
    .CLK(clknet_leaf_11_clk),
    .Q(net132));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][27]$_DFFE_PN0P_  (.D(_0570_),
    .RN(net1),
    .CLK(clknet_leaf_10_clk),
    .Q(net133));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][28]$_DFFE_PN0P_  (.D(_0571_),
    .RN(net1),
    .CLK(clknet_leaf_7_clk),
    .Q(net135));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][29]$_DFFE_PN0P_  (.D(_0572_),
    .RN(net1),
    .CLK(clknet_leaf_7_clk),
    .Q(net136));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][2]$_DFFE_PN0P_  (.D(_0573_),
    .RN(net1),
    .CLK(clknet_leaf_6_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][30]$_DFFE_PN0P_  (.D(_0574_),
    .RN(net1),
    .CLK(clknet_leaf_6_clk),
    .Q(net137));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][31]$_DFFE_PN0P_  (.D(_0575_),
    .RN(net1),
    .CLK(clknet_leaf_8_clk),
    .Q(net138));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][3]$_DFFE_PN0P_  (.D(_0576_),
    .RN(net1),
    .CLK(clknet_leaf_2_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][4]$_DFFE_PN0P_  (.D(_0577_),
    .RN(net1),
    .CLK(clknet_leaf_8_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][5]$_DFFE_PN0P_  (.D(_0578_),
    .RN(net1),
    .CLK(clknet_leaf_1_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][6]$_DFFE_PN0P_  (.D(_0579_),
    .RN(net1),
    .CLK(clknet_leaf_1_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][7]$_DFFE_PN0P_  (.D(_0580_),
    .RN(net1),
    .CLK(clknet_leaf_0_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][8]$_DFFE_PN0P_  (.D(_0581_),
    .RN(net1),
    .CLK(clknet_leaf_21_clk),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data_regs[1][9]$_DFFE_PN0P_  (.D(_0582_),
    .RN(net1),
    .CLK(clknet_leaf_0_clk),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[0]$_DFFE_PN0N_  (.D(_0583_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(\rd_ptr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \rd_ptr[1]$_DFFE_PN0N_  (.D(_0584_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(\rd_ptr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[2]$_DFFE_PN0N_  (.D(_0585_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(\rd_ptr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr[3]$_DFFE_PN0N_  (.D(_0586_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(\rd_ptr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_valid_regs[0]$_DFF_PN0_  (.D(_0001_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net143));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_valid_regs[1]$_DFF_PN0_  (.D(_2731_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(net144));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[0]$_DFFE_PN0N_  (.D(_0587_),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(\wr_ptr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[1]$_DFFE_PN0N_  (.D(_0588_),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(\wr_ptr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[2]$_DFFE_PN0N_  (.D(_0589_),
    .RN(net1),
    .CLK(clknet_leaf_24_clk),
    .Q(\wr_ptr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr[3]$_DFFE_PN0N_  (.D(_0590_),
    .RN(net1),
    .CLK(clknet_leaf_23_clk),
    .Q(\wr_ptr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net147),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_640 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input1 (.I(rd_en[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(rd_en[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input3 (.I(net233),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input4 (.I(net219),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input5 (.I(net207),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input6 (.I(net201),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(net204),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(net210),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(net227),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input10 (.I(net216),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input11 (.I(net234),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(net222),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input13 (.I(net173),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(net166),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input15 (.I(net192),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input16 (.I(net156),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input17 (.I(net213),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input18 (.I(net153),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input19 (.I(net240),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(net191),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input21 (.I(net150),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(net170),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input23 (.I(net197),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input24 (.I(net177),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input25 (.I(net198),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input26 (.I(net169),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input27 (.I(net165),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input28 (.I(net225),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input29 (.I(net159),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input30 (.I(net195),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input31 (.I(net161),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input32 (.I(net183),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(net178),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input34 (.I(net185),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input35 (.I(net228),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input36 (.I(net174),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input37 (.I(net241),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input38 (.I(net235),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input39 (.I(net217),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input40 (.I(net205),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input41 (.I(net199),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input42 (.I(net202),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input43 (.I(net208),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(net223),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input45 (.I(net214),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input46 (.I(net231),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input47 (.I(net188),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input48 (.I(net220),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input49 (.I(net171),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input50 (.I(net189),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input51 (.I(net154),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input52 (.I(net211),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input53 (.I(net151),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input54 (.I(net238),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input55 (.I(net180),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input56 (.I(net148),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input57 (.I(net163),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input58 (.I(net182),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input59 (.I(net193),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input60 (.I(net175),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input61 (.I(net167),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input62 (.I(net157),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(net187),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input64 (.I(net230),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input65 (.I(net243),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input66 (.I(net237),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input67 (.I(wr_en[0]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input68 (.I(wr_en[1]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(almost_empty));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(almost_full));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net72),
    .Z(data_count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net73),
    .Z(data_count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net74),
    .Z(data_count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net75),
    .Z(data_count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net76),
    .Z(data_count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net77),
    .Z(empty));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net78),
    .Z(full));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net79),
    .Z(rd_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net80),
    .Z(rd_data[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net81),
    .Z(rd_data[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net82),
    .Z(rd_data[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net83),
    .Z(rd_data[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net84),
    .Z(rd_data[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net85),
    .Z(rd_data[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net86),
    .Z(rd_data[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net87),
    .Z(rd_data[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net88),
    .Z(rd_data[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net89),
    .Z(rd_data[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net90),
    .Z(rd_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net91),
    .Z(rd_data[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net92),
    .Z(rd_data[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net93),
    .Z(rd_data[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net94),
    .Z(rd_data[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net95),
    .Z(rd_data[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net96),
    .Z(rd_data[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net97),
    .Z(rd_data[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net98),
    .Z(rd_data[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net99),
    .Z(rd_data[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net100),
    .Z(rd_data[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net101),
    .Z(rd_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net102),
    .Z(rd_data[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net103),
    .Z(rd_data[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net104),
    .Z(rd_data[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net105),
    .Z(rd_data[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net106),
    .Z(rd_data[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net107),
    .Z(rd_data[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net108),
    .Z(rd_data[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net109),
    .Z(rd_data[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net110),
    .Z(rd_data[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net111),
    .Z(rd_data[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net112),
    .Z(rd_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output112 (.I(net113),
    .Z(rd_data[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output113 (.I(net114),
    .Z(rd_data[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output114 (.I(net115),
    .Z(rd_data[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output115 (.I(net116),
    .Z(rd_data[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output116 (.I(net117),
    .Z(rd_data[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output117 (.I(net118),
    .Z(rd_data[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output118 (.I(net119),
    .Z(rd_data[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output119 (.I(net120),
    .Z(rd_data[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output120 (.I(net121),
    .Z(rd_data[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output121 (.I(net122),
    .Z(rd_data[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output122 (.I(net123),
    .Z(rd_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output123 (.I(net124),
    .Z(rd_data[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output124 (.I(net125),
    .Z(rd_data[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output125 (.I(net126),
    .Z(rd_data[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output126 (.I(net127),
    .Z(rd_data[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output127 (.I(net128),
    .Z(rd_data[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output128 (.I(net129),
    .Z(rd_data[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output129 (.I(net130),
    .Z(rd_data[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output130 (.I(net131),
    .Z(rd_data[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output131 (.I(net132),
    .Z(rd_data[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output132 (.I(net133),
    .Z(rd_data[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output133 (.I(net134),
    .Z(rd_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output134 (.I(net135),
    .Z(rd_data[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output135 (.I(net136),
    .Z(rd_data[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output136 (.I(net137),
    .Z(rd_data[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output137 (.I(net138),
    .Z(rd_data[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output138 (.I(net139),
    .Z(rd_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output139 (.I(net140),
    .Z(rd_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output140 (.I(net141),
    .Z(rd_data[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output141 (.I(net142),
    .Z(rd_data[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output142 (.I(net143),
    .Z(rd_valid[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output143 (.I(net144),
    .Z(rd_valid[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output144 (.I(net145),
    .Z(wr_ready[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net146),
    .Z(wr_ready[1]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload1 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload2 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload3 (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload4 (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload5 (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload6 (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload7 (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload8 (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload9 (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 clkload10 (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload11 (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload12 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload13 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload14 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload15 (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload16 (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload17 (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload18 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 clkload19 (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload20 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload21 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload22 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload23 (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(wr_data[58]),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold4 (.I(_0473_),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold5 (.I(wr_data[26]),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold6 (.I(wr_data[55]),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold7 (.I(_0438_),
    .Z(net152));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold8 (.I(wr_data[23]),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold9 (.I(wr_data[53]),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold10 (.I(_0404_),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold11 (.I(wr_data[21]),
    .Z(net156));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold12 (.I(wr_data[63]),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold13 (.I(_0351_),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold14 (.I(wr_data[33]),
    .Z(net159));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold15 (.I(_0370_),
    .Z(net160));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold16 (.I(wr_data[35]),
    .Z(net161));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold17 (.I(_0512_),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold18 (.I(wr_data[59]),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold19 (.I(_0378_),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold20 (.I(wr_data[31]),
    .Z(net165));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold21 (.I(wr_data[1]),
    .Z(net166));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold22 (.I(wr_data[62]),
    .Z(net167));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold23 (.I(_0446_),
    .Z(net168));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold24 (.I(wr_data[30]),
    .Z(net169));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold25 (.I(wr_data[27]),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold26 (.I(wr_data[51]),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold27 (.I(_0465_),
    .Z(net172));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold28 (.I(wr_data[19]),
    .Z(net173));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold29 (.I(wr_data[3]),
    .Z(net174));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold30 (.I(wr_data[61]),
    .Z(net175));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold31 (.I(_0412_),
    .Z(net176));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold32 (.I(wr_data[29]),
    .Z(net177));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold33 (.I(wr_data[37]),
    .Z(net178));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold34 (.I(_0514_),
    .Z(net179));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold35 (.I(wr_data[57]),
    .Z(net180));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold36 (.I(_0408_),
    .Z(net181));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold37 (.I(wr_data[5]),
    .Z(net182));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold38 (.I(wr_data[36]),
    .Z(net183));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold39 (.I(_0353_),
    .Z(net184));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold40 (.I(wr_data[38]),
    .Z(net185));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold41 (.I(_0387_),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold42 (.I(wr_data[6]),
    .Z(net187));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold43 (.I(wr_data[4]),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold44 (.I(wr_data[52]),
    .Z(net189));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold45 (.I(_0435_),
    .Z(net190));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold46 (.I(wr_data[25]),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold47 (.I(wr_data[20]),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold48 (.I(wr_data[60]),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold49 (.I(_0411_),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold50 (.I(wr_data[34]),
    .Z(net195));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold51 (.I(_0413_),
    .Z(net196));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold52 (.I(wr_data[28]),
    .Z(net197));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold53 (.I(wr_data[2]),
    .Z(net198));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold54 (.I(wr_data[44]),
    .Z(net199));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold55 (.I(_0362_),
    .Z(net200));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold56 (.I(wr_data[12]),
    .Z(net201));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold57 (.I(wr_data[45]),
    .Z(net202));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold58 (.I(_0331_),
    .Z(net203));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold59 (.I(wr_data[13]),
    .Z(net204));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold60 (.I(wr_data[43]),
    .Z(net205));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold61 (.I(_0361_),
    .Z(net206));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold62 (.I(wr_data[11]),
    .Z(net207));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold63 (.I(wr_data[46]),
    .Z(net208));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold64 (.I(_0332_),
    .Z(net209));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold65 (.I(wr_data[14]),
    .Z(net210));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold66 (.I(wr_data[54]),
    .Z(net211));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold67 (.I(_0373_),
    .Z(net212));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold68 (.I(wr_data[22]),
    .Z(net213));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold69 (.I(wr_data[48]),
    .Z(net214));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold70 (.I(_0334_),
    .Z(net215));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold71 (.I(wr_data[16]),
    .Z(net216));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold72 (.I(wr_data[42]),
    .Z(net217));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold73 (.I(_0392_),
    .Z(net218));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold74 (.I(wr_data[10]),
    .Z(net219));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold75 (.I(wr_data[50]),
    .Z(net220));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold76 (.I(_0464_),
    .Z(net221));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold77 (.I(wr_data[18]),
    .Z(net222));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold78 (.I(wr_data[47]),
    .Z(net223));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold79 (.I(_0397_),
    .Z(net224));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold80 (.I(wr_data[32]),
    .Z(net225));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold81 (.I(_0359_),
    .Z(net226));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold82 (.I(wr_data[15]),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold83 (.I(wr_data[39]),
    .Z(net228));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold84 (.I(_0516_),
    .Z(net229));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold85 (.I(wr_data[7]),
    .Z(net230));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold86 (.I(wr_data[49]),
    .Z(net231));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold87 (.I(_0463_),
    .Z(net232));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold88 (.I(wr_data[0]),
    .Z(net233));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold89 (.I(wr_data[17]),
    .Z(net234));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold90 (.I(wr_data[41]),
    .Z(net235));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold91 (.I(_0422_),
    .Z(net236));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold92 (.I(wr_data[9]),
    .Z(net237));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold93 (.I(wr_data[56]),
    .Z(net238));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold94 (.I(_0375_),
    .Z(net239));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold95 (.I(wr_data[24]),
    .Z(net240));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold96 (.I(wr_data[40]),
    .Z(net241));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold97 (.I(_0485_),
    .Z(net242));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold98 (.I(wr_data[8]),
    .Z(net243));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net113));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net127));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net138));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_11 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1154 ();
endmodule
