module register_file (clk,
    read_en1,
    read_en2,
    rst_n,
    write_en,
    read_addr1,
    read_addr2,
    read_data1,
    read_data2,
    write_addr,
    write_data);
 input clk;
 input read_en1;
 input read_en2;
 input rst_n;
 input write_en;
 input [4:0] read_addr1;
 input [4:0] read_addr2;
 output [31:0] read_data1;
 output [31:0] read_data2;
 input [4:0] write_addr;
 input [31:0] write_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire \registers[0][0] ;
 wire \registers[0][10] ;
 wire \registers[0][11] ;
 wire \registers[0][12] ;
 wire \registers[0][13] ;
 wire \registers[0][14] ;
 wire \registers[0][15] ;
 wire \registers[0][16] ;
 wire \registers[0][17] ;
 wire \registers[0][18] ;
 wire \registers[0][19] ;
 wire \registers[0][1] ;
 wire \registers[0][20] ;
 wire \registers[0][21] ;
 wire \registers[0][22] ;
 wire \registers[0][23] ;
 wire \registers[0][24] ;
 wire \registers[0][25] ;
 wire \registers[0][26] ;
 wire \registers[0][27] ;
 wire \registers[0][28] ;
 wire \registers[0][29] ;
 wire \registers[0][2] ;
 wire \registers[0][30] ;
 wire \registers[0][31] ;
 wire \registers[0][3] ;
 wire \registers[0][4] ;
 wire \registers[0][5] ;
 wire \registers[0][6] ;
 wire \registers[0][7] ;
 wire \registers[0][8] ;
 wire \registers[0][9] ;
 wire \registers[10][0] ;
 wire \registers[10][10] ;
 wire \registers[10][11] ;
 wire \registers[10][12] ;
 wire \registers[10][13] ;
 wire \registers[10][14] ;
 wire \registers[10][15] ;
 wire \registers[10][16] ;
 wire \registers[10][17] ;
 wire \registers[10][18] ;
 wire \registers[10][19] ;
 wire \registers[10][1] ;
 wire \registers[10][20] ;
 wire \registers[10][21] ;
 wire \registers[10][22] ;
 wire \registers[10][23] ;
 wire \registers[10][24] ;
 wire \registers[10][25] ;
 wire \registers[10][26] ;
 wire \registers[10][27] ;
 wire \registers[10][28] ;
 wire \registers[10][29] ;
 wire \registers[10][2] ;
 wire \registers[10][30] ;
 wire \registers[10][31] ;
 wire \registers[10][3] ;
 wire \registers[10][4] ;
 wire \registers[10][5] ;
 wire \registers[10][6] ;
 wire \registers[10][7] ;
 wire \registers[10][8] ;
 wire \registers[10][9] ;
 wire \registers[11][0] ;
 wire \registers[11][10] ;
 wire \registers[11][11] ;
 wire \registers[11][12] ;
 wire \registers[11][13] ;
 wire \registers[11][14] ;
 wire \registers[11][15] ;
 wire \registers[11][16] ;
 wire \registers[11][17] ;
 wire \registers[11][18] ;
 wire \registers[11][19] ;
 wire \registers[11][1] ;
 wire \registers[11][20] ;
 wire \registers[11][21] ;
 wire \registers[11][22] ;
 wire \registers[11][23] ;
 wire \registers[11][24] ;
 wire \registers[11][25] ;
 wire \registers[11][26] ;
 wire \registers[11][27] ;
 wire \registers[11][28] ;
 wire \registers[11][29] ;
 wire \registers[11][2] ;
 wire \registers[11][30] ;
 wire \registers[11][31] ;
 wire \registers[11][3] ;
 wire \registers[11][4] ;
 wire \registers[11][5] ;
 wire \registers[11][6] ;
 wire \registers[11][7] ;
 wire \registers[11][8] ;
 wire \registers[11][9] ;
 wire \registers[12][0] ;
 wire \registers[12][10] ;
 wire \registers[12][11] ;
 wire \registers[12][12] ;
 wire \registers[12][13] ;
 wire \registers[12][14] ;
 wire \registers[12][15] ;
 wire \registers[12][16] ;
 wire \registers[12][17] ;
 wire \registers[12][18] ;
 wire \registers[12][19] ;
 wire \registers[12][1] ;
 wire \registers[12][20] ;
 wire \registers[12][21] ;
 wire \registers[12][22] ;
 wire \registers[12][23] ;
 wire \registers[12][24] ;
 wire \registers[12][25] ;
 wire \registers[12][26] ;
 wire \registers[12][27] ;
 wire \registers[12][28] ;
 wire \registers[12][29] ;
 wire \registers[12][2] ;
 wire \registers[12][30] ;
 wire \registers[12][31] ;
 wire \registers[12][3] ;
 wire \registers[12][4] ;
 wire \registers[12][5] ;
 wire \registers[12][6] ;
 wire \registers[12][7] ;
 wire \registers[12][8] ;
 wire \registers[12][9] ;
 wire \registers[13][0] ;
 wire \registers[13][10] ;
 wire \registers[13][11] ;
 wire \registers[13][12] ;
 wire \registers[13][13] ;
 wire \registers[13][14] ;
 wire \registers[13][15] ;
 wire \registers[13][16] ;
 wire \registers[13][17] ;
 wire \registers[13][18] ;
 wire \registers[13][19] ;
 wire \registers[13][1] ;
 wire \registers[13][20] ;
 wire \registers[13][21] ;
 wire \registers[13][22] ;
 wire \registers[13][23] ;
 wire \registers[13][24] ;
 wire \registers[13][25] ;
 wire \registers[13][26] ;
 wire \registers[13][27] ;
 wire \registers[13][28] ;
 wire \registers[13][29] ;
 wire \registers[13][2] ;
 wire \registers[13][30] ;
 wire \registers[13][31] ;
 wire \registers[13][3] ;
 wire \registers[13][4] ;
 wire \registers[13][5] ;
 wire \registers[13][6] ;
 wire \registers[13][7] ;
 wire \registers[13][8] ;
 wire \registers[13][9] ;
 wire \registers[14][0] ;
 wire \registers[14][10] ;
 wire \registers[14][11] ;
 wire \registers[14][12] ;
 wire \registers[14][13] ;
 wire \registers[14][14] ;
 wire \registers[14][15] ;
 wire \registers[14][16] ;
 wire \registers[14][17] ;
 wire \registers[14][18] ;
 wire \registers[14][19] ;
 wire \registers[14][1] ;
 wire \registers[14][20] ;
 wire \registers[14][21] ;
 wire \registers[14][22] ;
 wire \registers[14][23] ;
 wire \registers[14][24] ;
 wire \registers[14][25] ;
 wire \registers[14][26] ;
 wire \registers[14][27] ;
 wire \registers[14][28] ;
 wire \registers[14][29] ;
 wire \registers[14][2] ;
 wire \registers[14][30] ;
 wire \registers[14][31] ;
 wire \registers[14][3] ;
 wire \registers[14][4] ;
 wire \registers[14][5] ;
 wire \registers[14][6] ;
 wire \registers[14][7] ;
 wire \registers[14][8] ;
 wire \registers[14][9] ;
 wire \registers[15][0] ;
 wire \registers[15][10] ;
 wire \registers[15][11] ;
 wire \registers[15][12] ;
 wire \registers[15][13] ;
 wire \registers[15][14] ;
 wire \registers[15][15] ;
 wire \registers[15][16] ;
 wire \registers[15][17] ;
 wire \registers[15][18] ;
 wire \registers[15][19] ;
 wire \registers[15][1] ;
 wire \registers[15][20] ;
 wire \registers[15][21] ;
 wire \registers[15][22] ;
 wire \registers[15][23] ;
 wire \registers[15][24] ;
 wire \registers[15][25] ;
 wire \registers[15][26] ;
 wire \registers[15][27] ;
 wire \registers[15][28] ;
 wire \registers[15][29] ;
 wire \registers[15][2] ;
 wire \registers[15][30] ;
 wire \registers[15][31] ;
 wire \registers[15][3] ;
 wire \registers[15][4] ;
 wire \registers[15][5] ;
 wire \registers[15][6] ;
 wire \registers[15][7] ;
 wire \registers[15][8] ;
 wire \registers[15][9] ;
 wire \registers[16][0] ;
 wire \registers[16][10] ;
 wire \registers[16][11] ;
 wire \registers[16][12] ;
 wire \registers[16][13] ;
 wire \registers[16][14] ;
 wire \registers[16][15] ;
 wire \registers[16][16] ;
 wire \registers[16][17] ;
 wire \registers[16][18] ;
 wire \registers[16][19] ;
 wire \registers[16][1] ;
 wire \registers[16][20] ;
 wire \registers[16][21] ;
 wire \registers[16][22] ;
 wire \registers[16][23] ;
 wire \registers[16][24] ;
 wire \registers[16][25] ;
 wire \registers[16][26] ;
 wire \registers[16][27] ;
 wire \registers[16][28] ;
 wire \registers[16][29] ;
 wire \registers[16][2] ;
 wire \registers[16][30] ;
 wire \registers[16][31] ;
 wire \registers[16][3] ;
 wire \registers[16][4] ;
 wire \registers[16][5] ;
 wire \registers[16][6] ;
 wire \registers[16][7] ;
 wire \registers[16][8] ;
 wire \registers[16][9] ;
 wire \registers[17][0] ;
 wire \registers[17][10] ;
 wire \registers[17][11] ;
 wire \registers[17][12] ;
 wire \registers[17][13] ;
 wire \registers[17][14] ;
 wire \registers[17][15] ;
 wire \registers[17][16] ;
 wire \registers[17][17] ;
 wire \registers[17][18] ;
 wire \registers[17][19] ;
 wire \registers[17][1] ;
 wire \registers[17][20] ;
 wire \registers[17][21] ;
 wire \registers[17][22] ;
 wire \registers[17][23] ;
 wire \registers[17][24] ;
 wire \registers[17][25] ;
 wire \registers[17][26] ;
 wire \registers[17][27] ;
 wire \registers[17][28] ;
 wire \registers[17][29] ;
 wire \registers[17][2] ;
 wire \registers[17][30] ;
 wire \registers[17][31] ;
 wire \registers[17][3] ;
 wire \registers[17][4] ;
 wire \registers[17][5] ;
 wire \registers[17][6] ;
 wire \registers[17][7] ;
 wire \registers[17][8] ;
 wire \registers[17][9] ;
 wire \registers[18][0] ;
 wire \registers[18][10] ;
 wire \registers[18][11] ;
 wire \registers[18][12] ;
 wire \registers[18][13] ;
 wire \registers[18][14] ;
 wire \registers[18][15] ;
 wire \registers[18][16] ;
 wire \registers[18][17] ;
 wire \registers[18][18] ;
 wire \registers[18][19] ;
 wire \registers[18][1] ;
 wire \registers[18][20] ;
 wire \registers[18][21] ;
 wire \registers[18][22] ;
 wire \registers[18][23] ;
 wire \registers[18][24] ;
 wire \registers[18][25] ;
 wire \registers[18][26] ;
 wire \registers[18][27] ;
 wire \registers[18][28] ;
 wire \registers[18][29] ;
 wire \registers[18][2] ;
 wire \registers[18][30] ;
 wire \registers[18][31] ;
 wire \registers[18][3] ;
 wire \registers[18][4] ;
 wire \registers[18][5] ;
 wire \registers[18][6] ;
 wire \registers[18][7] ;
 wire \registers[18][8] ;
 wire \registers[18][9] ;
 wire \registers[19][0] ;
 wire \registers[19][10] ;
 wire \registers[19][11] ;
 wire \registers[19][12] ;
 wire \registers[19][13] ;
 wire \registers[19][14] ;
 wire \registers[19][15] ;
 wire \registers[19][16] ;
 wire \registers[19][17] ;
 wire \registers[19][18] ;
 wire \registers[19][19] ;
 wire \registers[19][1] ;
 wire \registers[19][20] ;
 wire \registers[19][21] ;
 wire \registers[19][22] ;
 wire \registers[19][23] ;
 wire \registers[19][24] ;
 wire \registers[19][25] ;
 wire \registers[19][26] ;
 wire \registers[19][27] ;
 wire \registers[19][28] ;
 wire \registers[19][29] ;
 wire \registers[19][2] ;
 wire \registers[19][30] ;
 wire \registers[19][31] ;
 wire \registers[19][3] ;
 wire \registers[19][4] ;
 wire \registers[19][5] ;
 wire \registers[19][6] ;
 wire \registers[19][7] ;
 wire \registers[19][8] ;
 wire \registers[19][9] ;
 wire \registers[1][0] ;
 wire \registers[1][10] ;
 wire \registers[1][11] ;
 wire \registers[1][12] ;
 wire \registers[1][13] ;
 wire \registers[1][14] ;
 wire \registers[1][15] ;
 wire \registers[1][16] ;
 wire \registers[1][17] ;
 wire \registers[1][18] ;
 wire \registers[1][19] ;
 wire \registers[1][1] ;
 wire \registers[1][20] ;
 wire \registers[1][21] ;
 wire \registers[1][22] ;
 wire \registers[1][23] ;
 wire \registers[1][24] ;
 wire \registers[1][25] ;
 wire \registers[1][26] ;
 wire \registers[1][27] ;
 wire \registers[1][28] ;
 wire \registers[1][29] ;
 wire \registers[1][2] ;
 wire \registers[1][30] ;
 wire \registers[1][31] ;
 wire \registers[1][3] ;
 wire \registers[1][4] ;
 wire \registers[1][5] ;
 wire \registers[1][6] ;
 wire \registers[1][7] ;
 wire \registers[1][8] ;
 wire \registers[1][9] ;
 wire \registers[20][0] ;
 wire \registers[20][10] ;
 wire \registers[20][11] ;
 wire \registers[20][12] ;
 wire \registers[20][13] ;
 wire \registers[20][14] ;
 wire \registers[20][15] ;
 wire \registers[20][16] ;
 wire \registers[20][17] ;
 wire \registers[20][18] ;
 wire \registers[20][19] ;
 wire \registers[20][1] ;
 wire \registers[20][20] ;
 wire \registers[20][21] ;
 wire \registers[20][22] ;
 wire \registers[20][23] ;
 wire \registers[20][24] ;
 wire \registers[20][25] ;
 wire \registers[20][26] ;
 wire \registers[20][27] ;
 wire \registers[20][28] ;
 wire \registers[20][29] ;
 wire \registers[20][2] ;
 wire \registers[20][30] ;
 wire \registers[20][31] ;
 wire \registers[20][3] ;
 wire \registers[20][4] ;
 wire \registers[20][5] ;
 wire \registers[20][6] ;
 wire \registers[20][7] ;
 wire \registers[20][8] ;
 wire \registers[20][9] ;
 wire \registers[21][0] ;
 wire \registers[21][10] ;
 wire \registers[21][11] ;
 wire \registers[21][12] ;
 wire \registers[21][13] ;
 wire \registers[21][14] ;
 wire \registers[21][15] ;
 wire \registers[21][16] ;
 wire \registers[21][17] ;
 wire \registers[21][18] ;
 wire \registers[21][19] ;
 wire \registers[21][1] ;
 wire \registers[21][20] ;
 wire \registers[21][21] ;
 wire \registers[21][22] ;
 wire \registers[21][23] ;
 wire \registers[21][24] ;
 wire \registers[21][25] ;
 wire \registers[21][26] ;
 wire \registers[21][27] ;
 wire \registers[21][28] ;
 wire \registers[21][29] ;
 wire \registers[21][2] ;
 wire \registers[21][30] ;
 wire \registers[21][31] ;
 wire \registers[21][3] ;
 wire \registers[21][4] ;
 wire \registers[21][5] ;
 wire \registers[21][6] ;
 wire \registers[21][7] ;
 wire \registers[21][8] ;
 wire \registers[21][9] ;
 wire \registers[22][0] ;
 wire \registers[22][10] ;
 wire \registers[22][11] ;
 wire \registers[22][12] ;
 wire \registers[22][13] ;
 wire \registers[22][14] ;
 wire \registers[22][15] ;
 wire \registers[22][16] ;
 wire \registers[22][17] ;
 wire \registers[22][18] ;
 wire \registers[22][19] ;
 wire \registers[22][1] ;
 wire \registers[22][20] ;
 wire \registers[22][21] ;
 wire \registers[22][22] ;
 wire \registers[22][23] ;
 wire \registers[22][24] ;
 wire \registers[22][25] ;
 wire \registers[22][26] ;
 wire \registers[22][27] ;
 wire \registers[22][28] ;
 wire \registers[22][29] ;
 wire \registers[22][2] ;
 wire \registers[22][30] ;
 wire \registers[22][31] ;
 wire \registers[22][3] ;
 wire \registers[22][4] ;
 wire \registers[22][5] ;
 wire \registers[22][6] ;
 wire \registers[22][7] ;
 wire \registers[22][8] ;
 wire \registers[22][9] ;
 wire \registers[23][0] ;
 wire \registers[23][10] ;
 wire \registers[23][11] ;
 wire \registers[23][12] ;
 wire \registers[23][13] ;
 wire \registers[23][14] ;
 wire \registers[23][15] ;
 wire \registers[23][16] ;
 wire \registers[23][17] ;
 wire \registers[23][18] ;
 wire \registers[23][19] ;
 wire \registers[23][1] ;
 wire \registers[23][20] ;
 wire \registers[23][21] ;
 wire \registers[23][22] ;
 wire \registers[23][23] ;
 wire \registers[23][24] ;
 wire \registers[23][25] ;
 wire \registers[23][26] ;
 wire \registers[23][27] ;
 wire \registers[23][28] ;
 wire \registers[23][29] ;
 wire \registers[23][2] ;
 wire \registers[23][30] ;
 wire \registers[23][31] ;
 wire \registers[23][3] ;
 wire \registers[23][4] ;
 wire \registers[23][5] ;
 wire \registers[23][6] ;
 wire \registers[23][7] ;
 wire \registers[23][8] ;
 wire \registers[23][9] ;
 wire \registers[24][0] ;
 wire \registers[24][10] ;
 wire \registers[24][11] ;
 wire \registers[24][12] ;
 wire \registers[24][13] ;
 wire \registers[24][14] ;
 wire \registers[24][15] ;
 wire \registers[24][16] ;
 wire \registers[24][17] ;
 wire \registers[24][18] ;
 wire \registers[24][19] ;
 wire \registers[24][1] ;
 wire \registers[24][20] ;
 wire \registers[24][21] ;
 wire \registers[24][22] ;
 wire \registers[24][23] ;
 wire \registers[24][24] ;
 wire \registers[24][25] ;
 wire \registers[24][26] ;
 wire \registers[24][27] ;
 wire \registers[24][28] ;
 wire \registers[24][29] ;
 wire \registers[24][2] ;
 wire \registers[24][30] ;
 wire \registers[24][31] ;
 wire \registers[24][3] ;
 wire \registers[24][4] ;
 wire \registers[24][5] ;
 wire \registers[24][6] ;
 wire \registers[24][7] ;
 wire \registers[24][8] ;
 wire \registers[24][9] ;
 wire \registers[25][0] ;
 wire \registers[25][10] ;
 wire \registers[25][11] ;
 wire \registers[25][12] ;
 wire \registers[25][13] ;
 wire \registers[25][14] ;
 wire \registers[25][15] ;
 wire \registers[25][16] ;
 wire \registers[25][17] ;
 wire \registers[25][18] ;
 wire \registers[25][19] ;
 wire \registers[25][1] ;
 wire \registers[25][20] ;
 wire \registers[25][21] ;
 wire \registers[25][22] ;
 wire \registers[25][23] ;
 wire \registers[25][24] ;
 wire \registers[25][25] ;
 wire \registers[25][26] ;
 wire \registers[25][27] ;
 wire \registers[25][28] ;
 wire \registers[25][29] ;
 wire \registers[25][2] ;
 wire \registers[25][30] ;
 wire \registers[25][31] ;
 wire \registers[25][3] ;
 wire \registers[25][4] ;
 wire \registers[25][5] ;
 wire \registers[25][6] ;
 wire \registers[25][7] ;
 wire \registers[25][8] ;
 wire \registers[25][9] ;
 wire \registers[26][0] ;
 wire \registers[26][10] ;
 wire \registers[26][11] ;
 wire \registers[26][12] ;
 wire \registers[26][13] ;
 wire \registers[26][14] ;
 wire \registers[26][15] ;
 wire \registers[26][16] ;
 wire \registers[26][17] ;
 wire \registers[26][18] ;
 wire \registers[26][19] ;
 wire \registers[26][1] ;
 wire \registers[26][20] ;
 wire \registers[26][21] ;
 wire \registers[26][22] ;
 wire \registers[26][23] ;
 wire \registers[26][24] ;
 wire \registers[26][25] ;
 wire \registers[26][26] ;
 wire \registers[26][27] ;
 wire \registers[26][28] ;
 wire \registers[26][29] ;
 wire \registers[26][2] ;
 wire \registers[26][30] ;
 wire \registers[26][31] ;
 wire \registers[26][3] ;
 wire \registers[26][4] ;
 wire \registers[26][5] ;
 wire \registers[26][6] ;
 wire \registers[26][7] ;
 wire \registers[26][8] ;
 wire \registers[26][9] ;
 wire \registers[27][0] ;
 wire \registers[27][10] ;
 wire \registers[27][11] ;
 wire \registers[27][12] ;
 wire \registers[27][13] ;
 wire \registers[27][14] ;
 wire \registers[27][15] ;
 wire \registers[27][16] ;
 wire \registers[27][17] ;
 wire \registers[27][18] ;
 wire \registers[27][19] ;
 wire \registers[27][1] ;
 wire \registers[27][20] ;
 wire \registers[27][21] ;
 wire \registers[27][22] ;
 wire \registers[27][23] ;
 wire \registers[27][24] ;
 wire \registers[27][25] ;
 wire \registers[27][26] ;
 wire \registers[27][27] ;
 wire \registers[27][28] ;
 wire \registers[27][29] ;
 wire \registers[27][2] ;
 wire \registers[27][30] ;
 wire \registers[27][31] ;
 wire \registers[27][3] ;
 wire \registers[27][4] ;
 wire \registers[27][5] ;
 wire \registers[27][6] ;
 wire \registers[27][7] ;
 wire \registers[27][8] ;
 wire \registers[27][9] ;
 wire \registers[28][0] ;
 wire \registers[28][10] ;
 wire \registers[28][11] ;
 wire \registers[28][12] ;
 wire \registers[28][13] ;
 wire \registers[28][14] ;
 wire \registers[28][15] ;
 wire \registers[28][16] ;
 wire \registers[28][17] ;
 wire \registers[28][18] ;
 wire \registers[28][19] ;
 wire \registers[28][1] ;
 wire \registers[28][20] ;
 wire \registers[28][21] ;
 wire \registers[28][22] ;
 wire \registers[28][23] ;
 wire \registers[28][24] ;
 wire \registers[28][25] ;
 wire \registers[28][26] ;
 wire \registers[28][27] ;
 wire \registers[28][28] ;
 wire \registers[28][29] ;
 wire \registers[28][2] ;
 wire \registers[28][30] ;
 wire \registers[28][31] ;
 wire \registers[28][3] ;
 wire \registers[28][4] ;
 wire \registers[28][5] ;
 wire \registers[28][6] ;
 wire \registers[28][7] ;
 wire \registers[28][8] ;
 wire \registers[28][9] ;
 wire \registers[29][0] ;
 wire \registers[29][10] ;
 wire \registers[29][11] ;
 wire \registers[29][12] ;
 wire \registers[29][13] ;
 wire \registers[29][14] ;
 wire \registers[29][15] ;
 wire \registers[29][16] ;
 wire \registers[29][17] ;
 wire \registers[29][18] ;
 wire \registers[29][19] ;
 wire \registers[29][1] ;
 wire \registers[29][20] ;
 wire \registers[29][21] ;
 wire \registers[29][22] ;
 wire \registers[29][23] ;
 wire \registers[29][24] ;
 wire \registers[29][25] ;
 wire \registers[29][26] ;
 wire \registers[29][27] ;
 wire \registers[29][28] ;
 wire \registers[29][29] ;
 wire \registers[29][2] ;
 wire \registers[29][30] ;
 wire \registers[29][31] ;
 wire \registers[29][3] ;
 wire \registers[29][4] ;
 wire \registers[29][5] ;
 wire \registers[29][6] ;
 wire \registers[29][7] ;
 wire \registers[29][8] ;
 wire \registers[29][9] ;
 wire \registers[2][0] ;
 wire \registers[2][10] ;
 wire \registers[2][11] ;
 wire \registers[2][12] ;
 wire \registers[2][13] ;
 wire \registers[2][14] ;
 wire \registers[2][15] ;
 wire \registers[2][16] ;
 wire \registers[2][17] ;
 wire \registers[2][18] ;
 wire \registers[2][19] ;
 wire \registers[2][1] ;
 wire \registers[2][20] ;
 wire \registers[2][21] ;
 wire \registers[2][22] ;
 wire \registers[2][23] ;
 wire \registers[2][24] ;
 wire \registers[2][25] ;
 wire \registers[2][26] ;
 wire \registers[2][27] ;
 wire \registers[2][28] ;
 wire \registers[2][29] ;
 wire \registers[2][2] ;
 wire \registers[2][30] ;
 wire \registers[2][31] ;
 wire \registers[2][3] ;
 wire \registers[2][4] ;
 wire \registers[2][5] ;
 wire \registers[2][6] ;
 wire \registers[2][7] ;
 wire \registers[2][8] ;
 wire \registers[2][9] ;
 wire \registers[30][0] ;
 wire \registers[30][10] ;
 wire \registers[30][11] ;
 wire \registers[30][12] ;
 wire \registers[30][13] ;
 wire \registers[30][14] ;
 wire \registers[30][15] ;
 wire \registers[30][16] ;
 wire \registers[30][17] ;
 wire \registers[30][18] ;
 wire \registers[30][19] ;
 wire \registers[30][1] ;
 wire \registers[30][20] ;
 wire \registers[30][21] ;
 wire \registers[30][22] ;
 wire \registers[30][23] ;
 wire \registers[30][24] ;
 wire \registers[30][25] ;
 wire \registers[30][26] ;
 wire \registers[30][27] ;
 wire \registers[30][28] ;
 wire \registers[30][29] ;
 wire \registers[30][2] ;
 wire \registers[30][30] ;
 wire \registers[30][31] ;
 wire \registers[30][3] ;
 wire \registers[30][4] ;
 wire \registers[30][5] ;
 wire \registers[30][6] ;
 wire \registers[30][7] ;
 wire \registers[30][8] ;
 wire \registers[30][9] ;
 wire \registers[31][0] ;
 wire \registers[31][10] ;
 wire \registers[31][11] ;
 wire \registers[31][12] ;
 wire \registers[31][13] ;
 wire \registers[31][14] ;
 wire \registers[31][15] ;
 wire \registers[31][16] ;
 wire \registers[31][17] ;
 wire \registers[31][18] ;
 wire \registers[31][19] ;
 wire \registers[31][1] ;
 wire \registers[31][20] ;
 wire \registers[31][21] ;
 wire \registers[31][22] ;
 wire \registers[31][23] ;
 wire \registers[31][24] ;
 wire \registers[31][25] ;
 wire \registers[31][26] ;
 wire \registers[31][27] ;
 wire \registers[31][28] ;
 wire \registers[31][29] ;
 wire \registers[31][2] ;
 wire \registers[31][30] ;
 wire \registers[31][31] ;
 wire \registers[31][3] ;
 wire \registers[31][4] ;
 wire \registers[31][5] ;
 wire \registers[31][6] ;
 wire \registers[31][7] ;
 wire \registers[31][8] ;
 wire \registers[31][9] ;
 wire \registers[3][0] ;
 wire \registers[3][10] ;
 wire \registers[3][11] ;
 wire \registers[3][12] ;
 wire \registers[3][13] ;
 wire \registers[3][14] ;
 wire \registers[3][15] ;
 wire \registers[3][16] ;
 wire \registers[3][17] ;
 wire \registers[3][18] ;
 wire \registers[3][19] ;
 wire \registers[3][1] ;
 wire \registers[3][20] ;
 wire \registers[3][21] ;
 wire \registers[3][22] ;
 wire \registers[3][23] ;
 wire \registers[3][24] ;
 wire \registers[3][25] ;
 wire \registers[3][26] ;
 wire \registers[3][27] ;
 wire \registers[3][28] ;
 wire \registers[3][29] ;
 wire \registers[3][2] ;
 wire \registers[3][30] ;
 wire \registers[3][31] ;
 wire \registers[3][3] ;
 wire \registers[3][4] ;
 wire \registers[3][5] ;
 wire \registers[3][6] ;
 wire \registers[3][7] ;
 wire \registers[3][8] ;
 wire \registers[3][9] ;
 wire \registers[4][0] ;
 wire \registers[4][10] ;
 wire \registers[4][11] ;
 wire \registers[4][12] ;
 wire \registers[4][13] ;
 wire \registers[4][14] ;
 wire \registers[4][15] ;
 wire \registers[4][16] ;
 wire \registers[4][17] ;
 wire \registers[4][18] ;
 wire \registers[4][19] ;
 wire \registers[4][1] ;
 wire \registers[4][20] ;
 wire \registers[4][21] ;
 wire \registers[4][22] ;
 wire \registers[4][23] ;
 wire \registers[4][24] ;
 wire \registers[4][25] ;
 wire \registers[4][26] ;
 wire \registers[4][27] ;
 wire \registers[4][28] ;
 wire \registers[4][29] ;
 wire \registers[4][2] ;
 wire \registers[4][30] ;
 wire \registers[4][31] ;
 wire \registers[4][3] ;
 wire \registers[4][4] ;
 wire \registers[4][5] ;
 wire \registers[4][6] ;
 wire \registers[4][7] ;
 wire \registers[4][8] ;
 wire \registers[4][9] ;
 wire \registers[5][0] ;
 wire \registers[5][10] ;
 wire \registers[5][11] ;
 wire \registers[5][12] ;
 wire \registers[5][13] ;
 wire \registers[5][14] ;
 wire \registers[5][15] ;
 wire \registers[5][16] ;
 wire \registers[5][17] ;
 wire \registers[5][18] ;
 wire \registers[5][19] ;
 wire \registers[5][1] ;
 wire \registers[5][20] ;
 wire \registers[5][21] ;
 wire \registers[5][22] ;
 wire \registers[5][23] ;
 wire \registers[5][24] ;
 wire \registers[5][25] ;
 wire \registers[5][26] ;
 wire \registers[5][27] ;
 wire \registers[5][28] ;
 wire \registers[5][29] ;
 wire \registers[5][2] ;
 wire \registers[5][30] ;
 wire \registers[5][31] ;
 wire \registers[5][3] ;
 wire \registers[5][4] ;
 wire \registers[5][5] ;
 wire \registers[5][6] ;
 wire \registers[5][7] ;
 wire \registers[5][8] ;
 wire \registers[5][9] ;
 wire \registers[6][0] ;
 wire \registers[6][10] ;
 wire \registers[6][11] ;
 wire \registers[6][12] ;
 wire \registers[6][13] ;
 wire \registers[6][14] ;
 wire \registers[6][15] ;
 wire \registers[6][16] ;
 wire \registers[6][17] ;
 wire \registers[6][18] ;
 wire \registers[6][19] ;
 wire \registers[6][1] ;
 wire \registers[6][20] ;
 wire \registers[6][21] ;
 wire \registers[6][22] ;
 wire \registers[6][23] ;
 wire \registers[6][24] ;
 wire \registers[6][25] ;
 wire \registers[6][26] ;
 wire \registers[6][27] ;
 wire \registers[6][28] ;
 wire \registers[6][29] ;
 wire \registers[6][2] ;
 wire \registers[6][30] ;
 wire \registers[6][31] ;
 wire \registers[6][3] ;
 wire \registers[6][4] ;
 wire \registers[6][5] ;
 wire \registers[6][6] ;
 wire \registers[6][7] ;
 wire \registers[6][8] ;
 wire \registers[6][9] ;
 wire \registers[7][0] ;
 wire \registers[7][10] ;
 wire \registers[7][11] ;
 wire \registers[7][12] ;
 wire \registers[7][13] ;
 wire \registers[7][14] ;
 wire \registers[7][15] ;
 wire \registers[7][16] ;
 wire \registers[7][17] ;
 wire \registers[7][18] ;
 wire \registers[7][19] ;
 wire \registers[7][1] ;
 wire \registers[7][20] ;
 wire \registers[7][21] ;
 wire \registers[7][22] ;
 wire \registers[7][23] ;
 wire \registers[7][24] ;
 wire \registers[7][25] ;
 wire \registers[7][26] ;
 wire \registers[7][27] ;
 wire \registers[7][28] ;
 wire \registers[7][29] ;
 wire \registers[7][2] ;
 wire \registers[7][30] ;
 wire \registers[7][31] ;
 wire \registers[7][3] ;
 wire \registers[7][4] ;
 wire \registers[7][5] ;
 wire \registers[7][6] ;
 wire \registers[7][7] ;
 wire \registers[7][8] ;
 wire \registers[7][9] ;
 wire \registers[8][0] ;
 wire \registers[8][10] ;
 wire \registers[8][11] ;
 wire \registers[8][12] ;
 wire \registers[8][13] ;
 wire \registers[8][14] ;
 wire \registers[8][15] ;
 wire \registers[8][16] ;
 wire \registers[8][17] ;
 wire \registers[8][18] ;
 wire \registers[8][19] ;
 wire \registers[8][1] ;
 wire \registers[8][20] ;
 wire \registers[8][21] ;
 wire \registers[8][22] ;
 wire \registers[8][23] ;
 wire \registers[8][24] ;
 wire \registers[8][25] ;
 wire \registers[8][26] ;
 wire \registers[8][27] ;
 wire \registers[8][28] ;
 wire \registers[8][29] ;
 wire \registers[8][2] ;
 wire \registers[8][30] ;
 wire \registers[8][31] ;
 wire \registers[8][3] ;
 wire \registers[8][4] ;
 wire \registers[8][5] ;
 wire \registers[8][6] ;
 wire \registers[8][7] ;
 wire \registers[8][8] ;
 wire \registers[8][9] ;
 wire \registers[9][0] ;
 wire \registers[9][10] ;
 wire \registers[9][11] ;
 wire \registers[9][12] ;
 wire \registers[9][13] ;
 wire \registers[9][14] ;
 wire \registers[9][15] ;
 wire \registers[9][16] ;
 wire \registers[9][17] ;
 wire \registers[9][18] ;
 wire \registers[9][19] ;
 wire \registers[9][1] ;
 wire \registers[9][20] ;
 wire \registers[9][21] ;
 wire \registers[9][22] ;
 wire \registers[9][23] ;
 wire \registers[9][24] ;
 wire \registers[9][25] ;
 wire \registers[9][26] ;
 wire \registers[9][27] ;
 wire \registers[9][28] ;
 wire \registers[9][29] ;
 wire \registers[9][2] ;
 wire \registers[9][30] ;
 wire \registers[9][31] ;
 wire \registers[9][3] ;
 wire \registers[9][4] ;
 wire \registers[9][5] ;
 wire \registers[9][6] ;
 wire \registers[9][7] ;
 wire \registers[9][8] ;
 wire \registers[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;

 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4178_ (.I(net39),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4179_ (.I(net9),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4180_ (.I(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4181_ (.I(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4182_ (.A1(_1091_),
    .A2(\registers[29][31] ),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _4183_ (.A1(net13),
    .A2(net14),
    .A3(net12),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _4184_ (.A1(net9),
    .A2(net10),
    .A3(net47),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _4185_ (.A1(net11),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4186_ (.A1(_1093_),
    .A2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4187_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4188_ (.I0(_1088_),
    .I1(_1092_),
    .S(_1097_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4189_ (.I(net40),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4190_ (.A1(_1091_),
    .A2(\registers[29][3] ),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4191_ (.I0(_1098_),
    .I1(_1099_),
    .S(_1097_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4192_ (.I(net41),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4193_ (.A1(_1091_),
    .A2(\registers[29][4] ),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4194_ (.I0(_1100_),
    .I1(_1101_),
    .S(_1097_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4195_ (.I(net42),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4196_ (.A1(_1091_),
    .A2(\registers[29][5] ),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4197_ (.I0(_1102_),
    .I1(_1103_),
    .S(_1097_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4198_ (.I(net43),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4199_ (.A1(_1091_),
    .A2(\registers[29][6] ),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4200_ (.I0(_1104_),
    .I1(_1105_),
    .S(_1097_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4201_ (.I(net44),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4202_ (.A1(_1091_),
    .A2(\registers[29][7] ),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4203_ (.I0(_1106_),
    .I1(_1107_),
    .S(_1097_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4204_ (.I(net45),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4205_ (.A1(_1091_),
    .A2(\registers[29][8] ),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4206_ (.I0(_1108_),
    .I1(_1109_),
    .S(_1097_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4207_ (.I(net46),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4208_ (.A1(_1091_),
    .A2(\registers[29][9] ),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4209_ (.I0(_1110_),
    .I1(_1111_),
    .S(_1097_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4210_ (.I(_1089_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4211_ (.I(_1112_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4212_ (.A1(_1113_),
    .A2(\registers[2][0] ),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4213_ (.I(net15),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _4214_ (.A1(net13),
    .A2(net14),
    .A3(net12),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _4215_ (.A1(net9),
    .A2(net47),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _4216_ (.A1(net10),
    .A2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4217_ (.A1(net11),
    .A2(_1118_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4218_ (.A1(_1116_),
    .A2(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4219_ (.I(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4220_ (.I0(_1114_),
    .I1(_1115_),
    .S(_1121_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4221_ (.A1(_1113_),
    .A2(\registers[2][10] ),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4222_ (.I(net16),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4223_ (.I0(_1122_),
    .I1(_1123_),
    .S(_1121_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4224_ (.A1(_1113_),
    .A2(\registers[2][11] ),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4225_ (.I(net17),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4226_ (.I0(_1124_),
    .I1(_1125_),
    .S(_1121_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4227_ (.A1(_1113_),
    .A2(\registers[2][12] ),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4228_ (.I(net18),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4229_ (.I0(_1126_),
    .I1(_1127_),
    .S(_1121_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4230_ (.A1(_1113_),
    .A2(\registers[2][13] ),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4231_ (.I(net19),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4232_ (.I0(_1128_),
    .I1(_1129_),
    .S(_1121_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4233_ (.A1(_1113_),
    .A2(\registers[2][14] ),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4234_ (.I(net20),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4235_ (.I0(_1130_),
    .I1(_1131_),
    .S(_1121_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4236_ (.A1(_1113_),
    .A2(\registers[2][15] ),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4237_ (.I(net21),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4238_ (.I0(_1132_),
    .I1(_1133_),
    .S(_1121_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4239_ (.A1(_1113_),
    .A2(\registers[2][16] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4240_ (.I(net22),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4241_ (.I0(_1134_),
    .I1(_1135_),
    .S(_1121_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4242_ (.A1(_1113_),
    .A2(\registers[2][17] ),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4243_ (.I(net23),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4244_ (.I0(_1136_),
    .I1(_1137_),
    .S(_1121_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4245_ (.A1(_1113_),
    .A2(\registers[2][18] ),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4246_ (.I(net24),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4247_ (.I0(_1138_),
    .I1(_1139_),
    .S(_1121_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4248_ (.I(_1112_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4249_ (.A1(_1140_),
    .A2(\registers[2][19] ),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4250_ (.I(net25),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4251_ (.I(_1120_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4252_ (.I0(_1141_),
    .I1(_1142_),
    .S(_1143_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4253_ (.A1(_1140_),
    .A2(\registers[2][1] ),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4254_ (.I(net26),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4255_ (.I0(_1144_),
    .I1(_1145_),
    .S(_1143_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4256_ (.A1(_1140_),
    .A2(\registers[2][20] ),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4257_ (.I(net27),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4258_ (.I0(_1146_),
    .I1(_1147_),
    .S(_1143_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4259_ (.A1(_1140_),
    .A2(\registers[2][21] ),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4260_ (.I(net28),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4261_ (.I0(_1148_),
    .I1(_1149_),
    .S(_1143_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4262_ (.A1(_1140_),
    .A2(\registers[2][22] ),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4263_ (.I(net29),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4264_ (.I0(_1150_),
    .I1(_1151_),
    .S(_1143_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4265_ (.A1(_1140_),
    .A2(\registers[2][23] ),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4266_ (.I(net30),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4267_ (.I0(_1152_),
    .I1(_1153_),
    .S(_1143_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4268_ (.A1(_1140_),
    .A2(\registers[2][24] ),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4269_ (.I(net31),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4270_ (.I0(_1154_),
    .I1(_1155_),
    .S(_1143_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4271_ (.A1(_1140_),
    .A2(\registers[2][25] ),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4272_ (.I(net32),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4273_ (.I0(_1156_),
    .I1(_1157_),
    .S(_1143_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4274_ (.A1(_1140_),
    .A2(\registers[2][26] ),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4275_ (.I(net33),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4276_ (.I0(_1158_),
    .I1(_1159_),
    .S(_1143_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4277_ (.A1(_1140_),
    .A2(\registers[2][27] ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4278_ (.I(net34),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4279_ (.I0(_1160_),
    .I1(_1161_),
    .S(_1143_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4280_ (.I(_1112_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4281_ (.A1(_1162_),
    .A2(\registers[2][28] ),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4282_ (.I(net35),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4283_ (.I(_1120_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4284_ (.I0(_1163_),
    .I1(_1164_),
    .S(_1165_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4285_ (.A1(_1162_),
    .A2(\registers[2][29] ),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4286_ (.I(net36),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4287_ (.I0(_1166_),
    .I1(_1167_),
    .S(_1165_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4288_ (.A1(_1162_),
    .A2(\registers[2][2] ),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4289_ (.I(net37),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4290_ (.I0(_1168_),
    .I1(_1169_),
    .S(_1165_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4291_ (.A1(_1162_),
    .A2(\registers[2][30] ),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4292_ (.I(net38),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4293_ (.I0(_1170_),
    .I1(_1171_),
    .S(_1165_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4294_ (.A1(_1162_),
    .A2(\registers[2][31] ),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4295_ (.I(net39),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4296_ (.I0(_1172_),
    .I1(_1173_),
    .S(_1165_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4297_ (.A1(_1162_),
    .A2(\registers[2][3] ),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4298_ (.I(net40),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4299_ (.I0(_1174_),
    .I1(_1175_),
    .S(_1165_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4300_ (.A1(_1162_),
    .A2(\registers[2][4] ),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4301_ (.I(net41),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4302_ (.I0(_1176_),
    .I1(_1177_),
    .S(_1165_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4303_ (.A1(_1162_),
    .A2(\registers[2][5] ),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4304_ (.I(net42),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4305_ (.I0(_1178_),
    .I1(_1179_),
    .S(_1165_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4306_ (.A1(_1162_),
    .A2(\registers[2][6] ),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4307_ (.I(net43),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4308_ (.I0(_1180_),
    .I1(_1181_),
    .S(_1165_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4309_ (.A1(_1162_),
    .A2(\registers[2][7] ),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4310_ (.I(net44),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4311_ (.I0(_1182_),
    .I1(_1183_),
    .S(_1165_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4312_ (.I(_1112_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4313_ (.A1(_1184_),
    .A2(\registers[2][8] ),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4314_ (.I(net45),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4315_ (.I0(_1185_),
    .I1(_1186_),
    .S(_1120_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4316_ (.A1(_1184_),
    .A2(\registers[2][9] ),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4317_ (.I(net46),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4318_ (.I0(_1187_),
    .I1(_1188_),
    .S(_1120_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4319_ (.A1(_1184_),
    .A2(\registers[30][0] ),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4320_ (.A1(_1093_),
    .A2(_1119_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4321_ (.I(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4322_ (.I0(_1189_),
    .I1(_1115_),
    .S(_1191_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4323_ (.A1(_1184_),
    .A2(\registers[30][10] ),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4324_ (.I0(_1192_),
    .I1(_1123_),
    .S(_1191_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4325_ (.A1(_1184_),
    .A2(\registers[30][11] ),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4326_ (.I0(_1193_),
    .I1(_1125_),
    .S(_1191_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4327_ (.A1(_1184_),
    .A2(\registers[30][12] ),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4328_ (.I0(_1194_),
    .I1(_1127_),
    .S(_1191_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4329_ (.A1(_1184_),
    .A2(\registers[30][13] ),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4330_ (.I0(_1195_),
    .I1(_1129_),
    .S(_1191_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4331_ (.A1(_1184_),
    .A2(\registers[30][14] ),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4332_ (.I0(_1196_),
    .I1(_1131_),
    .S(_1191_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4333_ (.A1(_1184_),
    .A2(\registers[30][15] ),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4334_ (.I0(_1197_),
    .I1(_1133_),
    .S(_1191_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4335_ (.A1(_1184_),
    .A2(\registers[30][16] ),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4336_ (.I0(_1198_),
    .I1(_1135_),
    .S(_1191_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4337_ (.I(_1112_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4338_ (.A1(_1199_),
    .A2(\registers[30][17] ),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4339_ (.I0(_1200_),
    .I1(_1137_),
    .S(_1191_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4340_ (.A1(_1199_),
    .A2(\registers[30][18] ),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4341_ (.I0(_1201_),
    .I1(_1139_),
    .S(_1191_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4342_ (.A1(_1199_),
    .A2(\registers[30][19] ),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4343_ (.I(_1190_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4344_ (.I0(_1202_),
    .I1(_1142_),
    .S(_1203_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4345_ (.A1(_1199_),
    .A2(\registers[30][1] ),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4346_ (.I0(_1204_),
    .I1(_1145_),
    .S(_1203_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4347_ (.A1(_1199_),
    .A2(\registers[30][20] ),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4348_ (.I0(_1205_),
    .I1(_1147_),
    .S(_1203_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4349_ (.A1(_1199_),
    .A2(\registers[30][21] ),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4350_ (.I0(_1206_),
    .I1(_1149_),
    .S(_1203_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4351_ (.A1(_1199_),
    .A2(\registers[30][22] ),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4352_ (.I0(_1207_),
    .I1(_1151_),
    .S(_1203_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4353_ (.A1(_1199_),
    .A2(\registers[30][23] ),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4354_ (.I0(_1208_),
    .I1(_1153_),
    .S(_1203_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4355_ (.A1(_1199_),
    .A2(\registers[30][24] ),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4356_ (.I0(_1209_),
    .I1(_1155_),
    .S(_1203_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4357_ (.A1(_1199_),
    .A2(\registers[30][25] ),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4358_ (.I0(_1210_),
    .I1(_1157_),
    .S(_1203_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4359_ (.I(_1112_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4360_ (.A1(_1211_),
    .A2(\registers[30][26] ),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4361_ (.I0(_1212_),
    .I1(_1159_),
    .S(_1203_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4362_ (.A1(_1211_),
    .A2(\registers[30][27] ),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4363_ (.I0(_1213_),
    .I1(_1161_),
    .S(_1203_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4364_ (.A1(_1211_),
    .A2(\registers[30][28] ),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4365_ (.I(_1190_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4366_ (.I0(_1214_),
    .I1(_1164_),
    .S(_1215_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4367_ (.A1(_1211_),
    .A2(\registers[30][29] ),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4368_ (.I0(_1216_),
    .I1(_1167_),
    .S(_1215_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4369_ (.A1(_1211_),
    .A2(\registers[30][2] ),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4370_ (.I0(_1217_),
    .I1(_1169_),
    .S(_1215_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4371_ (.A1(_1211_),
    .A2(\registers[30][30] ),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4372_ (.I0(_1218_),
    .I1(_1171_),
    .S(_1215_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4373_ (.A1(_1211_),
    .A2(\registers[30][31] ),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4374_ (.I0(_1219_),
    .I1(_1173_),
    .S(_1215_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4375_ (.A1(_1211_),
    .A2(\registers[30][3] ),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4376_ (.I0(_1220_),
    .I1(_1175_),
    .S(_1215_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4377_ (.A1(_1211_),
    .A2(\registers[30][4] ),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4378_ (.I0(_1221_),
    .I1(_1177_),
    .S(_1215_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4379_ (.A1(_1211_),
    .A2(\registers[30][5] ),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4380_ (.I0(_1222_),
    .I1(_1179_),
    .S(_1215_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4381_ (.I(_1089_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4382_ (.I(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4383_ (.A1(_1224_),
    .A2(\registers[30][6] ),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4384_ (.I0(_1225_),
    .I1(_1181_),
    .S(_1215_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4385_ (.A1(_1224_),
    .A2(\registers[30][7] ),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4386_ (.I0(_1226_),
    .I1(_1183_),
    .S(_1215_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4387_ (.A1(_1224_),
    .A2(\registers[30][8] ),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4388_ (.I0(_1227_),
    .I1(_1186_),
    .S(_1190_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4389_ (.A1(_1224_),
    .A2(\registers[30][9] ),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4390_ (.I0(_1228_),
    .I1(_1188_),
    .S(_1190_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4391_ (.I(net15),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4392_ (.I(_1090_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4393_ (.A1(_1230_),
    .A2(\registers[31][0] ),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _4394_ (.A1(net9),
    .A2(net10),
    .A3(net11),
    .A4(net47),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4395_ (.A1(_1093_),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4396_ (.I(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4397_ (.I0(_1229_),
    .I1(_1231_),
    .S(_1234_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4398_ (.I(net16),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4399_ (.A1(_1230_),
    .A2(\registers[31][10] ),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4400_ (.I0(_1235_),
    .I1(_1236_),
    .S(_1234_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4401_ (.I(net17),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4402_ (.A1(_1230_),
    .A2(\registers[31][11] ),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4403_ (.I0(_1237_),
    .I1(_1238_),
    .S(_1234_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4404_ (.I(net18),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4405_ (.A1(_1230_),
    .A2(\registers[31][12] ),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4406_ (.I0(_1239_),
    .I1(_1240_),
    .S(_1234_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4407_ (.I(net19),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4408_ (.A1(_1230_),
    .A2(\registers[31][13] ),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4409_ (.I0(_1241_),
    .I1(_1242_),
    .S(_1234_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4410_ (.I(net20),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4411_ (.A1(_1230_),
    .A2(\registers[31][14] ),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4412_ (.I0(_1243_),
    .I1(_1244_),
    .S(_1234_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4413_ (.I(net21),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4414_ (.A1(_1230_),
    .A2(\registers[31][15] ),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4415_ (.I0(_1245_),
    .I1(_1246_),
    .S(_1234_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4416_ (.I(net22),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4417_ (.A1(_1230_),
    .A2(\registers[31][16] ),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4418_ (.I0(_1247_),
    .I1(_1248_),
    .S(_1234_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4419_ (.I(net23),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4420_ (.A1(_1230_),
    .A2(\registers[31][17] ),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4421_ (.I0(_1249_),
    .I1(_1250_),
    .S(_1234_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4422_ (.I(net24),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4423_ (.A1(_1230_),
    .A2(\registers[31][18] ),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4424_ (.I0(_1251_),
    .I1(_1252_),
    .S(_1234_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4425_ (.I(net25),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4426_ (.I(_1090_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4427_ (.A1(_1254_),
    .A2(\registers[31][19] ),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4428_ (.I(_1233_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4429_ (.I0(_1253_),
    .I1(_1255_),
    .S(_1256_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4430_ (.I(net26),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4431_ (.A1(_1254_),
    .A2(\registers[31][1] ),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4432_ (.I0(_1257_),
    .I1(_1258_),
    .S(_1256_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4433_ (.I(net27),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4434_ (.A1(_1254_),
    .A2(\registers[31][20] ),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4435_ (.I0(_1259_),
    .I1(_1260_),
    .S(_1256_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4436_ (.I(net28),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4437_ (.A1(_1254_),
    .A2(\registers[31][21] ),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4438_ (.I0(_1261_),
    .I1(_1262_),
    .S(_1256_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4439_ (.I(net29),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4440_ (.A1(_1254_),
    .A2(\registers[31][22] ),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4441_ (.I0(_1263_),
    .I1(_1264_),
    .S(_1256_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4442_ (.I(net30),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4443_ (.A1(_1254_),
    .A2(\registers[31][23] ),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4444_ (.I0(_1265_),
    .I1(_1266_),
    .S(_1256_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4445_ (.I(net31),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4446_ (.A1(_1254_),
    .A2(\registers[31][24] ),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4447_ (.I0(_1267_),
    .I1(_1268_),
    .S(_1256_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4448_ (.I(net32),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4449_ (.A1(_1254_),
    .A2(\registers[31][25] ),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4450_ (.I0(_1269_),
    .I1(_1270_),
    .S(_1256_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4451_ (.I(net33),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4452_ (.A1(_1254_),
    .A2(\registers[31][26] ),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4453_ (.I0(_1271_),
    .I1(_1272_),
    .S(_1256_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4454_ (.I(net34),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4455_ (.A1(_1254_),
    .A2(\registers[31][27] ),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4456_ (.I0(_1273_),
    .I1(_1274_),
    .S(_1256_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4457_ (.I(net35),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4458_ (.I(_1090_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4459_ (.A1(_1276_),
    .A2(\registers[31][28] ),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4460_ (.I(_1233_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4461_ (.I0(_1275_),
    .I1(_1277_),
    .S(_1278_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4462_ (.I(net36),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4463_ (.A1(_1276_),
    .A2(\registers[31][29] ),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4464_ (.I0(_1279_),
    .I1(_1280_),
    .S(_1278_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4465_ (.I(net37),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4466_ (.A1(_1276_),
    .A2(\registers[31][2] ),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4467_ (.I0(_1281_),
    .I1(_1282_),
    .S(_1278_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4468_ (.I(net38),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4469_ (.A1(_1276_),
    .A2(\registers[31][30] ),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4470_ (.I0(_1283_),
    .I1(_1284_),
    .S(_1278_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4471_ (.A1(_1276_),
    .A2(\registers[31][31] ),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4472_ (.I0(_1088_),
    .I1(_1285_),
    .S(_1278_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4473_ (.A1(_1276_),
    .A2(\registers[31][3] ),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4474_ (.I0(_1098_),
    .I1(_1286_),
    .S(_1278_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4475_ (.A1(_1276_),
    .A2(\registers[31][4] ),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4476_ (.I0(_1100_),
    .I1(_1287_),
    .S(_1278_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4477_ (.A1(_1276_),
    .A2(\registers[31][5] ),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4478_ (.I0(_1102_),
    .I1(_1288_),
    .S(_1278_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4479_ (.A1(_1276_),
    .A2(\registers[31][6] ),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4480_ (.I0(_1104_),
    .I1(_1289_),
    .S(_1278_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4481_ (.A1(_1276_),
    .A2(\registers[31][7] ),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4482_ (.I0(_1106_),
    .I1(_1290_),
    .S(_1278_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4483_ (.I(_1090_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4484_ (.A1(_1291_),
    .A2(\registers[31][8] ),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4485_ (.I0(_1108_),
    .I1(_1292_),
    .S(_1233_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4486_ (.A1(_1291_),
    .A2(\registers[31][9] ),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4487_ (.I0(_1110_),
    .I1(_1293_),
    .S(_1233_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4488_ (.A1(_1291_),
    .A2(\registers[3][0] ),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4489_ (.A1(_1116_),
    .A2(_1232_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4490_ (.I(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4491_ (.I0(_1229_),
    .I1(_1294_),
    .S(_1296_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4492_ (.A1(_1291_),
    .A2(\registers[3][10] ),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4493_ (.I0(_1235_),
    .I1(_1297_),
    .S(_1296_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4494_ (.A1(_1291_),
    .A2(\registers[3][11] ),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4495_ (.I0(_1237_),
    .I1(_1298_),
    .S(_1296_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4496_ (.A1(_1291_),
    .A2(\registers[3][12] ),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4497_ (.I0(_1239_),
    .I1(_1299_),
    .S(_1296_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4498_ (.A1(_1291_),
    .A2(\registers[3][13] ),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4499_ (.I0(_1241_),
    .I1(_1300_),
    .S(_1296_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4500_ (.A1(_1291_),
    .A2(\registers[3][14] ),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4501_ (.I0(_1243_),
    .I1(_1301_),
    .S(_1296_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4502_ (.A1(_1291_),
    .A2(\registers[3][15] ),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4503_ (.I0(_1245_),
    .I1(_1302_),
    .S(_1296_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4504_ (.A1(_1291_),
    .A2(\registers[3][16] ),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4505_ (.I0(_1247_),
    .I1(_1303_),
    .S(_1296_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4506_ (.I(_1090_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4507_ (.A1(_1304_),
    .A2(\registers[3][17] ),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4508_ (.I0(_1249_),
    .I1(_1305_),
    .S(_1296_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4509_ (.A1(_1304_),
    .A2(\registers[3][18] ),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4510_ (.I0(_1251_),
    .I1(_1306_),
    .S(_1296_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4511_ (.A1(_1304_),
    .A2(\registers[3][19] ),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4512_ (.I(_1295_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4513_ (.I0(_1253_),
    .I1(_1307_),
    .S(_1308_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4514_ (.A1(_1304_),
    .A2(\registers[3][1] ),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4515_ (.I0(_1257_),
    .I1(_1309_),
    .S(_1308_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4516_ (.A1(_1304_),
    .A2(\registers[3][20] ),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4517_ (.I0(_1259_),
    .I1(_1310_),
    .S(_1308_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4518_ (.A1(_1304_),
    .A2(\registers[3][21] ),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4519_ (.I0(_1261_),
    .I1(_1311_),
    .S(_1308_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4520_ (.A1(_1304_),
    .A2(\registers[3][22] ),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4521_ (.I0(_1263_),
    .I1(_1312_),
    .S(_1308_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4522_ (.A1(_1304_),
    .A2(\registers[3][23] ),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4523_ (.I0(_1265_),
    .I1(_1313_),
    .S(_1308_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4524_ (.A1(_1304_),
    .A2(\registers[3][24] ),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4525_ (.I0(_1267_),
    .I1(_1314_),
    .S(_1308_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4526_ (.A1(_1304_),
    .A2(\registers[3][25] ),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4527_ (.I0(_1269_),
    .I1(_1315_),
    .S(_1308_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4528_ (.I(_1090_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4529_ (.A1(_1316_),
    .A2(\registers[3][26] ),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4530_ (.I0(_1271_),
    .I1(_1317_),
    .S(_1308_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4531_ (.A1(_1316_),
    .A2(\registers[3][27] ),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4532_ (.I0(_1273_),
    .I1(_1318_),
    .S(_1308_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4533_ (.A1(_1316_),
    .A2(\registers[3][28] ),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4534_ (.I(_1295_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4535_ (.I0(_1275_),
    .I1(_1319_),
    .S(_1320_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4536_ (.A1(_1316_),
    .A2(\registers[3][29] ),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4537_ (.I0(_1279_),
    .I1(_1321_),
    .S(_1320_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4538_ (.A1(_1316_),
    .A2(\registers[3][2] ),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4539_ (.I0(_1281_),
    .I1(_1322_),
    .S(_1320_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4540_ (.A1(_1316_),
    .A2(\registers[3][30] ),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4541_ (.I0(_1283_),
    .I1(_1323_),
    .S(_1320_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4542_ (.A1(_1316_),
    .A2(\registers[3][31] ),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4543_ (.I0(_1088_),
    .I1(_1324_),
    .S(_1320_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4544_ (.A1(_1316_),
    .A2(\registers[3][3] ),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4545_ (.I0(_1098_),
    .I1(_1325_),
    .S(_1320_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4546_ (.A1(_1316_),
    .A2(\registers[3][4] ),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4547_ (.I0(_1100_),
    .I1(_1326_),
    .S(_1320_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4548_ (.A1(_1316_),
    .A2(\registers[3][5] ),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4549_ (.I0(_1102_),
    .I1(_1327_),
    .S(_1320_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4550_ (.I(_1089_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4551_ (.I(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4552_ (.A1(_1329_),
    .A2(\registers[3][6] ),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4553_ (.I0(_1104_),
    .I1(_1330_),
    .S(_1320_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4554_ (.A1(_1329_),
    .A2(\registers[3][7] ),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4555_ (.I0(_1106_),
    .I1(_1331_),
    .S(_1320_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4556_ (.A1(_1329_),
    .A2(\registers[3][8] ),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4557_ (.I0(_1108_),
    .I1(_1332_),
    .S(_1295_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4558_ (.A1(_1329_),
    .A2(\registers[3][9] ),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4559_ (.I0(_1110_),
    .I1(_1333_),
    .S(_1295_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4560_ (.A1(_1329_),
    .A2(\registers[4][0] ),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _4561_ (.I(net12),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _4562_ (.A1(net13),
    .A2(net14),
    .A3(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _4563_ (.I(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _4564_ (.A1(net10),
    .A2(net11),
    .A3(_1117_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4565_ (.A1(_1337_),
    .A2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4566_ (.I(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4567_ (.I0(_1229_),
    .I1(_1334_),
    .S(_1340_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4568_ (.A1(_1329_),
    .A2(\registers[4][10] ),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4569_ (.I0(_1235_),
    .I1(_1341_),
    .S(_1340_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4570_ (.A1(_1329_),
    .A2(\registers[4][11] ),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4571_ (.I0(_1237_),
    .I1(_1342_),
    .S(_1340_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4572_ (.A1(_1329_),
    .A2(\registers[4][12] ),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4573_ (.I0(_1239_),
    .I1(_1343_),
    .S(_1340_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4574_ (.A1(_1329_),
    .A2(\registers[4][13] ),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4575_ (.I0(_1241_),
    .I1(_1344_),
    .S(_1340_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4576_ (.A1(_1329_),
    .A2(\registers[4][14] ),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4577_ (.I0(_1243_),
    .I1(_1345_),
    .S(_1340_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4578_ (.I(_1328_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4579_ (.A1(_1346_),
    .A2(\registers[4][15] ),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4580_ (.I0(_1245_),
    .I1(_1347_),
    .S(_1340_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4581_ (.A1(_1346_),
    .A2(\registers[4][16] ),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4582_ (.I0(_1247_),
    .I1(_1348_),
    .S(_1340_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4583_ (.A1(_1346_),
    .A2(\registers[4][17] ),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4584_ (.I0(_1249_),
    .I1(_1349_),
    .S(_1340_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4585_ (.A1(_1346_),
    .A2(\registers[4][18] ),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4586_ (.I0(_1251_),
    .I1(_1350_),
    .S(_1340_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4587_ (.A1(_1346_),
    .A2(\registers[4][19] ),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4588_ (.I(_1339_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4589_ (.I0(_1253_),
    .I1(_1351_),
    .S(_1352_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4590_ (.A1(_1346_),
    .A2(\registers[4][1] ),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4591_ (.I0(_1257_),
    .I1(_1353_),
    .S(_1352_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4592_ (.A1(_1346_),
    .A2(\registers[4][20] ),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4593_ (.I0(_1259_),
    .I1(_1354_),
    .S(_1352_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4594_ (.A1(_1346_),
    .A2(\registers[4][21] ),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4595_ (.I0(_1261_),
    .I1(_1355_),
    .S(_1352_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4596_ (.A1(_1346_),
    .A2(\registers[4][22] ),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4597_ (.I0(_1263_),
    .I1(_1356_),
    .S(_1352_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4598_ (.A1(_1346_),
    .A2(\registers[4][23] ),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4599_ (.I0(_1265_),
    .I1(_1357_),
    .S(_1352_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4600_ (.I(_1328_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4601_ (.A1(_1358_),
    .A2(\registers[4][24] ),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4602_ (.I0(_1267_),
    .I1(_1359_),
    .S(_1352_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4603_ (.A1(_1358_),
    .A2(\registers[4][25] ),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4604_ (.I0(_1269_),
    .I1(_1360_),
    .S(_1352_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4605_ (.A1(_1358_),
    .A2(\registers[4][26] ),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4606_ (.I0(_1271_),
    .I1(_1361_),
    .S(_1352_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4607_ (.A1(_1358_),
    .A2(\registers[4][27] ),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4608_ (.I0(_1273_),
    .I1(_1362_),
    .S(_1352_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4609_ (.A1(_1358_),
    .A2(\registers[4][28] ),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4610_ (.I(_1339_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4611_ (.I0(_1275_),
    .I1(_1363_),
    .S(_1364_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4612_ (.A1(_1358_),
    .A2(\registers[4][29] ),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4613_ (.I0(_1279_),
    .I1(_1365_),
    .S(_1364_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4614_ (.A1(_1358_),
    .A2(\registers[4][2] ),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4615_ (.I0(_1281_),
    .I1(_1366_),
    .S(_1364_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4616_ (.A1(_1358_),
    .A2(\registers[4][30] ),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4617_ (.I0(_1283_),
    .I1(_1367_),
    .S(_1364_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4618_ (.A1(_1358_),
    .A2(\registers[4][31] ),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4619_ (.I0(_1088_),
    .I1(_1368_),
    .S(_1364_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4620_ (.A1(_1358_),
    .A2(\registers[4][3] ),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4621_ (.I0(_1098_),
    .I1(_1369_),
    .S(_1364_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4622_ (.I(_1328_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4623_ (.A1(_1370_),
    .A2(\registers[4][4] ),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4624_ (.I0(_1100_),
    .I1(_1371_),
    .S(_1364_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4625_ (.A1(_1370_),
    .A2(\registers[4][5] ),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4626_ (.I0(_1102_),
    .I1(_1372_),
    .S(_1364_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4627_ (.A1(_1370_),
    .A2(\registers[4][6] ),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4628_ (.I0(_1104_),
    .I1(_1373_),
    .S(_1364_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4629_ (.A1(_1370_),
    .A2(\registers[4][7] ),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4630_ (.I0(_1106_),
    .I1(_1374_),
    .S(_1364_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4631_ (.A1(_1370_),
    .A2(\registers[4][8] ),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4632_ (.I0(_1108_),
    .I1(_1375_),
    .S(_1339_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4633_ (.A1(_1370_),
    .A2(\registers[4][9] ),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4634_ (.I0(_1110_),
    .I1(_1376_),
    .S(_1339_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4635_ (.A1(_1370_),
    .A2(\registers[5][0] ),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4636_ (.A1(_1095_),
    .A2(_1337_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4637_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4638_ (.I0(_1229_),
    .I1(_1377_),
    .S(_1379_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4639_ (.A1(_1370_),
    .A2(\registers[5][10] ),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4640_ (.I0(_1235_),
    .I1(_1380_),
    .S(_1379_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4641_ (.A1(_1370_),
    .A2(\registers[5][11] ),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4642_ (.I0(_1237_),
    .I1(_1381_),
    .S(_1379_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4643_ (.A1(_1370_),
    .A2(\registers[5][12] ),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4644_ (.I0(_1239_),
    .I1(_1382_),
    .S(_1379_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4645_ (.I(_1328_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4646_ (.A1(_1383_),
    .A2(\registers[5][13] ),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4647_ (.I0(_1241_),
    .I1(_1384_),
    .S(_1379_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4648_ (.A1(_1383_),
    .A2(\registers[5][14] ),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4649_ (.I0(_1243_),
    .I1(_1385_),
    .S(_1379_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4650_ (.A1(_1383_),
    .A2(\registers[5][15] ),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4651_ (.I0(_1245_),
    .I1(_1386_),
    .S(_1379_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4652_ (.A1(_1383_),
    .A2(\registers[5][16] ),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4653_ (.I0(_1247_),
    .I1(_1387_),
    .S(_1379_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4654_ (.A1(_1383_),
    .A2(\registers[5][17] ),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4655_ (.I0(_1249_),
    .I1(_1388_),
    .S(_1379_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4656_ (.A1(_1383_),
    .A2(\registers[5][18] ),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4657_ (.I0(_1251_),
    .I1(_1389_),
    .S(_1379_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4658_ (.A1(_1383_),
    .A2(\registers[5][19] ),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4659_ (.I(_1378_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4660_ (.I0(_1253_),
    .I1(_1390_),
    .S(_1391_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4661_ (.A1(_1383_),
    .A2(\registers[5][1] ),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4662_ (.I0(_1257_),
    .I1(_1392_),
    .S(_1391_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4663_ (.A1(_1383_),
    .A2(\registers[5][20] ),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4664_ (.I0(_1259_),
    .I1(_1393_),
    .S(_1391_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4665_ (.A1(_1383_),
    .A2(\registers[5][21] ),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4666_ (.I0(_1261_),
    .I1(_1394_),
    .S(_1391_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4667_ (.I(_1328_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4668_ (.A1(_1395_),
    .A2(\registers[5][22] ),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4669_ (.I0(_1263_),
    .I1(_1396_),
    .S(_1391_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4670_ (.A1(_1395_),
    .A2(\registers[5][23] ),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4671_ (.I0(_1265_),
    .I1(_1397_),
    .S(_1391_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4672_ (.A1(_1395_),
    .A2(\registers[5][24] ),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4673_ (.I0(_1267_),
    .I1(_1398_),
    .S(_1391_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4674_ (.A1(_1395_),
    .A2(\registers[5][25] ),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4675_ (.I0(_1269_),
    .I1(_1399_),
    .S(_1391_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4676_ (.A1(_1395_),
    .A2(\registers[5][26] ),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4677_ (.I0(_1271_),
    .I1(_1400_),
    .S(_1391_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4678_ (.A1(_1395_),
    .A2(\registers[5][27] ),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4679_ (.I0(_1273_),
    .I1(_1401_),
    .S(_1391_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4680_ (.A1(_1395_),
    .A2(\registers[5][28] ),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4681_ (.I(_1378_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4682_ (.I0(_1275_),
    .I1(_1402_),
    .S(_1403_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4683_ (.A1(_1395_),
    .A2(\registers[5][29] ),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4684_ (.I0(_1279_),
    .I1(_1404_),
    .S(_1403_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4685_ (.A1(_1395_),
    .A2(\registers[5][2] ),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4686_ (.I0(_1281_),
    .I1(_1405_),
    .S(_1403_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4687_ (.A1(_1395_),
    .A2(\registers[5][30] ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4688_ (.I0(_1283_),
    .I1(_1406_),
    .S(_1403_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4689_ (.I(_1328_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4690_ (.A1(_1407_),
    .A2(\registers[5][31] ),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4691_ (.I0(_1088_),
    .I1(_1408_),
    .S(_1403_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4692_ (.A1(_1407_),
    .A2(\registers[5][3] ),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4693_ (.I0(_1098_),
    .I1(_1409_),
    .S(_1403_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4694_ (.A1(_1407_),
    .A2(\registers[5][4] ),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4695_ (.I0(_1100_),
    .I1(_1410_),
    .S(_1403_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4696_ (.A1(_1407_),
    .A2(\registers[5][5] ),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4697_ (.I0(_1102_),
    .I1(_1411_),
    .S(_1403_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4698_ (.A1(_1407_),
    .A2(\registers[5][6] ),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4699_ (.I0(_1104_),
    .I1(_1412_),
    .S(_1403_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4700_ (.A1(_1407_),
    .A2(\registers[5][7] ),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4701_ (.I0(_1106_),
    .I1(_1413_),
    .S(_1403_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4702_ (.A1(_1407_),
    .A2(\registers[5][8] ),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4703_ (.I0(_1108_),
    .I1(_1414_),
    .S(_1378_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4704_ (.A1(_1407_),
    .A2(\registers[5][9] ),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4705_ (.I0(_1110_),
    .I1(_1415_),
    .S(_1378_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4706_ (.A1(_1407_),
    .A2(\registers[6][0] ),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4707_ (.A1(_1119_),
    .A2(_1337_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4708_ (.I(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4709_ (.I0(_1229_),
    .I1(_1416_),
    .S(_1418_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4710_ (.A1(_1407_),
    .A2(\registers[6][10] ),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4711_ (.I0(_1235_),
    .I1(_1419_),
    .S(_1418_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4712_ (.I(_1328_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4713_ (.A1(_1420_),
    .A2(\registers[6][11] ),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4714_ (.I0(_1237_),
    .I1(_1421_),
    .S(_1418_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4715_ (.A1(_1420_),
    .A2(\registers[6][12] ),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4716_ (.I0(_1239_),
    .I1(_1422_),
    .S(_1418_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4717_ (.A1(_1420_),
    .A2(\registers[6][13] ),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4718_ (.I0(_1241_),
    .I1(_1423_),
    .S(_1418_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4719_ (.A1(_1420_),
    .A2(\registers[6][14] ),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4720_ (.I0(_1243_),
    .I1(_1424_),
    .S(_1418_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4721_ (.A1(_1420_),
    .A2(\registers[6][15] ),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4722_ (.I0(_1245_),
    .I1(_1425_),
    .S(_1418_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4723_ (.A1(_1420_),
    .A2(\registers[6][16] ),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4724_ (.I0(_1247_),
    .I1(_1426_),
    .S(_1418_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4725_ (.A1(_1420_),
    .A2(\registers[6][17] ),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4726_ (.I0(_1249_),
    .I1(_1427_),
    .S(_1418_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4727_ (.A1(_1420_),
    .A2(\registers[6][18] ),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4728_ (.I0(_1251_),
    .I1(_1428_),
    .S(_1418_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4729_ (.A1(_1420_),
    .A2(\registers[6][19] ),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4730_ (.I(_1417_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4731_ (.I0(_1253_),
    .I1(_1429_),
    .S(_1430_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4732_ (.A1(_1420_),
    .A2(\registers[6][1] ),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4733_ (.I0(_1257_),
    .I1(_1431_),
    .S(_1430_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4734_ (.I(_1328_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4735_ (.A1(_1432_),
    .A2(\registers[6][20] ),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4736_ (.I0(_1259_),
    .I1(_1433_),
    .S(_1430_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4737_ (.A1(_1432_),
    .A2(\registers[6][21] ),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4738_ (.I0(_1261_),
    .I1(_1434_),
    .S(_1430_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4739_ (.A1(_1432_),
    .A2(\registers[6][22] ),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4740_ (.I0(_1263_),
    .I1(_1435_),
    .S(_1430_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4741_ (.A1(_1432_),
    .A2(\registers[6][23] ),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4742_ (.I0(_1265_),
    .I1(_1436_),
    .S(_1430_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4743_ (.A1(_1432_),
    .A2(\registers[6][24] ),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4744_ (.I0(_1267_),
    .I1(_1437_),
    .S(_1430_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4745_ (.A1(_1432_),
    .A2(\registers[6][25] ),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4746_ (.I0(_1269_),
    .I1(_1438_),
    .S(_1430_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4747_ (.A1(_1432_),
    .A2(\registers[6][26] ),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4748_ (.I0(_1271_),
    .I1(_1439_),
    .S(_1430_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4749_ (.A1(_1432_),
    .A2(\registers[6][27] ),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4750_ (.I0(_1273_),
    .I1(_1440_),
    .S(_1430_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4751_ (.A1(_1432_),
    .A2(\registers[6][28] ),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4752_ (.I(_1417_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4753_ (.I0(_1275_),
    .I1(_1441_),
    .S(_1442_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4754_ (.A1(_1432_),
    .A2(\registers[6][29] ),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4755_ (.I0(_1279_),
    .I1(_1443_),
    .S(_1442_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4756_ (.I(_1328_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4757_ (.A1(_1444_),
    .A2(\registers[6][2] ),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4758_ (.I0(_1281_),
    .I1(_1445_),
    .S(_1442_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4759_ (.A1(_1444_),
    .A2(\registers[6][30] ),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4760_ (.I0(_1283_),
    .I1(_1446_),
    .S(_1442_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4761_ (.A1(_1444_),
    .A2(\registers[6][31] ),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4762_ (.I0(_1088_),
    .I1(_1447_),
    .S(_1442_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4763_ (.A1(_1444_),
    .A2(\registers[6][3] ),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4764_ (.I0(_1098_),
    .I1(_1448_),
    .S(_1442_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4765_ (.A1(_1444_),
    .A2(\registers[6][4] ),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4766_ (.I0(_1100_),
    .I1(_1449_),
    .S(_1442_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4767_ (.A1(_1444_),
    .A2(\registers[6][5] ),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4768_ (.I0(_1102_),
    .I1(_1450_),
    .S(_1442_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4769_ (.A1(_1444_),
    .A2(\registers[6][6] ),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4770_ (.I0(_1104_),
    .I1(_1451_),
    .S(_1442_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4771_ (.A1(_1444_),
    .A2(\registers[6][7] ),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4772_ (.I0(_1106_),
    .I1(_1452_),
    .S(_1442_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4773_ (.A1(_1444_),
    .A2(\registers[6][8] ),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4774_ (.I0(_1108_),
    .I1(_1453_),
    .S(_1417_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4775_ (.A1(_1444_),
    .A2(\registers[6][9] ),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4776_ (.I0(_1110_),
    .I1(_1454_),
    .S(_1417_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4777_ (.I(_1089_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4778_ (.I(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4779_ (.A1(_1456_),
    .A2(\registers[7][0] ),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4780_ (.A1(_1232_),
    .A2(_1337_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4781_ (.I(_1458_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4782_ (.I0(_1229_),
    .I1(_1457_),
    .S(_1459_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4783_ (.A1(_1456_),
    .A2(\registers[7][10] ),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4784_ (.I0(_1235_),
    .I1(_1460_),
    .S(_1459_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4785_ (.A1(_1456_),
    .A2(\registers[7][11] ),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4786_ (.I0(_1237_),
    .I1(_1461_),
    .S(_1459_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4787_ (.A1(_1456_),
    .A2(\registers[7][12] ),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4788_ (.I0(_1239_),
    .I1(_1462_),
    .S(_1459_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4789_ (.A1(_1456_),
    .A2(\registers[7][13] ),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4790_ (.I0(_1241_),
    .I1(_1463_),
    .S(_1459_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4791_ (.A1(_1456_),
    .A2(\registers[7][14] ),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4792_ (.I0(_1243_),
    .I1(_1464_),
    .S(_1459_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4793_ (.A1(_1456_),
    .A2(\registers[7][15] ),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4794_ (.I0(_1245_),
    .I1(_1465_),
    .S(_1459_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4795_ (.A1(_1456_),
    .A2(\registers[7][16] ),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4796_ (.I0(_1247_),
    .I1(_1466_),
    .S(_1459_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4797_ (.A1(_1456_),
    .A2(\registers[7][17] ),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4798_ (.I0(_1249_),
    .I1(_1467_),
    .S(_1459_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4799_ (.A1(_1456_),
    .A2(\registers[7][18] ),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4800_ (.I0(_1251_),
    .I1(_1468_),
    .S(_1459_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4801_ (.I(_1455_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4802_ (.A1(_1469_),
    .A2(\registers[7][19] ),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4803_ (.I(_1458_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4804_ (.I0(_1253_),
    .I1(_1470_),
    .S(_1471_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4805_ (.A1(_1469_),
    .A2(\registers[7][1] ),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4806_ (.I0(_1257_),
    .I1(_1472_),
    .S(_1471_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4807_ (.A1(_1469_),
    .A2(\registers[7][20] ),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4808_ (.I0(_1259_),
    .I1(_1473_),
    .S(_1471_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4809_ (.A1(_1469_),
    .A2(\registers[7][21] ),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4810_ (.I0(_1261_),
    .I1(_1474_),
    .S(_1471_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4811_ (.A1(_1469_),
    .A2(\registers[7][22] ),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4812_ (.I0(_1263_),
    .I1(_1475_),
    .S(_1471_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4813_ (.A1(_1469_),
    .A2(\registers[7][23] ),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4814_ (.I0(_1265_),
    .I1(_1476_),
    .S(_1471_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4815_ (.A1(_1469_),
    .A2(\registers[7][24] ),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4816_ (.I0(_1267_),
    .I1(_1477_),
    .S(_1471_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4817_ (.A1(_1469_),
    .A2(\registers[7][25] ),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4818_ (.I0(_1269_),
    .I1(_1478_),
    .S(_1471_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4819_ (.A1(_1469_),
    .A2(\registers[7][26] ),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4820_ (.I0(_1271_),
    .I1(_1479_),
    .S(_1471_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4821_ (.A1(_1469_),
    .A2(\registers[7][27] ),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4822_ (.I0(_1273_),
    .I1(_1480_),
    .S(_1471_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _4823_ (.I(_1455_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4824_ (.A1(_1481_),
    .A2(\registers[7][28] ),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4825_ (.I(_1458_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4826_ (.I0(_1275_),
    .I1(_1482_),
    .S(_1483_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4827_ (.A1(_1481_),
    .A2(\registers[7][29] ),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4828_ (.I0(_1279_),
    .I1(_1484_),
    .S(_1483_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4829_ (.A1(_1481_),
    .A2(\registers[7][2] ),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4830_ (.I0(_1281_),
    .I1(_1485_),
    .S(_1483_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4831_ (.A1(_1481_),
    .A2(\registers[7][30] ),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4832_ (.I0(_1283_),
    .I1(_1486_),
    .S(_1483_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4833_ (.A1(_1481_),
    .A2(\registers[7][31] ),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4834_ (.I0(_1088_),
    .I1(_1487_),
    .S(_1483_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4835_ (.A1(_1481_),
    .A2(\registers[7][3] ),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4836_ (.I0(_1098_),
    .I1(_1488_),
    .S(_1483_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4837_ (.A1(_1481_),
    .A2(\registers[7][4] ),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4838_ (.I0(_1100_),
    .I1(_1489_),
    .S(_1483_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4839_ (.A1(_1481_),
    .A2(\registers[7][5] ),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4840_ (.I0(_1102_),
    .I1(_1490_),
    .S(_1483_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4841_ (.A1(_1481_),
    .A2(\registers[7][6] ),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4842_ (.I0(_1104_),
    .I1(_1491_),
    .S(_1483_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4843_ (.A1(_1481_),
    .A2(\registers[7][7] ),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4844_ (.I0(_1106_),
    .I1(_1492_),
    .S(_1483_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4845_ (.I(_1455_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4846_ (.A1(_1493_),
    .A2(\registers[7][8] ),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4847_ (.I0(_1108_),
    .I1(_1494_),
    .S(_1458_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4848_ (.A1(_1493_),
    .A2(\registers[7][9] ),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4849_ (.I0(_1110_),
    .I1(_1495_),
    .S(_1458_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4850_ (.A1(_1493_),
    .A2(\registers[8][0] ),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _4851_ (.I(net14),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _4852_ (.A1(net13),
    .A2(_1497_),
    .A3(_1335_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _4853_ (.A1(_1338_),
    .A2(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4854_ (.I(_1499_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4855_ (.I0(_1229_),
    .I1(_1496_),
    .S(_1500_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4856_ (.A1(_1493_),
    .A2(\registers[8][10] ),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4857_ (.I0(_1235_),
    .I1(_1501_),
    .S(_1500_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4858_ (.A1(_1493_),
    .A2(\registers[8][11] ),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4859_ (.I0(_1237_),
    .I1(_1502_),
    .S(_1500_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4860_ (.A1(_1493_),
    .A2(\registers[8][12] ),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4861_ (.I0(_1239_),
    .I1(_1503_),
    .S(_1500_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4862_ (.A1(_1493_),
    .A2(\registers[8][13] ),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4863_ (.I0(_1241_),
    .I1(_1504_),
    .S(_1500_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4864_ (.A1(_1493_),
    .A2(\registers[8][14] ),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4865_ (.I0(_1243_),
    .I1(_1505_),
    .S(_1500_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4866_ (.A1(_1493_),
    .A2(\registers[8][15] ),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4867_ (.I0(_1245_),
    .I1(_1506_),
    .S(_1500_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4868_ (.A1(_1493_),
    .A2(\registers[8][16] ),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4869_ (.I0(_1247_),
    .I1(_1507_),
    .S(_1500_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4870_ (.I(_1455_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4871_ (.A1(_1508_),
    .A2(\registers[8][17] ),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4872_ (.I0(_1249_),
    .I1(_1509_),
    .S(_1500_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4873_ (.A1(_1508_),
    .A2(\registers[8][18] ),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4874_ (.I0(_1251_),
    .I1(_1510_),
    .S(_1500_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4875_ (.A1(_1508_),
    .A2(\registers[8][19] ),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4876_ (.I(_1499_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4877_ (.I0(_1253_),
    .I1(_1511_),
    .S(_1512_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4878_ (.A1(_1508_),
    .A2(\registers[8][1] ),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4879_ (.I0(_1257_),
    .I1(_1513_),
    .S(_1512_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4880_ (.A1(_1508_),
    .A2(\registers[8][20] ),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4881_ (.I0(_1259_),
    .I1(_1514_),
    .S(_1512_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4882_ (.A1(_1508_),
    .A2(\registers[8][21] ),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4883_ (.I0(_1261_),
    .I1(_1515_),
    .S(_1512_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4884_ (.A1(_1508_),
    .A2(\registers[8][22] ),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4885_ (.I0(_1263_),
    .I1(_1516_),
    .S(_1512_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4886_ (.A1(_1508_),
    .A2(\registers[8][23] ),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4887_ (.I0(_1265_),
    .I1(_1517_),
    .S(_1512_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4888_ (.A1(_1508_),
    .A2(\registers[8][24] ),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4889_ (.I0(_1267_),
    .I1(_1518_),
    .S(_1512_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4890_ (.A1(_1508_),
    .A2(\registers[8][25] ),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4891_ (.I0(_1269_),
    .I1(_1519_),
    .S(_1512_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4892_ (.I(_1455_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4893_ (.A1(_1520_),
    .A2(\registers[8][26] ),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4894_ (.I0(_1271_),
    .I1(_1521_),
    .S(_1512_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4895_ (.A1(_1520_),
    .A2(\registers[8][27] ),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4896_ (.I0(_1273_),
    .I1(_1522_),
    .S(_1512_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4897_ (.A1(_1520_),
    .A2(\registers[8][28] ),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4898_ (.I(_1499_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4899_ (.I0(_1275_),
    .I1(_1523_),
    .S(_1524_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4900_ (.A1(_1520_),
    .A2(\registers[8][29] ),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4901_ (.I0(_1279_),
    .I1(_1525_),
    .S(_1524_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4902_ (.A1(_1520_),
    .A2(\registers[8][2] ),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4903_ (.I0(_1281_),
    .I1(_1526_),
    .S(_1524_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4904_ (.A1(_1520_),
    .A2(\registers[8][30] ),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4905_ (.I0(_1283_),
    .I1(_1527_),
    .S(_1524_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4906_ (.A1(_1520_),
    .A2(\registers[8][31] ),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4907_ (.I0(_1088_),
    .I1(_1528_),
    .S(_1524_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4908_ (.A1(_1520_),
    .A2(\registers[8][3] ),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4909_ (.I0(_1098_),
    .I1(_1529_),
    .S(_1524_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4910_ (.A1(_1520_),
    .A2(\registers[8][4] ),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4911_ (.I0(_1100_),
    .I1(_1530_),
    .S(_1524_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4912_ (.A1(_1520_),
    .A2(\registers[8][5] ),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4913_ (.I0(_1102_),
    .I1(_1531_),
    .S(_1524_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4914_ (.I(_1455_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4915_ (.A1(_1532_),
    .A2(\registers[8][6] ),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4916_ (.I0(_1104_),
    .I1(_1533_),
    .S(_1524_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4917_ (.A1(_1532_),
    .A2(\registers[8][7] ),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4918_ (.I0(_1106_),
    .I1(_1534_),
    .S(_1524_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4919_ (.A1(_1532_),
    .A2(\registers[8][8] ),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4920_ (.I0(_1108_),
    .I1(_1535_),
    .S(_1499_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4921_ (.A1(_1532_),
    .A2(\registers[8][9] ),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4922_ (.I0(_1110_),
    .I1(_1536_),
    .S(_1499_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4923_ (.A1(_1224_),
    .A2(\registers[9][0] ),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _4924_ (.A1(_1095_),
    .A2(_1498_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4925_ (.I(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4926_ (.I0(_1537_),
    .I1(_1115_),
    .S(_1539_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4927_ (.A1(_1224_),
    .A2(\registers[9][10] ),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4928_ (.I0(_1540_),
    .I1(_1123_),
    .S(_1539_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4929_ (.A1(_1224_),
    .A2(\registers[9][11] ),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4930_ (.I0(_1541_),
    .I1(_1125_),
    .S(_1539_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4931_ (.A1(_1224_),
    .A2(\registers[9][12] ),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4932_ (.I0(_1542_),
    .I1(_1127_),
    .S(_1539_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4933_ (.A1(_1224_),
    .A2(\registers[9][13] ),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4934_ (.I0(_1543_),
    .I1(_1129_),
    .S(_1539_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4935_ (.A1(_1224_),
    .A2(\registers[9][14] ),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4936_ (.I0(_1544_),
    .I1(_1131_),
    .S(_1539_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4937_ (.I(_1223_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4938_ (.A1(_1545_),
    .A2(\registers[9][15] ),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4939_ (.I0(_1546_),
    .I1(_1133_),
    .S(_1539_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4940_ (.A1(_1545_),
    .A2(\registers[9][16] ),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4941_ (.I0(_1547_),
    .I1(_1135_),
    .S(_1539_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4942_ (.A1(_1545_),
    .A2(\registers[9][17] ),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4943_ (.I0(_1548_),
    .I1(_1137_),
    .S(_1539_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4944_ (.A1(_1545_),
    .A2(\registers[9][18] ),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4945_ (.I0(_1549_),
    .I1(_1139_),
    .S(_1539_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4946_ (.A1(_1545_),
    .A2(\registers[9][19] ),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4947_ (.I(_1538_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4948_ (.I0(_1550_),
    .I1(_1142_),
    .S(_1551_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4949_ (.A1(_1545_),
    .A2(\registers[9][1] ),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4950_ (.I0(_1552_),
    .I1(_1145_),
    .S(_1551_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4951_ (.A1(_1545_),
    .A2(\registers[9][20] ),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4952_ (.I0(_1553_),
    .I1(_1147_),
    .S(_1551_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4953_ (.A1(_1545_),
    .A2(\registers[9][21] ),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4954_ (.I0(_1554_),
    .I1(_1149_),
    .S(_1551_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4955_ (.A1(_1545_),
    .A2(\registers[9][22] ),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4956_ (.I0(_1555_),
    .I1(_1151_),
    .S(_1551_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4957_ (.A1(_1545_),
    .A2(\registers[9][23] ),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4958_ (.I0(_1556_),
    .I1(_1153_),
    .S(_1551_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4959_ (.I(_1223_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4960_ (.A1(_1557_),
    .A2(\registers[9][24] ),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4961_ (.I0(_1558_),
    .I1(_1155_),
    .S(_1551_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4962_ (.A1(_1557_),
    .A2(\registers[9][25] ),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4963_ (.I0(_1559_),
    .I1(_1157_),
    .S(_1551_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4964_ (.A1(_1557_),
    .A2(\registers[9][26] ),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4965_ (.I0(_1560_),
    .I1(_1159_),
    .S(_1551_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4966_ (.A1(_1557_),
    .A2(\registers[9][27] ),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4967_ (.I0(_1561_),
    .I1(_1161_),
    .S(_1551_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4968_ (.A1(_1557_),
    .A2(\registers[9][28] ),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4969_ (.I(_1538_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4970_ (.I0(_1562_),
    .I1(_1164_),
    .S(_1563_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4971_ (.A1(_1557_),
    .A2(\registers[9][29] ),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4972_ (.I0(_1564_),
    .I1(_1167_),
    .S(_1563_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4973_ (.A1(_1557_),
    .A2(\registers[9][2] ),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4974_ (.I0(_1565_),
    .I1(_1169_),
    .S(_1563_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4975_ (.A1(_1557_),
    .A2(\registers[9][30] ),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4976_ (.I0(_1566_),
    .I1(_1171_),
    .S(_1563_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4977_ (.A1(_1557_),
    .A2(\registers[9][31] ),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4978_ (.I0(_1567_),
    .I1(_1173_),
    .S(_1563_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4979_ (.A1(_1557_),
    .A2(\registers[9][3] ),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4980_ (.I0(_1568_),
    .I1(_1175_),
    .S(_1563_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _4981_ (.I(_1223_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4982_ (.A1(_1569_),
    .A2(\registers[9][4] ),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4983_ (.I0(_1570_),
    .I1(_1177_),
    .S(_1563_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4984_ (.A1(_1569_),
    .A2(\registers[9][5] ),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4985_ (.I0(_1571_),
    .I1(_1179_),
    .S(_1563_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4986_ (.A1(_1569_),
    .A2(\registers[9][6] ),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4987_ (.I0(_1572_),
    .I1(_1181_),
    .S(_1563_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4988_ (.A1(_1569_),
    .A2(\registers[9][7] ),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4989_ (.I0(_1573_),
    .I1(_1183_),
    .S(_1563_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4990_ (.A1(_1569_),
    .A2(\registers[9][8] ),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4991_ (.I0(_1574_),
    .I1(_1186_),
    .S(_1538_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _4992_ (.A1(_1569_),
    .A2(\registers[9][9] ),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _4993_ (.I0(_1575_),
    .I1(_1188_),
    .S(_1538_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4994_ (.I(net2),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _4995_ (.I(_1576_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4996_ (.I(read_addr1[0]),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _4997_ (.I(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _4998_ (.I(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _4999_ (.I(read_addr1[1]),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5000_ (.I(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5001_ (.I0(\registers[28][0] ),
    .I1(\registers[29][0] ),
    .I2(\registers[30][0] ),
    .I3(\registers[31][0] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5002_ (.I(_1578_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5003_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5004_ (.I(_1581_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5005_ (.I0(\registers[24][0] ),
    .I1(\registers[25][0] ),
    .I2(\registers[26][0] ),
    .I3(\registers[27][0] ),
    .S0(_1585_),
    .S1(_1586_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _5006_ (.I(net1),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5007_ (.I(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5008_ (.I(_1589_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5009_ (.I0(_1583_),
    .I1(_1587_),
    .S(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5010_ (.I(read_addr1[1]),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5011_ (.A1(_1592_),
    .A2(_1588_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5012_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5013_ (.I(_1578_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5014_ (.I(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5015_ (.I0(\registers[18][0] ),
    .I1(\registers[19][0] ),
    .S(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5016_ (.I(_1597_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _5017_ (.A1(_1581_),
    .A2(net1),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5018_ (.I(_1599_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5019_ (.I(_1584_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5020_ (.I0(\registers[16][0] ),
    .I1(\registers[17][0] ),
    .S(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _5021_ (.A1(_1581_),
    .A2(net1),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5022_ (.I(_1603_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5023_ (.I(_1584_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5024_ (.I0(\registers[22][0] ),
    .I1(\registers[23][0] ),
    .S(_1605_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5025_ (.A1(_1600_),
    .A2(_1602_),
    .B1(_1604_),
    .B2(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5026_ (.A1(_1594_),
    .A2(_1598_),
    .B(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _5027_ (.A1(_1592_),
    .A2(_1588_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5028_ (.I(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5029_ (.I(_1595_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5030_ (.I0(\registers[20][0] ),
    .I1(\registers[21][0] ),
    .S(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5031_ (.I(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5032_ (.I(net2),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5033_ (.A1(_1610_),
    .A2(_1613_),
    .B(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _5034_ (.I(net3),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5035_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5036_ (.A1(_1577_),
    .A2(_1591_),
    .B1(_1608_),
    .B2(_1615_),
    .C(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5037_ (.A1(_1576_),
    .A2(_1616_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5038_ (.I(_1619_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5039_ (.I(_1579_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5040_ (.I(_1592_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5041_ (.I0(\registers[12][0] ),
    .I1(\registers[13][0] ),
    .I2(\registers[14][0] ),
    .I3(\registers[15][0] ),
    .S0(_1621_),
    .S1(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5042_ (.I(_1579_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5043_ (.I(_1592_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5044_ (.I0(\registers[8][0] ),
    .I1(\registers[9][0] ),
    .I2(\registers[10][0] ),
    .I3(\registers[11][0] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5045_ (.I(_1589_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5046_ (.I0(_1623_),
    .I1(_1626_),
    .S(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5047_ (.A1(net2),
    .A2(net3),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5048_ (.I(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5049_ (.I(_1578_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5050_ (.I0(\registers[0][0] ),
    .I1(\registers[1][0] ),
    .S(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _5051_ (.I(_1578_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5052_ (.I(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5053_ (.I0(\registers[2][0] ),
    .I1(\registers[3][0] ),
    .S(_1634_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5054_ (.I0(\registers[4][0] ),
    .I1(\registers[5][0] ),
    .S(_1595_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5055_ (.I0(\registers[6][0] ),
    .I1(\registers[7][0] ),
    .S(_1595_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5056_ (.I0(_1632_),
    .I1(_1635_),
    .I2(_1636_),
    .I3(_1637_),
    .S0(_1622_),
    .S1(net1),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5057_ (.I(net9),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5058_ (.A1(net7),
    .A2(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5059_ (.I(_1640_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5060_ (.A1(_1620_),
    .A2(_1628_),
    .B1(_1630_),
    .B2(_1638_),
    .C(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5061_ (.I(net7),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5062_ (.A1(_1643_),
    .A2(_1639_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5063_ (.I(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5064_ (.A1(net48),
    .A2(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5065_ (.A1(_1618_),
    .A2(_1642_),
    .B(_1646_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5066_ (.I0(\registers[12][10] ),
    .I1(\registers[13][10] ),
    .I2(\registers[14][10] ),
    .I3(\registers[15][10] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5067_ (.I0(\registers[8][10] ),
    .I1(\registers[9][10] ),
    .I2(\registers[10][10] ),
    .I3(\registers[11][10] ),
    .S0(_1585_),
    .S1(_1586_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5068_ (.I0(_1647_),
    .I1(_1648_),
    .S(_1590_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5069_ (.I0(\registers[2][10] ),
    .I1(\registers[3][10] ),
    .S(_1596_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5070_ (.I(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5071_ (.I0(\registers[0][10] ),
    .I1(\registers[1][10] ),
    .S(_1601_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5072_ (.I(_1584_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5073_ (.I0(\registers[6][10] ),
    .I1(\registers[7][10] ),
    .S(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5074_ (.A1(_1600_),
    .A2(_1652_),
    .B1(_1654_),
    .B2(_1604_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5075_ (.A1(_1594_),
    .A2(_1651_),
    .B(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5076_ (.I0(\registers[4][10] ),
    .I1(\registers[5][10] ),
    .S(_1611_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5077_ (.I(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5078_ (.A1(_1610_),
    .A2(_1658_),
    .B(_1614_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5079_ (.I(net3),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5080_ (.A1(_1577_),
    .A2(_1649_),
    .B1(_1656_),
    .B2(_1659_),
    .C(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _5081_ (.A1(_1576_),
    .A2(net3),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5082_ (.I(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5083_ (.I0(\registers[28][10] ),
    .I1(\registers[29][10] ),
    .I2(\registers[30][10] ),
    .I3(\registers[31][10] ),
    .S0(_1621_),
    .S1(_1622_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5084_ (.I0(\registers[24][10] ),
    .I1(\registers[25][10] ),
    .I2(\registers[26][10] ),
    .I3(\registers[27][10] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5085_ (.I0(_1664_),
    .I1(_1665_),
    .S(_1627_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5086_ (.A1(net2),
    .A2(_1616_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5087_ (.I(_1667_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5088_ (.I0(\registers[16][10] ),
    .I1(\registers[17][10] ),
    .S(_1631_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5089_ (.I0(\registers[18][10] ),
    .I1(\registers[19][10] ),
    .S(_1634_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5090_ (.I0(\registers[20][10] ),
    .I1(\registers[21][10] ),
    .S(_1595_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5091_ (.I0(\registers[22][10] ),
    .I1(\registers[23][10] ),
    .S(_1595_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5092_ (.I0(_1669_),
    .I1(_1670_),
    .I2(_1671_),
    .I3(_1672_),
    .S0(_1622_),
    .S1(net1),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5093_ (.A1(_1663_),
    .A2(_1666_),
    .B1(_1668_),
    .B2(_1673_),
    .C(_1641_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5094_ (.A1(net49),
    .A2(_1645_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5095_ (.A1(_1661_),
    .A2(_1674_),
    .B(_1675_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5096_ (.I(_1579_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5097_ (.I0(\registers[12][11] ),
    .I1(\registers[13][11] ),
    .I2(\registers[14][11] ),
    .I3(\registers[15][11] ),
    .S0(_1676_),
    .S1(_1582_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5098_ (.I(_1581_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5099_ (.I0(\registers[8][11] ),
    .I1(\registers[9][11] ),
    .I2(\registers[10][11] ),
    .I3(\registers[11][11] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5100_ (.I0(_1677_),
    .I1(_1679_),
    .S(_1590_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5101_ (.I0(\registers[2][11] ),
    .I1(\registers[3][11] ),
    .S(_1596_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5102_ (.I(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5103_ (.I0(\registers[0][11] ),
    .I1(\registers[1][11] ),
    .S(_1601_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5104_ (.I0(\registers[6][11] ),
    .I1(\registers[7][11] ),
    .S(_1653_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5105_ (.A1(_1600_),
    .A2(_1683_),
    .B1(_1684_),
    .B2(_1604_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5106_ (.A1(_1594_),
    .A2(_1682_),
    .B(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5107_ (.I0(\registers[4][11] ),
    .I1(\registers[5][11] ),
    .S(_1611_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5108_ (.I(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5109_ (.A1(_1610_),
    .A2(_1688_),
    .B(_1614_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5110_ (.A1(_1577_),
    .A2(_1680_),
    .B1(_1686_),
    .B2(_1689_),
    .C(_1660_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5111_ (.I0(\registers[28][11] ),
    .I1(\registers[29][11] ),
    .I2(\registers[30][11] ),
    .I3(\registers[31][11] ),
    .S0(_1621_),
    .S1(_1622_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5112_ (.I0(\registers[24][11] ),
    .I1(\registers[25][11] ),
    .I2(\registers[26][11] ),
    .I3(\registers[27][11] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5113_ (.I0(_1691_),
    .I1(_1692_),
    .S(_1627_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5114_ (.I(_1633_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5115_ (.I0(\registers[16][11] ),
    .I1(\registers[17][11] ),
    .S(_1694_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5116_ (.I0(\registers[18][11] ),
    .I1(\registers[19][11] ),
    .S(_1605_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5117_ (.I0(\registers[20][11] ),
    .I1(\registers[21][11] ),
    .S(_1634_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5118_ (.I(_1633_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5119_ (.I0(\registers[22][11] ),
    .I1(\registers[23][11] ),
    .S(_1698_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5120_ (.I(_1592_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5121_ (.I(net1),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5122_ (.I0(_1695_),
    .I1(_1696_),
    .I2(_1697_),
    .I3(_1699_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5123_ (.A1(_1663_),
    .A2(_1693_),
    .B1(_1702_),
    .B2(_1668_),
    .C(_1641_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5124_ (.A1(net50),
    .A2(_1645_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5125_ (.A1(_1690_),
    .A2(_1703_),
    .B(_1704_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5126_ (.I0(\registers[12][12] ),
    .I1(\registers[13][12] ),
    .I2(\registers[14][12] ),
    .I3(\registers[15][12] ),
    .S0(_1676_),
    .S1(_1582_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5127_ (.I0(\registers[8][12] ),
    .I1(\registers[9][12] ),
    .I2(\registers[10][12] ),
    .I3(\registers[11][12] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5128_ (.I0(_1705_),
    .I1(_1706_),
    .S(_1590_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5129_ (.I0(\registers[2][12] ),
    .I1(\registers[3][12] ),
    .S(_1596_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5130_ (.I(_1708_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5131_ (.I0(\registers[0][12] ),
    .I1(\registers[1][12] ),
    .S(_1601_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5132_ (.I0(\registers[6][12] ),
    .I1(\registers[7][12] ),
    .S(_1653_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5133_ (.A1(_1600_),
    .A2(_1710_),
    .B1(_1711_),
    .B2(_1604_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5134_ (.A1(_1594_),
    .A2(_1709_),
    .B(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5135_ (.I0(\registers[4][12] ),
    .I1(\registers[5][12] ),
    .S(_1611_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5136_ (.I(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5137_ (.A1(_1610_),
    .A2(_1715_),
    .B(_1614_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5138_ (.A1(_1577_),
    .A2(_1707_),
    .B1(_1713_),
    .B2(_1716_),
    .C(_1660_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5139_ (.I0(\registers[28][12] ),
    .I1(\registers[29][12] ),
    .I2(\registers[30][12] ),
    .I3(\registers[31][12] ),
    .S0(_1621_),
    .S1(_1622_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5140_ (.I0(\registers[24][12] ),
    .I1(\registers[25][12] ),
    .I2(\registers[26][12] ),
    .I3(\registers[27][12] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5141_ (.I0(_1718_),
    .I1(_1719_),
    .S(_1627_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5142_ (.I0(\registers[16][12] ),
    .I1(\registers[17][12] ),
    .S(_1694_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5143_ (.I0(\registers[18][12] ),
    .I1(\registers[19][12] ),
    .S(_1605_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5144_ (.I0(\registers[20][12] ),
    .I1(\registers[21][12] ),
    .S(_1634_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5145_ (.I0(\registers[22][12] ),
    .I1(\registers[23][12] ),
    .S(_1698_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5146_ (.I0(_1721_),
    .I1(_1722_),
    .I2(_1723_),
    .I3(_1724_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5147_ (.A1(_1663_),
    .A2(_1720_),
    .B1(_1725_),
    .B2(_1668_),
    .C(_1641_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5148_ (.A1(net51),
    .A2(_1645_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5149_ (.A1(_1717_),
    .A2(_1726_),
    .B(_1727_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5150_ (.I(_1581_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5151_ (.I0(\registers[12][13] ),
    .I1(\registers[13][13] ),
    .I2(\registers[14][13] ),
    .I3(\registers[15][13] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5152_ (.I0(\registers[8][13] ),
    .I1(\registers[9][13] ),
    .I2(\registers[10][13] ),
    .I3(\registers[11][13] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5153_ (.I0(_1729_),
    .I1(_1730_),
    .S(_1590_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5154_ (.I0(\registers[2][13] ),
    .I1(\registers[3][13] ),
    .S(_1596_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5155_ (.I(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5156_ (.I0(\registers[0][13] ),
    .I1(\registers[1][13] ),
    .S(_1601_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5157_ (.I0(\registers[6][13] ),
    .I1(\registers[7][13] ),
    .S(_1653_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5158_ (.A1(_1600_),
    .A2(_1734_),
    .B1(_1735_),
    .B2(_1604_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5159_ (.A1(_1594_),
    .A2(_1733_),
    .B(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5160_ (.I0(\registers[4][13] ),
    .I1(\registers[5][13] ),
    .S(_1611_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5161_ (.I(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5162_ (.A1(_1610_),
    .A2(_1739_),
    .B(_1614_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5163_ (.A1(_1577_),
    .A2(_1731_),
    .B1(_1737_),
    .B2(_1740_),
    .C(_1660_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5164_ (.I0(\registers[28][13] ),
    .I1(\registers[29][13] ),
    .I2(\registers[30][13] ),
    .I3(\registers[31][13] ),
    .S0(_1621_),
    .S1(_1622_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5165_ (.I(_1579_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5166_ (.I0(\registers[24][13] ),
    .I1(\registers[25][13] ),
    .I2(\registers[26][13] ),
    .I3(\registers[27][13] ),
    .S0(_1743_),
    .S1(_1625_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5167_ (.I0(_1742_),
    .I1(_1744_),
    .S(_1627_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5168_ (.I0(\registers[16][13] ),
    .I1(\registers[17][13] ),
    .S(_1694_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5169_ (.I0(\registers[18][13] ),
    .I1(\registers[19][13] ),
    .S(_1605_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5170_ (.I(_1633_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5171_ (.I0(\registers[20][13] ),
    .I1(\registers[21][13] ),
    .S(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5172_ (.I0(\registers[22][13] ),
    .I1(\registers[23][13] ),
    .S(_1698_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5173_ (.I0(_1746_),
    .I1(_1747_),
    .I2(_1749_),
    .I3(_1750_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5174_ (.A1(_1663_),
    .A2(_1745_),
    .B1(_1751_),
    .B2(_1668_),
    .C(_1641_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5175_ (.A1(net52),
    .A2(_1645_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5176_ (.A1(_1741_),
    .A2(_1752_),
    .B(_1753_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5177_ (.I0(\registers[28][14] ),
    .I1(\registers[29][14] ),
    .I2(\registers[30][14] ),
    .I3(\registers[31][14] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5178_ (.I0(\registers[24][14] ),
    .I1(\registers[25][14] ),
    .I2(\registers[26][14] ),
    .I3(\registers[27][14] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5179_ (.I0(_1754_),
    .I1(_1755_),
    .S(_1590_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5180_ (.I0(\registers[18][14] ),
    .I1(\registers[19][14] ),
    .S(_1596_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5181_ (.I(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5182_ (.I0(\registers[16][14] ),
    .I1(\registers[17][14] ),
    .S(_1601_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5183_ (.I0(\registers[22][14] ),
    .I1(\registers[23][14] ),
    .S(_1653_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5184_ (.A1(_1600_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(_1604_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5185_ (.A1(_1594_),
    .A2(_1758_),
    .B(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5186_ (.I0(\registers[20][14] ),
    .I1(\registers[21][14] ),
    .S(_1611_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5187_ (.I(_1763_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5188_ (.A1(_1610_),
    .A2(_1764_),
    .B(_1614_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5189_ (.A1(_1577_),
    .A2(_1756_),
    .B1(_1762_),
    .B2(_1765_),
    .C(_1617_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5190_ (.I0(\registers[12][14] ),
    .I1(\registers[13][14] ),
    .I2(\registers[14][14] ),
    .I3(\registers[15][14] ),
    .S0(_1621_),
    .S1(_1622_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5191_ (.I0(\registers[8][14] ),
    .I1(\registers[9][14] ),
    .I2(\registers[10][14] ),
    .I3(\registers[11][14] ),
    .S0(_1743_),
    .S1(_1625_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5192_ (.I0(_1767_),
    .I1(_1768_),
    .S(_1627_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5193_ (.I0(\registers[0][14] ),
    .I1(\registers[1][14] ),
    .S(_1694_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5194_ (.I0(\registers[2][14] ),
    .I1(\registers[3][14] ),
    .S(_1605_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5195_ (.I0(\registers[4][14] ),
    .I1(\registers[5][14] ),
    .S(_1748_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5196_ (.I0(\registers[6][14] ),
    .I1(\registers[7][14] ),
    .S(_1698_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5197_ (.I0(_1770_),
    .I1(_1771_),
    .I2(_1772_),
    .I3(_1773_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5198_ (.A1(_1620_),
    .A2(_1769_),
    .B1(_1774_),
    .B2(_1630_),
    .C(_1641_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5199_ (.A1(net53),
    .A2(_1645_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5200_ (.A1(_1766_),
    .A2(_1775_),
    .B(_1776_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5201_ (.I0(\registers[12][15] ),
    .I1(\registers[13][15] ),
    .I2(\registers[14][15] ),
    .I3(\registers[15][15] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5202_ (.I0(\registers[8][15] ),
    .I1(\registers[9][15] ),
    .I2(\registers[10][15] ),
    .I3(\registers[11][15] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5203_ (.I0(_1777_),
    .I1(_1778_),
    .S(_1590_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5204_ (.I0(\registers[2][15] ),
    .I1(\registers[3][15] ),
    .S(_1596_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5205_ (.I(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5206_ (.I0(\registers[0][15] ),
    .I1(\registers[1][15] ),
    .S(_1601_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5207_ (.I0(\registers[6][15] ),
    .I1(\registers[7][15] ),
    .S(_1653_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5208_ (.A1(_1600_),
    .A2(_1782_),
    .B1(_1783_),
    .B2(_1604_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5209_ (.A1(_1594_),
    .A2(_1781_),
    .B(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5210_ (.I0(\registers[4][15] ),
    .I1(\registers[5][15] ),
    .S(_1611_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5211_ (.I(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5212_ (.A1(_1610_),
    .A2(_1787_),
    .B(_1614_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5213_ (.A1(_1577_),
    .A2(_1779_),
    .B1(_1785_),
    .B2(_1788_),
    .C(_1660_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5214_ (.I(_1579_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5215_ (.I0(\registers[28][15] ),
    .I1(\registers[29][15] ),
    .I2(\registers[30][15] ),
    .I3(\registers[31][15] ),
    .S0(_1790_),
    .S1(_1622_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5216_ (.I(_1592_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5217_ (.I0(\registers[24][15] ),
    .I1(\registers[25][15] ),
    .I2(\registers[26][15] ),
    .I3(\registers[27][15] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5218_ (.I0(_1791_),
    .I1(_1793_),
    .S(_1627_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5219_ (.I(_1633_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5220_ (.I0(\registers[16][15] ),
    .I1(\registers[17][15] ),
    .S(_1795_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5221_ (.I(_1633_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5222_ (.I0(\registers[18][15] ),
    .I1(\registers[19][15] ),
    .S(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5223_ (.I0(\registers[20][15] ),
    .I1(\registers[21][15] ),
    .S(_1748_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5224_ (.I(_1633_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5225_ (.I0(\registers[22][15] ),
    .I1(\registers[23][15] ),
    .S(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5226_ (.I0(_1796_),
    .I1(_1798_),
    .I2(_1799_),
    .I3(_1801_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5227_ (.A1(_1663_),
    .A2(_1794_),
    .B1(_1802_),
    .B2(_1668_),
    .C(_1641_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5228_ (.A1(net54),
    .A2(_1645_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5229_ (.A1(_1789_),
    .A2(_1803_),
    .B(_1804_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5230_ (.I0(\registers[28][16] ),
    .I1(\registers[29][16] ),
    .I2(\registers[30][16] ),
    .I3(\registers[31][16] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5231_ (.I0(\registers[24][16] ),
    .I1(\registers[25][16] ),
    .I2(\registers[26][16] ),
    .I3(\registers[27][16] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5232_ (.I0(_1805_),
    .I1(_1806_),
    .S(_1590_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5233_ (.I0(\registers[18][16] ),
    .I1(\registers[19][16] ),
    .S(_1596_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5234_ (.I(_1808_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5235_ (.I0(\registers[16][16] ),
    .I1(\registers[17][16] ),
    .S(_1601_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5236_ (.I(_1584_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5237_ (.I0(\registers[22][16] ),
    .I1(\registers[23][16] ),
    .S(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5238_ (.A1(_1600_),
    .A2(_1810_),
    .B1(_1812_),
    .B2(_1604_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5239_ (.A1(_1594_),
    .A2(_1809_),
    .B(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5240_ (.I0(\registers[20][16] ),
    .I1(\registers[21][16] ),
    .S(_1611_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5241_ (.I(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5242_ (.A1(_1610_),
    .A2(_1816_),
    .B(_1614_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5243_ (.A1(_1577_),
    .A2(_1807_),
    .B1(_1814_),
    .B2(_1817_),
    .C(_1617_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5244_ (.I0(\registers[12][16] ),
    .I1(\registers[13][16] ),
    .I2(\registers[14][16] ),
    .I3(\registers[15][16] ),
    .S0(_1790_),
    .S1(_1622_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5245_ (.I0(\registers[8][16] ),
    .I1(\registers[9][16] ),
    .I2(\registers[10][16] ),
    .I3(\registers[11][16] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5246_ (.I0(_1819_),
    .I1(_1820_),
    .S(_1627_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5247_ (.I0(\registers[0][16] ),
    .I1(\registers[1][16] ),
    .S(_1795_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5248_ (.I0(\registers[2][16] ),
    .I1(\registers[3][16] ),
    .S(_1797_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5249_ (.I0(\registers[4][16] ),
    .I1(\registers[5][16] ),
    .S(_1748_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5250_ (.I0(\registers[6][16] ),
    .I1(\registers[7][16] ),
    .S(_1800_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5251_ (.I0(_1822_),
    .I1(_1823_),
    .I2(_1824_),
    .I3(_1825_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5252_ (.A1(_1620_),
    .A2(_1821_),
    .B1(_1826_),
    .B2(_1630_),
    .C(_1641_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5253_ (.A1(net55),
    .A2(_1645_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5254_ (.A1(_1818_),
    .A2(_1827_),
    .B(_1828_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5255_ (.I0(\registers[28][17] ),
    .I1(\registers[29][17] ),
    .I2(\registers[30][17] ),
    .I3(\registers[31][17] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5256_ (.I0(\registers[24][17] ),
    .I1(\registers[25][17] ),
    .I2(\registers[26][17] ),
    .I3(\registers[27][17] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5257_ (.I(_1589_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5258_ (.I0(_1829_),
    .I1(_1830_),
    .S(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5259_ (.I0(\registers[18][17] ),
    .I1(\registers[19][17] ),
    .S(_1596_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5260_ (.I(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5261_ (.I(_1584_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5262_ (.I0(\registers[16][17] ),
    .I1(\registers[17][17] ),
    .S(_1835_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5263_ (.I0(\registers[22][17] ),
    .I1(\registers[23][17] ),
    .S(_1811_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5264_ (.A1(_1600_),
    .A2(_1836_),
    .B1(_1837_),
    .B2(_1604_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5265_ (.A1(_1594_),
    .A2(_1834_),
    .B(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5266_ (.I(_1595_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5267_ (.I0(\registers[20][17] ),
    .I1(\registers[21][17] ),
    .S(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5268_ (.I(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5269_ (.I(_1576_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5270_ (.A1(_1610_),
    .A2(_1842_),
    .B(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5271_ (.A1(_1577_),
    .A2(_1832_),
    .B1(_1839_),
    .B2(_1844_),
    .C(_1617_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5272_ (.I(_1592_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5273_ (.I0(\registers[12][17] ),
    .I1(\registers[13][17] ),
    .I2(\registers[14][17] ),
    .I3(\registers[15][17] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5274_ (.I0(\registers[8][17] ),
    .I1(\registers[9][17] ),
    .I2(\registers[10][17] ),
    .I3(\registers[11][17] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5275_ (.I0(_1847_),
    .I1(_1848_),
    .S(_1627_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5276_ (.I0(\registers[0][17] ),
    .I1(\registers[1][17] ),
    .S(_1795_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5277_ (.I0(\registers[2][17] ),
    .I1(\registers[3][17] ),
    .S(_1797_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5278_ (.I0(\registers[4][17] ),
    .I1(\registers[5][17] ),
    .S(_1748_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5279_ (.I0(\registers[6][17] ),
    .I1(\registers[7][17] ),
    .S(_1800_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5280_ (.I0(_1850_),
    .I1(_1851_),
    .I2(_1852_),
    .I3(_1853_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5281_ (.A1(_1620_),
    .A2(_1849_),
    .B1(_1854_),
    .B2(_1630_),
    .C(_1641_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5282_ (.A1(net56),
    .A2(_1645_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5283_ (.A1(_1845_),
    .A2(_1855_),
    .B(_1856_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5284_ (.I0(\registers[12][18] ),
    .I1(\registers[13][18] ),
    .I2(\registers[14][18] ),
    .I3(\registers[15][18] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5285_ (.I0(\registers[8][18] ),
    .I1(\registers[9][18] ),
    .I2(\registers[10][18] ),
    .I3(\registers[11][18] ),
    .S0(_1585_),
    .S1(_1678_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5286_ (.I0(_1857_),
    .I1(_1858_),
    .S(_1831_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5287_ (.I0(\registers[2][18] ),
    .I1(\registers[3][18] ),
    .S(_1596_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5288_ (.I(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5289_ (.I0(\registers[0][18] ),
    .I1(\registers[1][18] ),
    .S(_1835_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5290_ (.I0(\registers[6][18] ),
    .I1(\registers[7][18] ),
    .S(_1811_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5291_ (.A1(_1600_),
    .A2(_1862_),
    .B1(_1863_),
    .B2(_1604_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5292_ (.A1(_1594_),
    .A2(_1861_),
    .B(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5293_ (.I0(\registers[4][18] ),
    .I1(\registers[5][18] ),
    .S(_1840_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5294_ (.I(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5295_ (.A1(_1610_),
    .A2(_1867_),
    .B(_1843_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5296_ (.A1(_1577_),
    .A2(_1859_),
    .B1(_1865_),
    .B2(_1868_),
    .C(_1660_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5297_ (.I0(\registers[28][18] ),
    .I1(\registers[29][18] ),
    .I2(\registers[30][18] ),
    .I3(\registers[31][18] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5298_ (.I0(\registers[24][18] ),
    .I1(\registers[25][18] ),
    .I2(\registers[26][18] ),
    .I3(\registers[27][18] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5299_ (.I0(_1870_),
    .I1(_1871_),
    .S(_1627_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5300_ (.I0(\registers[16][18] ),
    .I1(\registers[17][18] ),
    .S(_1795_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5301_ (.I0(\registers[18][18] ),
    .I1(\registers[19][18] ),
    .S(_1797_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5302_ (.I0(\registers[20][18] ),
    .I1(\registers[21][18] ),
    .S(_1748_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5303_ (.I0(\registers[22][18] ),
    .I1(\registers[23][18] ),
    .S(_1800_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5304_ (.I0(_1873_),
    .I1(_1874_),
    .I2(_1875_),
    .I3(_1876_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5305_ (.A1(_1663_),
    .A2(_1872_),
    .B1(_1877_),
    .B2(_1668_),
    .C(_1641_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5306_ (.A1(net57),
    .A2(_1645_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5307_ (.A1(_1869_),
    .A2(_1878_),
    .B(_1879_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5308_ (.I(_1576_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5309_ (.I0(\registers[12][19] ),
    .I1(\registers[13][19] ),
    .I2(\registers[14][19] ),
    .I3(\registers[15][19] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5310_ (.I(_1584_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5311_ (.I0(\registers[8][19] ),
    .I1(\registers[9][19] ),
    .I2(\registers[10][19] ),
    .I3(\registers[11][19] ),
    .S0(_1882_),
    .S1(_1678_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5312_ (.I0(_1881_),
    .I1(_1883_),
    .S(_1831_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5313_ (.I(_1593_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5314_ (.I(_1595_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5315_ (.I0(\registers[2][19] ),
    .I1(\registers[3][19] ),
    .S(_1886_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5316_ (.I(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5317_ (.I(_1599_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5318_ (.I0(\registers[0][19] ),
    .I1(\registers[1][19] ),
    .S(_1835_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5319_ (.I0(\registers[6][19] ),
    .I1(\registers[7][19] ),
    .S(_1811_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5320_ (.I(_1603_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5321_ (.A1(_1889_),
    .A2(_1890_),
    .B1(_1891_),
    .B2(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5322_ (.A1(_1885_),
    .A2(_1888_),
    .B(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5323_ (.I(_1609_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5324_ (.I0(\registers[4][19] ),
    .I1(\registers[5][19] ),
    .S(_1840_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5325_ (.I(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5326_ (.A1(_1895_),
    .A2(_1897_),
    .B(_1843_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5327_ (.A1(_1880_),
    .A2(_1884_),
    .B1(_1894_),
    .B2(_1898_),
    .C(_1660_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5328_ (.I0(\registers[28][19] ),
    .I1(\registers[29][19] ),
    .I2(\registers[30][19] ),
    .I3(\registers[31][19] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5329_ (.I0(\registers[24][19] ),
    .I1(\registers[25][19] ),
    .I2(\registers[26][19] ),
    .I3(\registers[27][19] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5330_ (.I(_1589_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5331_ (.I0(_1900_),
    .I1(_1901_),
    .S(_1902_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5332_ (.I0(\registers[16][19] ),
    .I1(\registers[17][19] ),
    .S(_1795_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5333_ (.I0(\registers[18][19] ),
    .I1(\registers[19][19] ),
    .S(_1797_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5334_ (.I0(\registers[20][19] ),
    .I1(\registers[21][19] ),
    .S(_1748_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5335_ (.I0(\registers[22][19] ),
    .I1(\registers[23][19] ),
    .S(_1800_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5336_ (.I0(_1904_),
    .I1(_1905_),
    .I2(_1906_),
    .I3(_1907_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5337_ (.I(_1640_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5338_ (.A1(_1663_),
    .A2(_1903_),
    .B1(_1908_),
    .B2(_1668_),
    .C(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5339_ (.I(_1644_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5340_ (.A1(net58),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5341_ (.A1(_1899_),
    .A2(_1910_),
    .B(_1912_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5342_ (.I0(\registers[12][1] ),
    .I1(\registers[13][1] ),
    .I2(\registers[14][1] ),
    .I3(\registers[15][1] ),
    .S0(_1676_),
    .S1(_1728_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5343_ (.I0(\registers[8][1] ),
    .I1(\registers[9][1] ),
    .I2(\registers[10][1] ),
    .I3(\registers[11][1] ),
    .S0(_1882_),
    .S1(_1678_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5344_ (.I0(_1913_),
    .I1(_1914_),
    .S(_1831_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5345_ (.I0(\registers[2][1] ),
    .I1(\registers[3][1] ),
    .S(_1886_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5346_ (.I(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5347_ (.I0(\registers[0][1] ),
    .I1(\registers[1][1] ),
    .S(_1835_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5348_ (.I0(\registers[6][1] ),
    .I1(\registers[7][1] ),
    .S(_1811_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5349_ (.A1(_1889_),
    .A2(_1918_),
    .B1(_1919_),
    .B2(_1892_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5350_ (.A1(_1885_),
    .A2(_1917_),
    .B(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5351_ (.I0(\registers[4][1] ),
    .I1(\registers[5][1] ),
    .S(_1840_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5352_ (.I(_1922_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5353_ (.A1(_1895_),
    .A2(_1923_),
    .B(_1843_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5354_ (.A1(_1880_),
    .A2(_1915_),
    .B1(_1921_),
    .B2(_1924_),
    .C(_1660_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5355_ (.I0(\registers[28][1] ),
    .I1(\registers[29][1] ),
    .I2(\registers[30][1] ),
    .I3(\registers[31][1] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5356_ (.I0(\registers[24][1] ),
    .I1(\registers[25][1] ),
    .I2(\registers[26][1] ),
    .I3(\registers[27][1] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5357_ (.I0(_1926_),
    .I1(_1927_),
    .S(_1902_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5358_ (.I0(\registers[16][1] ),
    .I1(\registers[17][1] ),
    .S(_1795_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5359_ (.I0(\registers[18][1] ),
    .I1(\registers[19][1] ),
    .S(_1797_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5360_ (.I0(\registers[20][1] ),
    .I1(\registers[21][1] ),
    .S(_1748_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5361_ (.I0(\registers[22][1] ),
    .I1(\registers[23][1] ),
    .S(_1800_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5362_ (.I0(_1929_),
    .I1(_1930_),
    .I2(_1931_),
    .I3(_1932_),
    .S0(_1700_),
    .S1(_1701_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5363_ (.A1(_1663_),
    .A2(_1928_),
    .B1(_1933_),
    .B2(_1668_),
    .C(_1909_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5364_ (.A1(net59),
    .A2(_1911_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5365_ (.A1(_1925_),
    .A2(_1934_),
    .B(_1935_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5366_ (.I(_1579_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5367_ (.I0(\registers[12][20] ),
    .I1(\registers[13][20] ),
    .I2(\registers[14][20] ),
    .I3(\registers[15][20] ),
    .S0(_1936_),
    .S1(_1728_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5368_ (.I(_1581_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5369_ (.I0(\registers[8][20] ),
    .I1(\registers[9][20] ),
    .I2(\registers[10][20] ),
    .I3(\registers[11][20] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5370_ (.I0(_1937_),
    .I1(_1939_),
    .S(_1831_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5371_ (.I0(\registers[2][20] ),
    .I1(\registers[3][20] ),
    .S(_1886_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5372_ (.I(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5373_ (.I0(\registers[0][20] ),
    .I1(\registers[1][20] ),
    .S(_1835_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5374_ (.I0(\registers[6][20] ),
    .I1(\registers[7][20] ),
    .S(_1811_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5375_ (.A1(_1889_),
    .A2(_1943_),
    .B1(_1944_),
    .B2(_1892_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5376_ (.A1(_1885_),
    .A2(_1942_),
    .B(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5377_ (.I0(\registers[4][20] ),
    .I1(\registers[5][20] ),
    .S(_1840_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5378_ (.I(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5379_ (.A1(_1895_),
    .A2(_1948_),
    .B(_1843_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5380_ (.A1(_1880_),
    .A2(_1940_),
    .B1(_1946_),
    .B2(_1949_),
    .C(_1660_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5381_ (.I0(\registers[28][20] ),
    .I1(\registers[29][20] ),
    .I2(\registers[30][20] ),
    .I3(\registers[31][20] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5382_ (.I0(\registers[24][20] ),
    .I1(\registers[25][20] ),
    .I2(\registers[26][20] ),
    .I3(\registers[27][20] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5383_ (.I0(_1951_),
    .I1(_1952_),
    .S(_1902_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5384_ (.I0(\registers[16][20] ),
    .I1(\registers[17][20] ),
    .S(_1795_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5385_ (.I0(\registers[18][20] ),
    .I1(\registers[19][20] ),
    .S(_1797_),
    .Z(_1955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5386_ (.I0(\registers[20][20] ),
    .I1(\registers[21][20] ),
    .S(_1748_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5387_ (.I0(\registers[22][20] ),
    .I1(\registers[23][20] ),
    .S(_1800_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5388_ (.I(_1592_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5389_ (.I(net1),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5390_ (.I0(_1954_),
    .I1(_1955_),
    .I2(_1956_),
    .I3(_1957_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5391_ (.A1(_1663_),
    .A2(_1953_),
    .B1(_1960_),
    .B2(_1668_),
    .C(_1909_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5392_ (.A1(net60),
    .A2(_1911_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5393_ (.A1(_1950_),
    .A2(_1961_),
    .B(_1962_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5394_ (.I0(\registers[12][21] ),
    .I1(\registers[13][21] ),
    .I2(\registers[14][21] ),
    .I3(\registers[15][21] ),
    .S0(_1936_),
    .S1(_1728_),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5395_ (.I0(\registers[8][21] ),
    .I1(\registers[9][21] ),
    .I2(\registers[10][21] ),
    .I3(\registers[11][21] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5396_ (.I0(_1963_),
    .I1(_1964_),
    .S(_1831_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5397_ (.I0(\registers[2][21] ),
    .I1(\registers[3][21] ),
    .S(_1886_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5398_ (.I(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5399_ (.I0(\registers[0][21] ),
    .I1(\registers[1][21] ),
    .S(_1835_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5400_ (.I0(\registers[6][21] ),
    .I1(\registers[7][21] ),
    .S(_1811_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5401_ (.A1(_1889_),
    .A2(_1968_),
    .B1(_1969_),
    .B2(_1892_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5402_ (.A1(_1885_),
    .A2(_1967_),
    .B(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5403_ (.I0(\registers[4][21] ),
    .I1(\registers[5][21] ),
    .S(_1840_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5404_ (.I(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5405_ (.A1(_1895_),
    .A2(_1973_),
    .B(_1843_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5406_ (.A1(_1880_),
    .A2(_1965_),
    .B1(_1971_),
    .B2(_1974_),
    .C(_1660_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5407_ (.I0(\registers[28][21] ),
    .I1(\registers[29][21] ),
    .I2(\registers[30][21] ),
    .I3(\registers[31][21] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5408_ (.I0(\registers[24][21] ),
    .I1(\registers[25][21] ),
    .I2(\registers[26][21] ),
    .I3(\registers[27][21] ),
    .S0(_1743_),
    .S1(_1792_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5409_ (.I0(_1976_),
    .I1(_1977_),
    .S(_1902_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5410_ (.I0(\registers[16][21] ),
    .I1(\registers[17][21] ),
    .S(_1795_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5411_ (.I0(\registers[18][21] ),
    .I1(\registers[19][21] ),
    .S(_1797_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5412_ (.I0(\registers[20][21] ),
    .I1(\registers[21][21] ),
    .S(_1748_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5413_ (.I0(\registers[22][21] ),
    .I1(\registers[23][21] ),
    .S(_1800_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5414_ (.I0(_1979_),
    .I1(_1980_),
    .I2(_1981_),
    .I3(_1982_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5415_ (.A1(_1663_),
    .A2(_1978_),
    .B1(_1983_),
    .B2(_1668_),
    .C(_1909_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5416_ (.A1(net61),
    .A2(_1911_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5417_ (.A1(_1975_),
    .A2(_1984_),
    .B(_1985_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5418_ (.I(_1581_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5419_ (.I0(\registers[12][22] ),
    .I1(\registers[13][22] ),
    .I2(\registers[14][22] ),
    .I3(\registers[15][22] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5420_ (.I0(\registers[8][22] ),
    .I1(\registers[9][22] ),
    .I2(\registers[10][22] ),
    .I3(\registers[11][22] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5421_ (.I0(_1987_),
    .I1(_1988_),
    .S(_1831_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5422_ (.I0(\registers[2][22] ),
    .I1(\registers[3][22] ),
    .S(_1886_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5423_ (.I(_1990_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5424_ (.I0(\registers[0][22] ),
    .I1(\registers[1][22] ),
    .S(_1835_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5425_ (.I0(\registers[6][22] ),
    .I1(\registers[7][22] ),
    .S(_1811_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5426_ (.A1(_1889_),
    .A2(_1992_),
    .B1(_1993_),
    .B2(_1892_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5427_ (.A1(_1885_),
    .A2(_1991_),
    .B(_1994_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5428_ (.I0(\registers[4][22] ),
    .I1(\registers[5][22] ),
    .S(_1840_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5429_ (.I(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5430_ (.A1(_1895_),
    .A2(_1997_),
    .B(_1843_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5431_ (.I(net3),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5432_ (.A1(_1880_),
    .A2(_1989_),
    .B1(_1995_),
    .B2(_1998_),
    .C(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5433_ (.I(_1662_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5434_ (.I0(\registers[28][22] ),
    .I1(\registers[29][22] ),
    .I2(\registers[30][22] ),
    .I3(\registers[31][22] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5435_ (.I(_1579_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5436_ (.I0(\registers[24][22] ),
    .I1(\registers[25][22] ),
    .I2(\registers[26][22] ),
    .I3(\registers[27][22] ),
    .S0(_2003_),
    .S1(_1792_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5437_ (.I0(_2002_),
    .I1(_2004_),
    .S(_1902_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5438_ (.I0(\registers[16][22] ),
    .I1(\registers[17][22] ),
    .S(_1795_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5439_ (.I0(\registers[18][22] ),
    .I1(\registers[19][22] ),
    .S(_1797_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5440_ (.I(_1578_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5441_ (.I0(\registers[20][22] ),
    .I1(\registers[21][22] ),
    .S(_2008_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5442_ (.I0(\registers[22][22] ),
    .I1(\registers[23][22] ),
    .S(_1800_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5443_ (.I0(_2006_),
    .I1(_2007_),
    .I2(_2009_),
    .I3(_2010_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5444_ (.I(_1667_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5445_ (.A1(_2001_),
    .A2(_2005_),
    .B1(_2011_),
    .B2(_2012_),
    .C(_1909_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5446_ (.A1(net62),
    .A2(_1911_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5447_ (.A1(_2000_),
    .A2(_2013_),
    .B(_2014_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5448_ (.I0(\registers[12][23] ),
    .I1(\registers[13][23] ),
    .I2(\registers[14][23] ),
    .I3(\registers[15][23] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5449_ (.I0(\registers[8][23] ),
    .I1(\registers[9][23] ),
    .I2(\registers[10][23] ),
    .I3(\registers[11][23] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5450_ (.I0(_2015_),
    .I1(_2016_),
    .S(_1831_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5451_ (.I0(\registers[2][23] ),
    .I1(\registers[3][23] ),
    .S(_1886_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5452_ (.I(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5453_ (.I0(\registers[0][23] ),
    .I1(\registers[1][23] ),
    .S(_1835_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5454_ (.I0(\registers[6][23] ),
    .I1(\registers[7][23] ),
    .S(_1811_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5455_ (.A1(_1889_),
    .A2(_2020_),
    .B1(_2021_),
    .B2(_1892_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5456_ (.A1(_1885_),
    .A2(_2019_),
    .B(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5457_ (.I0(\registers[4][23] ),
    .I1(\registers[5][23] ),
    .S(_1840_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5458_ (.I(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5459_ (.A1(_1895_),
    .A2(_2025_),
    .B(_1843_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5460_ (.A1(_1880_),
    .A2(_2017_),
    .B1(_2023_),
    .B2(_2026_),
    .C(_1999_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5461_ (.I0(\registers[28][23] ),
    .I1(\registers[29][23] ),
    .I2(\registers[30][23] ),
    .I3(\registers[31][23] ),
    .S0(_1790_),
    .S1(_1846_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5462_ (.I0(\registers[24][23] ),
    .I1(\registers[25][23] ),
    .I2(\registers[26][23] ),
    .I3(\registers[27][23] ),
    .S0(_2003_),
    .S1(_1792_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5463_ (.I0(_2028_),
    .I1(_2029_),
    .S(_1902_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5464_ (.I0(\registers[16][23] ),
    .I1(\registers[17][23] ),
    .S(_1795_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5465_ (.I0(\registers[18][23] ),
    .I1(\registers[19][23] ),
    .S(_1797_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5466_ (.I0(\registers[20][23] ),
    .I1(\registers[21][23] ),
    .S(_2008_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5467_ (.I0(\registers[22][23] ),
    .I1(\registers[23][23] ),
    .S(_1800_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5468_ (.I0(_2031_),
    .I1(_2032_),
    .I2(_2033_),
    .I3(_2034_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5469_ (.A1(_2001_),
    .A2(_2030_),
    .B1(_2035_),
    .B2(_2012_),
    .C(_1909_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5470_ (.A1(net63),
    .A2(_1911_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5471_ (.A1(_2027_),
    .A2(_2036_),
    .B(_2037_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5472_ (.I0(\registers[12][24] ),
    .I1(\registers[13][24] ),
    .I2(\registers[14][24] ),
    .I3(\registers[15][24] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5473_ (.I0(\registers[8][24] ),
    .I1(\registers[9][24] ),
    .I2(\registers[10][24] ),
    .I3(\registers[11][24] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5474_ (.I0(_2038_),
    .I1(_2039_),
    .S(_1831_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5475_ (.I0(\registers[2][24] ),
    .I1(\registers[3][24] ),
    .S(_1886_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5476_ (.I(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5477_ (.I0(\registers[0][24] ),
    .I1(\registers[1][24] ),
    .S(_1835_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5478_ (.I0(\registers[6][24] ),
    .I1(\registers[7][24] ),
    .S(_1811_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5479_ (.A1(_1889_),
    .A2(_2043_),
    .B1(_2044_),
    .B2(_1892_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5480_ (.A1(_1885_),
    .A2(_2042_),
    .B(_2045_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5481_ (.I0(\registers[4][24] ),
    .I1(\registers[5][24] ),
    .S(_1840_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5482_ (.I(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5483_ (.A1(_1895_),
    .A2(_2048_),
    .B(_1843_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _5484_ (.A1(_1880_),
    .A2(_2040_),
    .B1(_2046_),
    .B2(_2049_),
    .C(_1999_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5485_ (.I(_1579_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5486_ (.I0(\registers[28][24] ),
    .I1(\registers[29][24] ),
    .I2(\registers[30][24] ),
    .I3(\registers[31][24] ),
    .S0(_2051_),
    .S1(_1846_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5487_ (.I(_1581_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5488_ (.I0(\registers[24][24] ),
    .I1(\registers[25][24] ),
    .I2(\registers[26][24] ),
    .I3(\registers[27][24] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5489_ (.I0(_2052_),
    .I1(_2054_),
    .S(_1902_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5490_ (.I(_1633_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5491_ (.I0(\registers[16][24] ),
    .I1(\registers[17][24] ),
    .S(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5492_ (.I(_1633_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5493_ (.I0(\registers[18][24] ),
    .I1(\registers[19][24] ),
    .S(_2058_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5494_ (.I0(\registers[20][24] ),
    .I1(\registers[21][24] ),
    .S(_2008_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5495_ (.I(_1633_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5496_ (.I0(\registers[22][24] ),
    .I1(\registers[23][24] ),
    .S(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5497_ (.I0(_2057_),
    .I1(_2059_),
    .I2(_2060_),
    .I3(_2062_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5498_ (.A1(_2001_),
    .A2(_2055_),
    .B1(_2063_),
    .B2(_2012_),
    .C(_1909_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5499_ (.A1(net64),
    .A2(_1911_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5500_ (.A1(_2050_),
    .A2(_2064_),
    .B(_2065_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5501_ (.I0(\registers[12][25] ),
    .I1(\registers[13][25] ),
    .I2(\registers[14][25] ),
    .I3(\registers[15][25] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5502_ (.I0(\registers[8][25] ),
    .I1(\registers[9][25] ),
    .I2(\registers[10][25] ),
    .I3(\registers[11][25] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5503_ (.I0(_2066_),
    .I1(_2067_),
    .S(_1831_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5504_ (.I0(\registers[2][25] ),
    .I1(\registers[3][25] ),
    .S(_1886_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5505_ (.I(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5506_ (.I0(\registers[0][25] ),
    .I1(\registers[1][25] ),
    .S(_1835_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5507_ (.I(_1584_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5508_ (.I0(\registers[6][25] ),
    .I1(\registers[7][25] ),
    .S(_2072_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5509_ (.A1(_1889_),
    .A2(_2071_),
    .B1(_2073_),
    .B2(_1892_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5510_ (.A1(_1885_),
    .A2(_2070_),
    .B(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5511_ (.I0(\registers[4][25] ),
    .I1(\registers[5][25] ),
    .S(_1840_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5512_ (.I(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5513_ (.A1(_1895_),
    .A2(_2077_),
    .B(_1843_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _5514_ (.A1(_1880_),
    .A2(_2068_),
    .B1(_2075_),
    .B2(_2078_),
    .C(_1999_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5515_ (.I0(\registers[28][25] ),
    .I1(\registers[29][25] ),
    .I2(\registers[30][25] ),
    .I3(\registers[31][25] ),
    .S0(_2051_),
    .S1(_1846_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5516_ (.I0(\registers[24][25] ),
    .I1(\registers[25][25] ),
    .I2(\registers[26][25] ),
    .I3(\registers[27][25] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5517_ (.I0(_2080_),
    .I1(_2081_),
    .S(_1902_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5518_ (.I0(\registers[16][25] ),
    .I1(\registers[17][25] ),
    .S(_2056_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5519_ (.I0(\registers[18][25] ),
    .I1(\registers[19][25] ),
    .S(_2058_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5520_ (.I0(\registers[20][25] ),
    .I1(\registers[21][25] ),
    .S(_2008_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5521_ (.I0(\registers[22][25] ),
    .I1(\registers[23][25] ),
    .S(_2061_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5522_ (.I0(_2083_),
    .I1(_2084_),
    .I2(_2085_),
    .I3(_2086_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5523_ (.A1(_2001_),
    .A2(_2082_),
    .B1(_2087_),
    .B2(_2012_),
    .C(_1909_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5524_ (.A1(net65),
    .A2(_1911_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5525_ (.A1(_2079_),
    .A2(_2088_),
    .B(_2089_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5526_ (.I0(\registers[28][26] ),
    .I1(\registers[29][26] ),
    .I2(\registers[30][26] ),
    .I3(\registers[31][26] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5527_ (.I0(\registers[24][26] ),
    .I1(\registers[25][26] ),
    .I2(\registers[26][26] ),
    .I3(\registers[27][26] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5528_ (.I(_1589_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5529_ (.I0(_2090_),
    .I1(_2091_),
    .S(_2092_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5530_ (.I0(\registers[18][26] ),
    .I1(\registers[19][26] ),
    .S(_1886_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5531_ (.I(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5532_ (.I(_1584_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5533_ (.I0(\registers[16][26] ),
    .I1(\registers[17][26] ),
    .S(_2096_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5534_ (.I0(\registers[22][26] ),
    .I1(\registers[23][26] ),
    .S(_2072_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5535_ (.A1(_1889_),
    .A2(_2097_),
    .B1(_2098_),
    .B2(_1892_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5536_ (.A1(_1885_),
    .A2(_2095_),
    .B(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5537_ (.I(_1595_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5538_ (.I0(\registers[20][26] ),
    .I1(\registers[21][26] ),
    .S(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5539_ (.I(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5540_ (.I(net2),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5541_ (.A1(_1895_),
    .A2(_2103_),
    .B(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5542_ (.A1(_1880_),
    .A2(_2093_),
    .B1(_2100_),
    .B2(_2105_),
    .C(_1617_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5543_ (.I(_1592_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5544_ (.I0(\registers[12][26] ),
    .I1(\registers[13][26] ),
    .I2(\registers[14][26] ),
    .I3(\registers[15][26] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5545_ (.I0(\registers[8][26] ),
    .I1(\registers[9][26] ),
    .I2(\registers[10][26] ),
    .I3(\registers[11][26] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5546_ (.I0(_2108_),
    .I1(_2109_),
    .S(_1902_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5547_ (.I0(\registers[0][26] ),
    .I1(\registers[1][26] ),
    .S(_2056_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5548_ (.I0(\registers[2][26] ),
    .I1(\registers[3][26] ),
    .S(_2058_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5549_ (.I0(\registers[4][26] ),
    .I1(\registers[5][26] ),
    .S(_2008_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5550_ (.I0(\registers[6][26] ),
    .I1(\registers[7][26] ),
    .S(_2061_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5551_ (.I0(_2111_),
    .I1(_2112_),
    .I2(_2113_),
    .I3(_2114_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5552_ (.A1(_1620_),
    .A2(_2110_),
    .B1(_2115_),
    .B2(_1630_),
    .C(_1909_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5553_ (.A1(net66),
    .A2(_1911_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5554_ (.A1(_2106_),
    .A2(_2116_),
    .B(_2117_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5555_ (.I0(\registers[12][27] ),
    .I1(\registers[13][27] ),
    .I2(\registers[14][27] ),
    .I3(\registers[15][27] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5556_ (.I0(\registers[8][27] ),
    .I1(\registers[9][27] ),
    .I2(\registers[10][27] ),
    .I3(\registers[11][27] ),
    .S0(_1882_),
    .S1(_1938_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5557_ (.I0(_2118_),
    .I1(_2119_),
    .S(_2092_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5558_ (.I0(\registers[2][27] ),
    .I1(\registers[3][27] ),
    .S(_1886_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5559_ (.I(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5560_ (.I0(\registers[0][27] ),
    .I1(\registers[1][27] ),
    .S(_2096_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5561_ (.I0(\registers[6][27] ),
    .I1(\registers[7][27] ),
    .S(_2072_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5562_ (.A1(_1889_),
    .A2(_2123_),
    .B1(_2124_),
    .B2(_1892_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5563_ (.A1(_1885_),
    .A2(_2122_),
    .B(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5564_ (.I0(\registers[4][27] ),
    .I1(\registers[5][27] ),
    .S(_2101_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5565_ (.I(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5566_ (.A1(_1895_),
    .A2(_2128_),
    .B(_2104_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _5567_ (.A1(_1880_),
    .A2(_2120_),
    .B1(_2126_),
    .B2(_2129_),
    .C(_1999_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5568_ (.I0(\registers[28][27] ),
    .I1(\registers[29][27] ),
    .I2(\registers[30][27] ),
    .I3(\registers[31][27] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5569_ (.I0(\registers[24][27] ),
    .I1(\registers[25][27] ),
    .I2(\registers[26][27] ),
    .I3(\registers[27][27] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5570_ (.I0(_2131_),
    .I1(_2132_),
    .S(_1902_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5571_ (.I0(\registers[16][27] ),
    .I1(\registers[17][27] ),
    .S(_2056_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5572_ (.I0(\registers[18][27] ),
    .I1(\registers[19][27] ),
    .S(_2058_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5573_ (.I0(\registers[20][27] ),
    .I1(\registers[21][27] ),
    .S(_2008_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5574_ (.I0(\registers[22][27] ),
    .I1(\registers[23][27] ),
    .S(_2061_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5575_ (.I0(_2134_),
    .I1(_2135_),
    .I2(_2136_),
    .I3(_2137_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5576_ (.A1(_2001_),
    .A2(_2133_),
    .B1(_2138_),
    .B2(_2012_),
    .C(_1909_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5577_ (.A1(net67),
    .A2(_1911_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5578_ (.A1(_2130_),
    .A2(_2139_),
    .B(_2140_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5579_ (.I(_1576_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5580_ (.I0(\registers[12][28] ),
    .I1(\registers[13][28] ),
    .I2(\registers[14][28] ),
    .I3(\registers[15][28] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5581_ (.I(_1584_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5582_ (.I0(\registers[8][28] ),
    .I1(\registers[9][28] ),
    .I2(\registers[10][28] ),
    .I3(\registers[11][28] ),
    .S0(_2143_),
    .S1(_1938_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5583_ (.I0(_2142_),
    .I1(_2144_),
    .S(_2092_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5584_ (.I(_1593_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5585_ (.I(_1595_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5586_ (.I0(\registers[2][28] ),
    .I1(\registers[3][28] ),
    .S(_2147_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5587_ (.I(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5588_ (.I(_1599_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5589_ (.I0(\registers[0][28] ),
    .I1(\registers[1][28] ),
    .S(_2096_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5590_ (.I0(\registers[6][28] ),
    .I1(\registers[7][28] ),
    .S(_2072_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5591_ (.I(_1603_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5592_ (.A1(_2150_),
    .A2(_2151_),
    .B1(_2152_),
    .B2(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5593_ (.A1(_2146_),
    .A2(_2149_),
    .B(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5594_ (.I(_1609_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5595_ (.I0(\registers[4][28] ),
    .I1(\registers[5][28] ),
    .S(_2101_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5596_ (.I(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5597_ (.A1(_2156_),
    .A2(_2158_),
    .B(_2104_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _5598_ (.A1(_2141_),
    .A2(_2145_),
    .B1(_2155_),
    .B2(_2159_),
    .C(_1999_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5599_ (.I0(\registers[28][28] ),
    .I1(\registers[29][28] ),
    .I2(\registers[30][28] ),
    .I3(\registers[31][28] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5600_ (.I0(\registers[24][28] ),
    .I1(\registers[25][28] ),
    .I2(\registers[26][28] ),
    .I3(\registers[27][28] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5601_ (.I(_1589_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5602_ (.I0(_2161_),
    .I1(_2162_),
    .S(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5603_ (.I0(\registers[16][28] ),
    .I1(\registers[17][28] ),
    .S(_2056_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5604_ (.I0(\registers[18][28] ),
    .I1(\registers[19][28] ),
    .S(_2058_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5605_ (.I0(\registers[20][28] ),
    .I1(\registers[21][28] ),
    .S(_2008_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5606_ (.I0(\registers[22][28] ),
    .I1(\registers[23][28] ),
    .S(_2061_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5607_ (.I0(_2165_),
    .I1(_2166_),
    .I2(_2167_),
    .I3(_2168_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5608_ (.I(_1640_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5609_ (.A1(_2001_),
    .A2(_2164_),
    .B1(_2169_),
    .B2(_2012_),
    .C(_2170_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5610_ (.I(_1644_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5611_ (.A1(net68),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5612_ (.A1(_2160_),
    .A2(_2171_),
    .B(_2173_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5613_ (.I0(\registers[28][29] ),
    .I1(\registers[29][29] ),
    .I2(\registers[30][29] ),
    .I3(\registers[31][29] ),
    .S0(_1936_),
    .S1(_1986_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5614_ (.I0(\registers[24][29] ),
    .I1(\registers[25][29] ),
    .I2(\registers[26][29] ),
    .I3(\registers[27][29] ),
    .S0(_2143_),
    .S1(_1938_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5615_ (.I0(_2174_),
    .I1(_2175_),
    .S(_2092_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5616_ (.I0(\registers[18][29] ),
    .I1(\registers[19][29] ),
    .S(_2147_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5617_ (.I(_2177_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5618_ (.I0(\registers[16][29] ),
    .I1(\registers[17][29] ),
    .S(_2096_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5619_ (.I0(\registers[22][29] ),
    .I1(\registers[23][29] ),
    .S(_2072_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5620_ (.A1(_2150_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(_2153_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5621_ (.A1(_2146_),
    .A2(_2178_),
    .B(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5622_ (.I0(\registers[20][29] ),
    .I1(\registers[21][29] ),
    .S(_2101_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5623_ (.I(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5624_ (.A1(_2156_),
    .A2(_2184_),
    .B(_2104_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5625_ (.A1(_2141_),
    .A2(_2176_),
    .B1(_2182_),
    .B2(_2185_),
    .C(_1617_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5626_ (.I0(\registers[12][29] ),
    .I1(\registers[13][29] ),
    .I2(\registers[14][29] ),
    .I3(\registers[15][29] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5627_ (.I0(\registers[8][29] ),
    .I1(\registers[9][29] ),
    .I2(\registers[10][29] ),
    .I3(\registers[11][29] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5628_ (.I0(_2187_),
    .I1(_2188_),
    .S(_2163_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5629_ (.I0(\registers[0][29] ),
    .I1(\registers[1][29] ),
    .S(_2056_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5630_ (.I0(\registers[2][29] ),
    .I1(\registers[3][29] ),
    .S(_2058_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5631_ (.I0(\registers[4][29] ),
    .I1(\registers[5][29] ),
    .S(_2008_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5632_ (.I0(\registers[6][29] ),
    .I1(\registers[7][29] ),
    .S(_2061_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5633_ (.I0(_2190_),
    .I1(_2191_),
    .I2(_2192_),
    .I3(_2193_),
    .S0(_1958_),
    .S1(_1959_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5634_ (.A1(_1620_),
    .A2(_2189_),
    .B1(_2194_),
    .B2(_1630_),
    .C(_2170_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5635_ (.A1(net69),
    .A2(_2172_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5636_ (.A1(_2186_),
    .A2(_2195_),
    .B(_2196_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5637_ (.I(_1579_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5638_ (.I0(\registers[28][2] ),
    .I1(\registers[29][2] ),
    .I2(\registers[30][2] ),
    .I3(\registers[31][2] ),
    .S0(_2197_),
    .S1(_1986_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5639_ (.I(_1581_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5640_ (.I0(\registers[24][2] ),
    .I1(\registers[25][2] ),
    .I2(\registers[26][2] ),
    .I3(\registers[27][2] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5641_ (.I0(_2198_),
    .I1(_2200_),
    .S(_2092_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5642_ (.I0(\registers[18][2] ),
    .I1(\registers[19][2] ),
    .S(_2147_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5643_ (.I(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5644_ (.I0(\registers[16][2] ),
    .I1(\registers[17][2] ),
    .S(_2096_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5645_ (.I0(\registers[22][2] ),
    .I1(\registers[23][2] ),
    .S(_2072_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5646_ (.A1(_2150_),
    .A2(_2204_),
    .B1(_2205_),
    .B2(_2153_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5647_ (.A1(_2146_),
    .A2(_2203_),
    .B(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5648_ (.I0(\registers[20][2] ),
    .I1(\registers[21][2] ),
    .S(_2101_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5649_ (.I(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5650_ (.A1(_2156_),
    .A2(_2209_),
    .B(_2104_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5651_ (.A1(_2141_),
    .A2(_2201_),
    .B1(_2207_),
    .B2(_2210_),
    .C(_1617_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5652_ (.I0(\registers[12][2] ),
    .I1(\registers[13][2] ),
    .I2(\registers[14][2] ),
    .I3(\registers[15][2] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5653_ (.I0(\registers[8][2] ),
    .I1(\registers[9][2] ),
    .I2(\registers[10][2] ),
    .I3(\registers[11][2] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5654_ (.I0(_2212_),
    .I1(_2213_),
    .S(_2163_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5655_ (.I0(\registers[0][2] ),
    .I1(\registers[1][2] ),
    .S(_2056_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5656_ (.I0(\registers[2][2] ),
    .I1(\registers[3][2] ),
    .S(_2058_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5657_ (.I0(\registers[4][2] ),
    .I1(\registers[5][2] ),
    .S(_2008_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5658_ (.I0(\registers[6][2] ),
    .I1(\registers[7][2] ),
    .S(_2061_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5659_ (.I(_1592_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5660_ (.I(net1),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5661_ (.I0(_2215_),
    .I1(_2216_),
    .I2(_2217_),
    .I3(_2218_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5662_ (.A1(_1620_),
    .A2(_2214_),
    .B1(_2221_),
    .B2(_1630_),
    .C(_2170_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5663_ (.A1(net70),
    .A2(_2172_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5664_ (.A1(_2211_),
    .A2(_2222_),
    .B(_2223_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5665_ (.I0(\registers[12][30] ),
    .I1(\registers[13][30] ),
    .I2(\registers[14][30] ),
    .I3(\registers[15][30] ),
    .S0(_2197_),
    .S1(_1986_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5666_ (.I0(\registers[8][30] ),
    .I1(\registers[9][30] ),
    .I2(\registers[10][30] ),
    .I3(\registers[11][30] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5667_ (.I0(_2224_),
    .I1(_2225_),
    .S(_2092_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5668_ (.I0(\registers[2][30] ),
    .I1(\registers[3][30] ),
    .S(_2147_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5669_ (.I(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5670_ (.I0(\registers[0][30] ),
    .I1(\registers[1][30] ),
    .S(_2096_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5671_ (.I0(\registers[6][30] ),
    .I1(\registers[7][30] ),
    .S(_2072_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5672_ (.A1(_2150_),
    .A2(_2229_),
    .B1(_2230_),
    .B2(_2153_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5673_ (.A1(_2146_),
    .A2(_2228_),
    .B(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5674_ (.I0(\registers[4][30] ),
    .I1(\registers[5][30] ),
    .S(_2101_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5675_ (.I(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5676_ (.A1(_2156_),
    .A2(_2234_),
    .B(_2104_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _5677_ (.A1(_2141_),
    .A2(_2226_),
    .B1(_2232_),
    .B2(_2235_),
    .C(_1999_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5678_ (.I0(\registers[28][30] ),
    .I1(\registers[29][30] ),
    .I2(\registers[30][30] ),
    .I3(\registers[31][30] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5679_ (.I0(\registers[24][30] ),
    .I1(\registers[25][30] ),
    .I2(\registers[26][30] ),
    .I3(\registers[27][30] ),
    .S0(_2003_),
    .S1(_2053_),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5680_ (.I0(_2237_),
    .I1(_2238_),
    .S(_2163_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5681_ (.I0(\registers[16][30] ),
    .I1(\registers[17][30] ),
    .S(_2056_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5682_ (.I0(\registers[18][30] ),
    .I1(\registers[19][30] ),
    .S(_2058_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5683_ (.I0(\registers[20][30] ),
    .I1(\registers[21][30] ),
    .S(_2008_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5684_ (.I0(\registers[22][30] ),
    .I1(\registers[23][30] ),
    .S(_2061_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5685_ (.I0(_2240_),
    .I1(_2241_),
    .I2(_2242_),
    .I3(_2243_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5686_ (.A1(_2001_),
    .A2(_2239_),
    .B1(_2244_),
    .B2(_2012_),
    .C(_2170_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5687_ (.A1(net71),
    .A2(_2172_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5688_ (.A1(_2236_),
    .A2(_2245_),
    .B(_2246_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5689_ (.I0(\registers[12][31] ),
    .I1(\registers[13][31] ),
    .I2(\registers[14][31] ),
    .I3(\registers[15][31] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5690_ (.I0(\registers[8][31] ),
    .I1(\registers[9][31] ),
    .I2(\registers[10][31] ),
    .I3(\registers[11][31] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5691_ (.I0(_2247_),
    .I1(_2248_),
    .S(_2092_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5692_ (.I0(\registers[2][31] ),
    .I1(\registers[3][31] ),
    .S(_2147_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5693_ (.I(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5694_ (.I0(\registers[0][31] ),
    .I1(\registers[1][31] ),
    .S(_2096_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5695_ (.I0(\registers[6][31] ),
    .I1(\registers[7][31] ),
    .S(_2072_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5696_ (.A1(_2150_),
    .A2(_2252_),
    .B1(_2253_),
    .B2(_2153_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5697_ (.A1(_2146_),
    .A2(_2251_),
    .B(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5698_ (.I0(\registers[4][31] ),
    .I1(\registers[5][31] ),
    .S(_2101_),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5699_ (.I(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5700_ (.A1(_2156_),
    .A2(_2257_),
    .B(_2104_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _5701_ (.A1(_2141_),
    .A2(_2249_),
    .B1(_2255_),
    .B2(_2258_),
    .C(_1999_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5702_ (.I0(\registers[28][31] ),
    .I1(\registers[29][31] ),
    .I2(\registers[30][31] ),
    .I3(\registers[31][31] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5703_ (.I0(\registers[24][31] ),
    .I1(\registers[25][31] ),
    .I2(\registers[26][31] ),
    .I3(\registers[27][31] ),
    .S0(_1580_),
    .S1(_2053_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5704_ (.I0(_2260_),
    .I1(_2261_),
    .S(_2163_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5705_ (.I0(\registers[16][31] ),
    .I1(\registers[17][31] ),
    .S(_2056_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5706_ (.I0(\registers[18][31] ),
    .I1(\registers[19][31] ),
    .S(_2058_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5707_ (.I0(\registers[20][31] ),
    .I1(\registers[21][31] ),
    .S(_1631_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5708_ (.I0(\registers[22][31] ),
    .I1(\registers[23][31] ),
    .S(_2061_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5709_ (.I0(_2263_),
    .I1(_2264_),
    .I2(_2265_),
    .I3(_2266_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5710_ (.A1(_2001_),
    .A2(_2262_),
    .B1(_2267_),
    .B2(_2012_),
    .C(_2170_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5711_ (.A1(net72),
    .A2(_2172_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5712_ (.A1(_2259_),
    .A2(_2268_),
    .B(_2269_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5713_ (.I0(\registers[12][3] ),
    .I1(\registers[13][3] ),
    .I2(\registers[14][3] ),
    .I3(\registers[15][3] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5714_ (.I0(\registers[8][3] ),
    .I1(\registers[9][3] ),
    .I2(\registers[10][3] ),
    .I3(\registers[11][3] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5715_ (.I0(_2270_),
    .I1(_2271_),
    .S(_2092_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5716_ (.I0(\registers[2][3] ),
    .I1(\registers[3][3] ),
    .S(_2147_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5717_ (.I(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5718_ (.I0(\registers[0][3] ),
    .I1(\registers[1][3] ),
    .S(_2096_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5719_ (.I0(\registers[6][3] ),
    .I1(\registers[7][3] ),
    .S(_2072_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5720_ (.A1(_2150_),
    .A2(_2275_),
    .B1(_2276_),
    .B2(_2153_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5721_ (.A1(_2146_),
    .A2(_2274_),
    .B(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5722_ (.I0(\registers[4][3] ),
    .I1(\registers[5][3] ),
    .S(_2101_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5723_ (.I(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5724_ (.A1(_2156_),
    .A2(_2280_),
    .B(_2104_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5725_ (.A1(_2141_),
    .A2(_2272_),
    .B1(_2278_),
    .B2(_2281_),
    .C(_1999_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5726_ (.I0(\registers[28][3] ),
    .I1(\registers[29][3] ),
    .I2(\registers[30][3] ),
    .I3(\registers[31][3] ),
    .S0(_2051_),
    .S1(_2107_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5727_ (.I0(\registers[24][3] ),
    .I1(\registers[25][3] ),
    .I2(\registers[26][3] ),
    .I3(\registers[27][3] ),
    .S0(_1580_),
    .S1(_2053_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5728_ (.I0(_2283_),
    .I1(_2284_),
    .S(_2163_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5729_ (.I0(\registers[16][3] ),
    .I1(\registers[17][3] ),
    .S(_2056_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5730_ (.I0(\registers[18][3] ),
    .I1(\registers[19][3] ),
    .S(_2058_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5731_ (.I0(\registers[20][3] ),
    .I1(\registers[21][3] ),
    .S(_1631_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5732_ (.I0(\registers[22][3] ),
    .I1(\registers[23][3] ),
    .S(_2061_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5733_ (.I0(_2286_),
    .I1(_2287_),
    .I2(_2288_),
    .I3(_2289_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5734_ (.A1(_2001_),
    .A2(_2285_),
    .B1(_2290_),
    .B2(_2012_),
    .C(_2170_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5735_ (.A1(net73),
    .A2(_2172_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5736_ (.A1(_2282_),
    .A2(_2291_),
    .B(_2292_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5737_ (.I0(\registers[12][4] ),
    .I1(\registers[13][4] ),
    .I2(\registers[14][4] ),
    .I3(\registers[15][4] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5738_ (.I0(\registers[8][4] ),
    .I1(\registers[9][4] ),
    .I2(\registers[10][4] ),
    .I3(\registers[11][4] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5739_ (.I0(_2293_),
    .I1(_2294_),
    .S(_2092_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5740_ (.I0(\registers[2][4] ),
    .I1(\registers[3][4] ),
    .S(_2147_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5741_ (.I(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5742_ (.I0(\registers[0][4] ),
    .I1(\registers[1][4] ),
    .S(_2096_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5743_ (.I0(\registers[6][4] ),
    .I1(\registers[7][4] ),
    .S(_2072_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5744_ (.A1(_2150_),
    .A2(_2298_),
    .B1(_2299_),
    .B2(_2153_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5745_ (.A1(_2146_),
    .A2(_2297_),
    .B(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5746_ (.I0(\registers[4][4] ),
    .I1(\registers[5][4] ),
    .S(_2101_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5747_ (.I(_2302_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5748_ (.A1(_2156_),
    .A2(_2303_),
    .B(_2104_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5749_ (.A1(_2141_),
    .A2(_2295_),
    .B1(_2301_),
    .B2(_2304_),
    .C(_1999_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5750_ (.I0(\registers[28][4] ),
    .I1(\registers[29][4] ),
    .I2(\registers[30][4] ),
    .I3(\registers[31][4] ),
    .S0(_1624_),
    .S1(_2107_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5751_ (.I0(\registers[24][4] ),
    .I1(\registers[25][4] ),
    .I2(\registers[26][4] ),
    .I3(\registers[27][4] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5752_ (.I0(_2306_),
    .I1(_2307_),
    .S(_2163_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5753_ (.I0(\registers[16][4] ),
    .I1(\registers[17][4] ),
    .S(_1698_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5754_ (.I0(\registers[18][4] ),
    .I1(\registers[19][4] ),
    .S(_1694_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5755_ (.I0(\registers[20][4] ),
    .I1(\registers[21][4] ),
    .S(_1631_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5756_ (.I0(\registers[22][4] ),
    .I1(\registers[23][4] ),
    .S(_1634_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5757_ (.I0(_2309_),
    .I1(_2310_),
    .I2(_2311_),
    .I3(_2312_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5758_ (.A1(_2001_),
    .A2(_2308_),
    .B1(_2313_),
    .B2(_2012_),
    .C(_2170_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5759_ (.A1(net74),
    .A2(_2172_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5760_ (.A1(_2305_),
    .A2(_2314_),
    .B(_2315_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5761_ (.I0(\registers[28][5] ),
    .I1(\registers[29][5] ),
    .I2(\registers[30][5] ),
    .I3(\registers[31][5] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5762_ (.I0(\registers[24][5] ),
    .I1(\registers[25][5] ),
    .I2(\registers[26][5] ),
    .I3(\registers[27][5] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5763_ (.I0(_2316_),
    .I1(_2317_),
    .S(_2092_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5764_ (.I0(\registers[18][5] ),
    .I1(\registers[19][5] ),
    .S(_2147_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5765_ (.I(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5766_ (.I0(\registers[16][5] ),
    .I1(\registers[17][5] ),
    .S(_2096_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5767_ (.I0(\registers[22][5] ),
    .I1(\registers[23][5] ),
    .S(_1605_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5768_ (.A1(_2150_),
    .A2(_2321_),
    .B1(_2322_),
    .B2(_2153_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5769_ (.A1(_2146_),
    .A2(_2320_),
    .B(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5770_ (.I0(\registers[20][5] ),
    .I1(\registers[21][5] ),
    .S(_2101_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5771_ (.I(_2325_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5772_ (.A1(_2156_),
    .A2(_2326_),
    .B(_2104_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5773_ (.A1(_2141_),
    .A2(_2318_),
    .B1(_2324_),
    .B2(_2327_),
    .C(_1617_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5774_ (.I0(\registers[12][5] ),
    .I1(\registers[13][5] ),
    .I2(\registers[14][5] ),
    .I3(\registers[15][5] ),
    .S0(_1624_),
    .S1(_2107_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5775_ (.I0(\registers[8][5] ),
    .I1(\registers[9][5] ),
    .I2(\registers[10][5] ),
    .I3(\registers[11][5] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5776_ (.I0(_2329_),
    .I1(_2330_),
    .S(_2163_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5777_ (.I0(\registers[0][5] ),
    .I1(\registers[1][5] ),
    .S(_1698_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5778_ (.I0(\registers[2][5] ),
    .I1(\registers[3][5] ),
    .S(_1694_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5779_ (.I0(\registers[4][5] ),
    .I1(\registers[5][5] ),
    .S(_1631_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5780_ (.I0(\registers[6][5] ),
    .I1(\registers[7][5] ),
    .S(_1634_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5781_ (.I0(_2332_),
    .I1(_2333_),
    .I2(_2334_),
    .I3(_2335_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5782_ (.A1(_1620_),
    .A2(_2331_),
    .B1(_2336_),
    .B2(_1630_),
    .C(_2170_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5783_ (.A1(net75),
    .A2(_2172_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5784_ (.A1(_2328_),
    .A2(_2337_),
    .B(_2338_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5785_ (.I0(\registers[28][6] ),
    .I1(\registers[29][6] ),
    .I2(\registers[30][6] ),
    .I3(\registers[31][6] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5786_ (.I0(\registers[24][6] ),
    .I1(\registers[25][6] ),
    .I2(\registers[26][6] ),
    .I3(\registers[27][6] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5787_ (.I0(_2339_),
    .I1(_2340_),
    .S(_1589_),
    .Z(_2341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5788_ (.I0(\registers[18][6] ),
    .I1(\registers[19][6] ),
    .S(_2147_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5789_ (.I(_2342_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5790_ (.I0(\registers[16][6] ),
    .I1(\registers[17][6] ),
    .S(_1653_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5791_ (.I0(\registers[22][6] ),
    .I1(\registers[23][6] ),
    .S(_1605_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5792_ (.A1(_2150_),
    .A2(_2344_),
    .B1(_2345_),
    .B2(_2153_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5793_ (.A1(_2146_),
    .A2(_2343_),
    .B(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5794_ (.I0(\registers[20][6] ),
    .I1(\registers[21][6] ),
    .S(_1621_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5795_ (.I(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5796_ (.A1(_2156_),
    .A2(_2349_),
    .B(_1576_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5797_ (.A1(_2141_),
    .A2(_2341_),
    .B1(_2347_),
    .B2(_2350_),
    .C(_1617_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5798_ (.I0(\registers[12][6] ),
    .I1(\registers[13][6] ),
    .I2(\registers[14][6] ),
    .I3(\registers[15][6] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5799_ (.I0(\registers[8][6] ),
    .I1(\registers[9][6] ),
    .I2(\registers[10][6] ),
    .I3(\registers[11][6] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5800_ (.I0(_2352_),
    .I1(_2353_),
    .S(_2163_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5801_ (.I0(\registers[0][6] ),
    .I1(\registers[1][6] ),
    .S(_1698_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5802_ (.I0(\registers[2][6] ),
    .I1(\registers[3][6] ),
    .S(_1694_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5803_ (.I0(\registers[4][6] ),
    .I1(\registers[5][6] ),
    .S(_1631_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5804_ (.I0(\registers[6][6] ),
    .I1(\registers[7][6] ),
    .S(_1634_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5805_ (.I0(_2355_),
    .I1(_2356_),
    .I2(_2357_),
    .I3(_2358_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5806_ (.A1(_1620_),
    .A2(_2354_),
    .B1(_2359_),
    .B2(_1630_),
    .C(_2170_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5807_ (.A1(net76),
    .A2(_2172_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5808_ (.A1(_2351_),
    .A2(_2360_),
    .B(_2361_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5809_ (.I0(\registers[28][7] ),
    .I1(\registers[29][7] ),
    .I2(\registers[30][7] ),
    .I3(\registers[31][7] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5810_ (.I0(\registers[24][7] ),
    .I1(\registers[25][7] ),
    .I2(\registers[26][7] ),
    .I3(\registers[27][7] ),
    .S0(_2143_),
    .S1(_2199_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5811_ (.I0(_2362_),
    .I1(_2363_),
    .S(_1589_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5812_ (.I0(\registers[18][7] ),
    .I1(\registers[19][7] ),
    .S(_2147_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5813_ (.I(_2365_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5814_ (.I0(\registers[16][7] ),
    .I1(\registers[17][7] ),
    .S(_1653_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5815_ (.I0(\registers[22][7] ),
    .I1(\registers[23][7] ),
    .S(_1605_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5816_ (.A1(_2150_),
    .A2(_2367_),
    .B1(_2368_),
    .B2(_2153_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5817_ (.A1(_2146_),
    .A2(_2366_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5818_ (.I0(\registers[20][7] ),
    .I1(\registers[21][7] ),
    .S(_1621_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5819_ (.I(_2371_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5820_ (.A1(_2156_),
    .A2(_2372_),
    .B(_1576_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5821_ (.A1(_2141_),
    .A2(_2364_),
    .B1(_2370_),
    .B2(_2373_),
    .C(_1617_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5822_ (.I0(\registers[12][7] ),
    .I1(\registers[13][7] ),
    .I2(\registers[14][7] ),
    .I3(\registers[15][7] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5823_ (.I0(\registers[8][7] ),
    .I1(\registers[9][7] ),
    .I2(\registers[10][7] ),
    .I3(\registers[11][7] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5824_ (.I0(_2375_),
    .I1(_2376_),
    .S(_2163_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5825_ (.I0(\registers[0][7] ),
    .I1(\registers[1][7] ),
    .S(_1698_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5826_ (.I0(\registers[2][7] ),
    .I1(\registers[3][7] ),
    .S(_1694_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5827_ (.I0(\registers[4][7] ),
    .I1(\registers[5][7] ),
    .S(_1631_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5828_ (.I0(\registers[6][7] ),
    .I1(\registers[7][7] ),
    .S(_1634_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5829_ (.I0(_2378_),
    .I1(_2379_),
    .I2(_2380_),
    .I3(_2381_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5830_ (.A1(_1620_),
    .A2(_2377_),
    .B1(_2382_),
    .B2(_1630_),
    .C(_2170_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5831_ (.A1(net77),
    .A2(_2172_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5832_ (.A1(_2374_),
    .A2(_2383_),
    .B(_2384_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5833_ (.I0(\registers[12][8] ),
    .I1(\registers[13][8] ),
    .I2(\registers[14][8] ),
    .I3(\registers[15][8] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5834_ (.I0(\registers[8][8] ),
    .I1(\registers[9][8] ),
    .I2(\registers[10][8] ),
    .I3(\registers[11][8] ),
    .S0(_1601_),
    .S1(_2199_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5835_ (.I0(_2385_),
    .I1(_2386_),
    .S(_1589_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5836_ (.I0(\registers[2][8] ),
    .I1(\registers[3][8] ),
    .S(_1611_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5837_ (.I(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5838_ (.I0(\registers[0][8] ),
    .I1(\registers[1][8] ),
    .S(_1653_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5839_ (.I0(\registers[6][8] ),
    .I1(\registers[7][8] ),
    .S(_1605_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5840_ (.A1(_1599_),
    .A2(_2390_),
    .B1(_2391_),
    .B2(_1603_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5841_ (.A1(_1593_),
    .A2(_2389_),
    .B(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5842_ (.I0(\registers[4][8] ),
    .I1(\registers[5][8] ),
    .S(_1621_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5843_ (.I(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5844_ (.A1(_1609_),
    .A2(_2395_),
    .B(_1576_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5845_ (.A1(_1614_),
    .A2(_2387_),
    .B1(_2393_),
    .B2(_2396_),
    .C(net3),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5846_ (.I0(\registers[28][8] ),
    .I1(\registers[29][8] ),
    .I2(\registers[30][8] ),
    .I3(\registers[31][8] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_2398_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5847_ (.I0(\registers[24][8] ),
    .I1(\registers[25][8] ),
    .I2(\registers[26][8] ),
    .I3(\registers[27][8] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5848_ (.I0(_2398_),
    .I1(_2399_),
    .S(_1590_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5849_ (.I0(\registers[16][8] ),
    .I1(\registers[17][8] ),
    .S(_1698_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5850_ (.I0(\registers[18][8] ),
    .I1(\registers[19][8] ),
    .S(_1694_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5851_ (.I0(\registers[20][8] ),
    .I1(\registers[21][8] ),
    .S(_1631_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5852_ (.I0(\registers[22][8] ),
    .I1(\registers[23][8] ),
    .S(_1634_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5853_ (.I0(_2401_),
    .I1(_2402_),
    .I2(_2403_),
    .I3(_2404_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5854_ (.A1(_1662_),
    .A2(_2400_),
    .B1(_2405_),
    .B2(_1667_),
    .C(_1640_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5855_ (.A1(net78),
    .A2(_1644_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5856_ (.A1(_2397_),
    .A2(_2406_),
    .B(_2407_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5857_ (.I0(\registers[28][9] ),
    .I1(\registers[29][9] ),
    .I2(\registers[30][9] ),
    .I3(\registers[31][9] ),
    .S0(_2197_),
    .S1(_1586_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5858_ (.I0(\registers[24][9] ),
    .I1(\registers[25][9] ),
    .I2(\registers[26][9] ),
    .I3(\registers[27][9] ),
    .S0(_1601_),
    .S1(_2199_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5859_ (.I0(_2408_),
    .I1(_2409_),
    .S(_1589_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5860_ (.I0(\registers[18][9] ),
    .I1(\registers[19][9] ),
    .S(_1611_),
    .Z(_2411_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5861_ (.I(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5862_ (.I0(\registers[16][9] ),
    .I1(\registers[17][9] ),
    .S(_1653_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5863_ (.I0(\registers[22][9] ),
    .I1(\registers[23][9] ),
    .S(_1605_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5864_ (.A1(_1599_),
    .A2(_2413_),
    .B1(_2414_),
    .B2(_1603_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5865_ (.A1(_1593_),
    .A2(_2412_),
    .B(_2415_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5866_ (.I0(\registers[20][9] ),
    .I1(\registers[21][9] ),
    .S(_1621_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5867_ (.I(_2417_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5868_ (.A1(_1609_),
    .A2(_2418_),
    .B(_1576_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5869_ (.A1(_1614_),
    .A2(_2410_),
    .B1(_2416_),
    .B2(_2419_),
    .C(_1616_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5870_ (.I0(\registers[12][9] ),
    .I1(\registers[13][9] ),
    .I2(\registers[14][9] ),
    .I3(\registers[15][9] ),
    .S0(_1624_),
    .S1(_1625_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5871_ (.I0(\registers[8][9] ),
    .I1(\registers[9][9] ),
    .I2(\registers[10][9] ),
    .I3(\registers[11][9] ),
    .S0(_1580_),
    .S1(_1582_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5872_ (.I0(_2421_),
    .I1(_2422_),
    .S(_1590_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5873_ (.I0(\registers[0][9] ),
    .I1(\registers[1][9] ),
    .S(_1698_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5874_ (.I0(\registers[2][9] ),
    .I1(\registers[3][9] ),
    .S(_1694_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5875_ (.I0(\registers[4][9] ),
    .I1(\registers[5][9] ),
    .S(_1631_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5876_ (.I0(\registers[6][9] ),
    .I1(\registers[7][9] ),
    .S(_1634_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5877_ (.I0(_2424_),
    .I1(_2425_),
    .I2(_2426_),
    .I3(_2427_),
    .S0(_2219_),
    .S1(_2220_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5878_ (.A1(_1619_),
    .A2(_2423_),
    .B1(_2428_),
    .B2(_1629_),
    .C(_1640_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5879_ (.A1(net79),
    .A2(_1644_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5880_ (.A1(_2420_),
    .A2(_2429_),
    .B(_2430_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5881_ (.I(net5),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5882_ (.I(_2431_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5883_ (.I(read_addr2[0]),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _5884_ (.I(_2433_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5885_ (.I(_2434_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5886_ (.I(read_addr2[1]),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5887_ (.I(_2436_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5888_ (.I0(\registers[28][0] ),
    .I1(\registers[29][0] ),
    .I2(\registers[30][0] ),
    .I3(\registers[31][0] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5889_ (.I(_2433_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5890_ (.I(_2439_),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5891_ (.I(_2436_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5892_ (.I0(\registers[24][0] ),
    .I1(\registers[25][0] ),
    .I2(\registers[26][0] ),
    .I3(\registers[27][0] ),
    .S0(_2440_),
    .S1(_2441_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _5893_ (.I(net4),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _5894_ (.I(_2443_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5895_ (.I(_2444_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5896_ (.I0(_2438_),
    .I1(_2442_),
    .S(_2445_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5897_ (.I(read_addr2[1]),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5898_ (.A1(_2447_),
    .A2(_2443_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5899_ (.I(_2448_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5900_ (.I(_2433_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5901_ (.I(_2450_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5902_ (.I0(\registers[18][0] ),
    .I1(\registers[19][0] ),
    .S(_2451_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5903_ (.I(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _5904_ (.A1(_2436_),
    .A2(net4),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5905_ (.I(_2454_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5906_ (.I(_2439_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5907_ (.I0(\registers[16][0] ),
    .I1(\registers[17][0] ),
    .S(_2456_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _5908_ (.A1(_2436_),
    .A2(net4),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5909_ (.I(_2458_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5910_ (.I(_2439_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5911_ (.I0(\registers[22][0] ),
    .I1(\registers[23][0] ),
    .S(_2460_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5912_ (.A1(_2455_),
    .A2(_2457_),
    .B1(_2459_),
    .B2(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5913_ (.A1(_2449_),
    .A2(_2453_),
    .B(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _5914_ (.A1(_2447_),
    .A2(_2443_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5915_ (.I(_2464_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5916_ (.I(_2450_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5917_ (.I0(\registers[20][0] ),
    .I1(\registers[21][0] ),
    .S(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5918_ (.I(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5919_ (.I(net5),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5920_ (.A1(_2465_),
    .A2(_2468_),
    .B(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _5921_ (.I(net6),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5922_ (.I(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5923_ (.A1(_2432_),
    .A2(_2446_),
    .B1(_2463_),
    .B2(_2470_),
    .C(_2472_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _5924_ (.A1(_2431_),
    .A2(_2471_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5925_ (.I(_2474_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5926_ (.I(_2434_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5927_ (.I(_2447_),
    .Z(_2477_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5928_ (.I0(\registers[12][0] ),
    .I1(\registers[13][0] ),
    .I2(\registers[14][0] ),
    .I3(\registers[15][0] ),
    .S0(_2476_),
    .S1(_2477_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5929_ (.I(_2434_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5930_ (.I(_2447_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5931_ (.I0(\registers[8][0] ),
    .I1(\registers[9][0] ),
    .I2(\registers[10][0] ),
    .I3(\registers[11][0] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5932_ (.I(_2444_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5933_ (.I0(_2478_),
    .I1(_2481_),
    .S(_2482_),
    .Z(_2483_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5934_ (.A1(net5),
    .A2(net6),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5935_ (.I(_2484_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5936_ (.I(_2433_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5937_ (.I0(\registers[0][0] ),
    .I1(\registers[1][0] ),
    .S(_2486_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 _5938_ (.I(_2433_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5939_ (.I(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5940_ (.I0(\registers[2][0] ),
    .I1(\registers[3][0] ),
    .S(_2489_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5941_ (.I0(\registers[4][0] ),
    .I1(\registers[5][0] ),
    .S(_2450_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5942_ (.I0(\registers[6][0] ),
    .I1(\registers[7][0] ),
    .S(_2450_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5943_ (.I0(_2487_),
    .I1(_2490_),
    .I2(_2491_),
    .I3(_2492_),
    .S0(_2477_),
    .S1(net4),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5944_ (.A1(_1639_),
    .A2(net8),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5945_ (.I(_2494_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5946_ (.A1(_2475_),
    .A2(_2483_),
    .B1(_2485_),
    .B2(_2493_),
    .C(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5947_ (.I(net8),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _5948_ (.A1(_1639_),
    .A2(_2497_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5949_ (.I(_2498_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5950_ (.A1(net80),
    .A2(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5951_ (.A1(_2473_),
    .A2(_2496_),
    .B(_2500_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5952_ (.I0(\registers[12][10] ),
    .I1(\registers[13][10] ),
    .I2(\registers[14][10] ),
    .I3(\registers[15][10] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5953_ (.I0(\registers[8][10] ),
    .I1(\registers[9][10] ),
    .I2(\registers[10][10] ),
    .I3(\registers[11][10] ),
    .S0(_2440_),
    .S1(_2441_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5954_ (.I0(_2501_),
    .I1(_2502_),
    .S(_2445_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5955_ (.I0(\registers[2][10] ),
    .I1(\registers[3][10] ),
    .S(_2451_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5956_ (.I(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5957_ (.I0(\registers[0][10] ),
    .I1(\registers[1][10] ),
    .S(_2456_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5958_ (.I(_2439_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5959_ (.I0(\registers[6][10] ),
    .I1(\registers[7][10] ),
    .S(_2507_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5960_ (.A1(_2455_),
    .A2(_2506_),
    .B1(_2508_),
    .B2(_2459_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5961_ (.A1(_2449_),
    .A2(_2505_),
    .B(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5962_ (.I0(\registers[4][10] ),
    .I1(\registers[5][10] ),
    .S(_2466_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5963_ (.I(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5964_ (.A1(_2465_),
    .A2(_2512_),
    .B(_2469_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5965_ (.I(net6),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5966_ (.A1(_2432_),
    .A2(_2503_),
    .B1(_2510_),
    .B2(_2513_),
    .C(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5967_ (.A1(_2431_),
    .A2(net6),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5968_ (.I(_2516_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5969_ (.I0(\registers[28][10] ),
    .I1(\registers[29][10] ),
    .I2(\registers[30][10] ),
    .I3(\registers[31][10] ),
    .S0(_2476_),
    .S1(_2477_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5970_ (.I0(\registers[24][10] ),
    .I1(\registers[25][10] ),
    .I2(\registers[26][10] ),
    .I3(\registers[27][10] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5971_ (.I0(_2518_),
    .I1(_2519_),
    .S(_2482_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5972_ (.A1(net5),
    .A2(_2471_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _5973_ (.I(_2521_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5974_ (.I0(\registers[16][10] ),
    .I1(\registers[17][10] ),
    .S(_2486_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5975_ (.I0(\registers[18][10] ),
    .I1(\registers[19][10] ),
    .S(_2489_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5976_ (.I0(\registers[20][10] ),
    .I1(\registers[21][10] ),
    .S(_2450_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5977_ (.I0(\registers[22][10] ),
    .I1(\registers[23][10] ),
    .S(_2450_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5978_ (.I0(_2523_),
    .I1(_2524_),
    .I2(_2525_),
    .I3(_2526_),
    .S0(_2477_),
    .S1(net4),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5979_ (.A1(_2517_),
    .A2(_2520_),
    .B1(_2522_),
    .B2(_2527_),
    .C(_2495_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5980_ (.A1(net81),
    .A2(_2499_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5981_ (.A1(_2515_),
    .A2(_2528_),
    .B(_2529_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _5982_ (.I(_2434_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5983_ (.I0(\registers[12][11] ),
    .I1(\registers[13][11] ),
    .I2(\registers[14][11] ),
    .I3(\registers[15][11] ),
    .S0(_2530_),
    .S1(_2437_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _5984_ (.I(_2436_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5985_ (.I0(\registers[8][11] ),
    .I1(\registers[9][11] ),
    .I2(\registers[10][11] ),
    .I3(\registers[11][11] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5986_ (.I0(_2531_),
    .I1(_2533_),
    .S(_2445_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5987_ (.I0(\registers[2][11] ),
    .I1(\registers[3][11] ),
    .S(_2451_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5988_ (.I(_2535_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5989_ (.I0(\registers[0][11] ),
    .I1(\registers[1][11] ),
    .S(_2456_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5990_ (.I0(\registers[6][11] ),
    .I1(\registers[7][11] ),
    .S(_2507_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _5991_ (.A1(_2455_),
    .A2(_2537_),
    .B1(_2538_),
    .B2(_2459_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5992_ (.A1(_2449_),
    .A2(_2536_),
    .B(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5993_ (.I0(\registers[4][11] ),
    .I1(\registers[5][11] ),
    .S(_2466_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _5994_ (.I(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5995_ (.A1(_2465_),
    .A2(_2542_),
    .B(_2469_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5996_ (.A1(_2432_),
    .A2(_2534_),
    .B1(_2540_),
    .B2(_2543_),
    .C(_2514_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5997_ (.I0(\registers[28][11] ),
    .I1(\registers[29][11] ),
    .I2(\registers[30][11] ),
    .I3(\registers[31][11] ),
    .S0(_2476_),
    .S1(_2477_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _5998_ (.I0(\registers[24][11] ),
    .I1(\registers[25][11] ),
    .I2(\registers[26][11] ),
    .I3(\registers[27][11] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _5999_ (.I0(_2545_),
    .I1(_2546_),
    .S(_2482_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6000_ (.I(_2488_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6001_ (.I0(\registers[16][11] ),
    .I1(\registers[17][11] ),
    .S(_2548_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6002_ (.I0(\registers[18][11] ),
    .I1(\registers[19][11] ),
    .S(_2460_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6003_ (.I0(\registers[20][11] ),
    .I1(\registers[21][11] ),
    .S(_2489_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6004_ (.I(_2488_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6005_ (.I0(\registers[22][11] ),
    .I1(\registers[23][11] ),
    .S(_2552_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6006_ (.I(_2447_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6007_ (.I(net4),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6008_ (.I0(_2549_),
    .I1(_2550_),
    .I2(_2551_),
    .I3(_2553_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2556_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6009_ (.A1(_2517_),
    .A2(_2547_),
    .B1(_2556_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6010_ (.A1(net82),
    .A2(_2499_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6011_ (.A1(_2544_),
    .A2(_2557_),
    .B(_2558_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6012_ (.I0(\registers[12][12] ),
    .I1(\registers[13][12] ),
    .I2(\registers[14][12] ),
    .I3(\registers[15][12] ),
    .S0(_2530_),
    .S1(_2437_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6013_ (.I0(\registers[8][12] ),
    .I1(\registers[9][12] ),
    .I2(\registers[10][12] ),
    .I3(\registers[11][12] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6014_ (.I0(_2559_),
    .I1(_2560_),
    .S(_2445_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6015_ (.I0(\registers[2][12] ),
    .I1(\registers[3][12] ),
    .S(_2451_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6016_ (.I(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6017_ (.I0(\registers[0][12] ),
    .I1(\registers[1][12] ),
    .S(_2456_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6018_ (.I0(\registers[6][12] ),
    .I1(\registers[7][12] ),
    .S(_2507_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6019_ (.A1(_2455_),
    .A2(_2564_),
    .B1(_2565_),
    .B2(_2459_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6020_ (.A1(_2449_),
    .A2(_2563_),
    .B(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6021_ (.I0(\registers[4][12] ),
    .I1(\registers[5][12] ),
    .S(_2466_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6022_ (.I(_2568_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6023_ (.A1(_2465_),
    .A2(_2569_),
    .B(_2469_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6024_ (.A1(_2432_),
    .A2(_2561_),
    .B1(_2567_),
    .B2(_2570_),
    .C(_2514_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6025_ (.I0(\registers[28][12] ),
    .I1(\registers[29][12] ),
    .I2(\registers[30][12] ),
    .I3(\registers[31][12] ),
    .S0(_2476_),
    .S1(_2477_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6026_ (.I0(\registers[24][12] ),
    .I1(\registers[25][12] ),
    .I2(\registers[26][12] ),
    .I3(\registers[27][12] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6027_ (.I0(_2572_),
    .I1(_2573_),
    .S(_2482_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6028_ (.I0(\registers[16][12] ),
    .I1(\registers[17][12] ),
    .S(_2548_),
    .Z(_2575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6029_ (.I0(\registers[18][12] ),
    .I1(\registers[19][12] ),
    .S(_2460_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6030_ (.I0(\registers[20][12] ),
    .I1(\registers[21][12] ),
    .S(_2489_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6031_ (.I0(\registers[22][12] ),
    .I1(\registers[23][12] ),
    .S(_2552_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6032_ (.I0(_2575_),
    .I1(_2576_),
    .I2(_2577_),
    .I3(_2578_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6033_ (.A1(_2517_),
    .A2(_2574_),
    .B1(_2579_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6034_ (.A1(net83),
    .A2(_2499_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6035_ (.A1(_2571_),
    .A2(_2580_),
    .B(_2581_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6036_ (.I(_2436_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6037_ (.I0(\registers[28][13] ),
    .I1(\registers[29][13] ),
    .I2(\registers[30][13] ),
    .I3(\registers[31][13] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6038_ (.I0(\registers[24][13] ),
    .I1(\registers[25][13] ),
    .I2(\registers[26][13] ),
    .I3(\registers[27][13] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6039_ (.I0(_2583_),
    .I1(_2584_),
    .S(_2445_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6040_ (.I0(\registers[18][13] ),
    .I1(\registers[19][13] ),
    .S(_2451_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6041_ (.I(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6042_ (.I0(\registers[16][13] ),
    .I1(\registers[17][13] ),
    .S(_2456_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6043_ (.I0(\registers[22][13] ),
    .I1(\registers[23][13] ),
    .S(_2507_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6044_ (.A1(_2455_),
    .A2(_2588_),
    .B1(_2589_),
    .B2(_2459_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6045_ (.A1(_2449_),
    .A2(_2587_),
    .B(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6046_ (.I0(\registers[20][13] ),
    .I1(\registers[21][13] ),
    .S(_2466_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6047_ (.I(_2592_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6048_ (.A1(_2465_),
    .A2(_2593_),
    .B(_2469_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6049_ (.A1(_2432_),
    .A2(_2585_),
    .B1(_2591_),
    .B2(_2594_),
    .C(_2472_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6050_ (.I0(\registers[12][13] ),
    .I1(\registers[13][13] ),
    .I2(\registers[14][13] ),
    .I3(\registers[15][13] ),
    .S0(_2476_),
    .S1(_2477_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6051_ (.I(_2434_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6052_ (.I0(\registers[8][13] ),
    .I1(\registers[9][13] ),
    .I2(\registers[10][13] ),
    .I3(\registers[11][13] ),
    .S0(_2597_),
    .S1(_2480_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6053_ (.I0(_2596_),
    .I1(_2598_),
    .S(_2482_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6054_ (.I0(\registers[0][13] ),
    .I1(\registers[1][13] ),
    .S(_2548_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6055_ (.I0(\registers[2][13] ),
    .I1(\registers[3][13] ),
    .S(_2460_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6056_ (.I(_2488_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6057_ (.I0(\registers[4][13] ),
    .I1(\registers[5][13] ),
    .S(_2602_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6058_ (.I0(\registers[6][13] ),
    .I1(\registers[7][13] ),
    .S(_2552_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6059_ (.I0(_2600_),
    .I1(_2601_),
    .I2(_2603_),
    .I3(_2604_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6060_ (.A1(_2475_),
    .A2(_2599_),
    .B1(_2605_),
    .B2(_2485_),
    .C(_2495_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6061_ (.A1(net84),
    .A2(_2499_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6062_ (.A1(_2595_),
    .A2(_2606_),
    .B(_2607_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6063_ (.I0(\registers[12][14] ),
    .I1(\registers[13][14] ),
    .I2(\registers[14][14] ),
    .I3(\registers[15][14] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6064_ (.I0(\registers[8][14] ),
    .I1(\registers[9][14] ),
    .I2(\registers[10][14] ),
    .I3(\registers[11][14] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6065_ (.I0(_2608_),
    .I1(_2609_),
    .S(_2445_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6066_ (.I0(\registers[2][14] ),
    .I1(\registers[3][14] ),
    .S(_2451_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6067_ (.I(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6068_ (.I0(\registers[0][14] ),
    .I1(\registers[1][14] ),
    .S(_2456_),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6069_ (.I0(\registers[6][14] ),
    .I1(\registers[7][14] ),
    .S(_2507_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6070_ (.A1(_2455_),
    .A2(_2613_),
    .B1(_2614_),
    .B2(_2459_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6071_ (.A1(_2449_),
    .A2(_2612_),
    .B(_2615_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6072_ (.I0(\registers[4][14] ),
    .I1(\registers[5][14] ),
    .S(_2466_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6073_ (.I(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6074_ (.A1(_2465_),
    .A2(_2618_),
    .B(_2469_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6075_ (.A1(_2432_),
    .A2(_2610_),
    .B1(_2616_),
    .B2(_2619_),
    .C(_2514_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6076_ (.I0(\registers[28][14] ),
    .I1(\registers[29][14] ),
    .I2(\registers[30][14] ),
    .I3(\registers[31][14] ),
    .S0(_2476_),
    .S1(_2477_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6077_ (.I0(\registers[24][14] ),
    .I1(\registers[25][14] ),
    .I2(\registers[26][14] ),
    .I3(\registers[27][14] ),
    .S0(_2597_),
    .S1(_2480_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6078_ (.I0(_2621_),
    .I1(_2622_),
    .S(_2482_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6079_ (.I0(\registers[16][14] ),
    .I1(\registers[17][14] ),
    .S(_2548_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6080_ (.I0(\registers[18][14] ),
    .I1(\registers[19][14] ),
    .S(_2460_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6081_ (.I0(\registers[20][14] ),
    .I1(\registers[21][14] ),
    .S(_2602_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6082_ (.I0(\registers[22][14] ),
    .I1(\registers[23][14] ),
    .S(_2552_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6083_ (.I0(_2624_),
    .I1(_2625_),
    .I2(_2626_),
    .I3(_2627_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6084_ (.A1(_2517_),
    .A2(_2623_),
    .B1(_2628_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6085_ (.A1(net85),
    .A2(_2499_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6086_ (.A1(_2620_),
    .A2(_2629_),
    .B(_2630_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6087_ (.I0(\registers[12][15] ),
    .I1(\registers[13][15] ),
    .I2(\registers[14][15] ),
    .I3(\registers[15][15] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6088_ (.I0(\registers[8][15] ),
    .I1(\registers[9][15] ),
    .I2(\registers[10][15] ),
    .I3(\registers[11][15] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6089_ (.I0(_2631_),
    .I1(_2632_),
    .S(_2445_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6090_ (.I0(\registers[2][15] ),
    .I1(\registers[3][15] ),
    .S(_2451_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6091_ (.I(_2634_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6092_ (.I0(\registers[0][15] ),
    .I1(\registers[1][15] ),
    .S(_2456_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6093_ (.I0(\registers[6][15] ),
    .I1(\registers[7][15] ),
    .S(_2507_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6094_ (.A1(_2455_),
    .A2(_2636_),
    .B1(_2637_),
    .B2(_2459_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6095_ (.A1(_2449_),
    .A2(_2635_),
    .B(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6096_ (.I0(\registers[4][15] ),
    .I1(\registers[5][15] ),
    .S(_2466_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6097_ (.I(_2640_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6098_ (.A1(_2465_),
    .A2(_2641_),
    .B(_2469_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6099_ (.A1(_2432_),
    .A2(_2633_),
    .B1(_2639_),
    .B2(_2642_),
    .C(_2514_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6100_ (.I(_2434_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6101_ (.I0(\registers[28][15] ),
    .I1(\registers[29][15] ),
    .I2(\registers[30][15] ),
    .I3(\registers[31][15] ),
    .S0(_2644_),
    .S1(_2477_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6102_ (.I(_2447_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6103_ (.I0(\registers[24][15] ),
    .I1(\registers[25][15] ),
    .I2(\registers[26][15] ),
    .I3(\registers[27][15] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6104_ (.I0(_2645_),
    .I1(_2647_),
    .S(_2482_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6105_ (.I(_2488_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6106_ (.I0(\registers[16][15] ),
    .I1(\registers[17][15] ),
    .S(_2649_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6107_ (.I(_2488_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6108_ (.I0(\registers[18][15] ),
    .I1(\registers[19][15] ),
    .S(_2651_),
    .Z(_2652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6109_ (.I0(\registers[20][15] ),
    .I1(\registers[21][15] ),
    .S(_2602_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6110_ (.I(_2488_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6111_ (.I0(\registers[22][15] ),
    .I1(\registers[23][15] ),
    .S(_2654_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6112_ (.I0(_2650_),
    .I1(_2652_),
    .I2(_2653_),
    .I3(_2655_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6113_ (.A1(_2517_),
    .A2(_2648_),
    .B1(_2656_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6114_ (.A1(net86),
    .A2(_2499_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6115_ (.A1(_2643_),
    .A2(_2657_),
    .B(_2658_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6116_ (.I0(\registers[12][16] ),
    .I1(\registers[13][16] ),
    .I2(\registers[14][16] ),
    .I3(\registers[15][16] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6117_ (.I0(\registers[8][16] ),
    .I1(\registers[9][16] ),
    .I2(\registers[10][16] ),
    .I3(\registers[11][16] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6118_ (.I0(_2659_),
    .I1(_2660_),
    .S(_2445_),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6119_ (.I0(\registers[2][16] ),
    .I1(\registers[3][16] ),
    .S(_2451_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6120_ (.I(_2662_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6121_ (.I0(\registers[0][16] ),
    .I1(\registers[1][16] ),
    .S(_2456_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6122_ (.I(_2439_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6123_ (.I0(\registers[6][16] ),
    .I1(\registers[7][16] ),
    .S(_2665_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6124_ (.A1(_2455_),
    .A2(_2664_),
    .B1(_2666_),
    .B2(_2459_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6125_ (.A1(_2449_),
    .A2(_2663_),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6126_ (.I0(\registers[4][16] ),
    .I1(\registers[5][16] ),
    .S(_2466_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6127_ (.I(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6128_ (.A1(_2465_),
    .A2(_2670_),
    .B(_2469_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6129_ (.A1(_2432_),
    .A2(_2661_),
    .B1(_2668_),
    .B2(_2671_),
    .C(_2514_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6130_ (.I0(\registers[28][16] ),
    .I1(\registers[29][16] ),
    .I2(\registers[30][16] ),
    .I3(\registers[31][16] ),
    .S0(_2644_),
    .S1(_2477_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6131_ (.I0(\registers[24][16] ),
    .I1(\registers[25][16] ),
    .I2(\registers[26][16] ),
    .I3(\registers[27][16] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6132_ (.I0(_2673_),
    .I1(_2674_),
    .S(_2482_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6133_ (.I0(\registers[16][16] ),
    .I1(\registers[17][16] ),
    .S(_2649_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6134_ (.I0(\registers[18][16] ),
    .I1(\registers[19][16] ),
    .S(_2651_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6135_ (.I0(\registers[20][16] ),
    .I1(\registers[21][16] ),
    .S(_2602_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6136_ (.I0(\registers[22][16] ),
    .I1(\registers[23][16] ),
    .S(_2654_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6137_ (.I0(_2676_),
    .I1(_2677_),
    .I2(_2678_),
    .I3(_2679_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6138_ (.A1(_2517_),
    .A2(_2675_),
    .B1(_2680_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6139_ (.A1(net87),
    .A2(_2499_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6140_ (.A1(_2672_),
    .A2(_2681_),
    .B(_2682_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6141_ (.I0(\registers[12][17] ),
    .I1(\registers[13][17] ),
    .I2(\registers[14][17] ),
    .I3(\registers[15][17] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6142_ (.I0(\registers[8][17] ),
    .I1(\registers[9][17] ),
    .I2(\registers[10][17] ),
    .I3(\registers[11][17] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6143_ (.I(_2444_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6144_ (.I0(_2683_),
    .I1(_2684_),
    .S(_2685_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6145_ (.I0(\registers[2][17] ),
    .I1(\registers[3][17] ),
    .S(_2451_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6146_ (.I(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6147_ (.I(_2439_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6148_ (.I0(\registers[0][17] ),
    .I1(\registers[1][17] ),
    .S(_2689_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6149_ (.I0(\registers[6][17] ),
    .I1(\registers[7][17] ),
    .S(_2665_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6150_ (.A1(_2455_),
    .A2(_2690_),
    .B1(_2691_),
    .B2(_2459_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6151_ (.A1(_2449_),
    .A2(_2688_),
    .B(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6152_ (.I(_2450_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6153_ (.I0(\registers[4][17] ),
    .I1(\registers[5][17] ),
    .S(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6154_ (.I(_2695_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6155_ (.I(_2431_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6156_ (.A1(_2465_),
    .A2(_2696_),
    .B(_2697_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6157_ (.A1(_2432_),
    .A2(_2686_),
    .B1(_2693_),
    .B2(_2698_),
    .C(_2514_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6158_ (.I(_2447_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6159_ (.I0(\registers[28][17] ),
    .I1(\registers[29][17] ),
    .I2(\registers[30][17] ),
    .I3(\registers[31][17] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6160_ (.I0(\registers[24][17] ),
    .I1(\registers[25][17] ),
    .I2(\registers[26][17] ),
    .I3(\registers[27][17] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6161_ (.I0(_2701_),
    .I1(_2702_),
    .S(_2482_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6162_ (.I0(\registers[16][17] ),
    .I1(\registers[17][17] ),
    .S(_2649_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6163_ (.I0(\registers[18][17] ),
    .I1(\registers[19][17] ),
    .S(_2651_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6164_ (.I0(\registers[20][17] ),
    .I1(\registers[21][17] ),
    .S(_2602_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6165_ (.I0(\registers[22][17] ),
    .I1(\registers[23][17] ),
    .S(_2654_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6166_ (.I0(_2704_),
    .I1(_2705_),
    .I2(_2706_),
    .I3(_2707_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6167_ (.A1(_2517_),
    .A2(_2703_),
    .B1(_2708_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6168_ (.A1(net88),
    .A2(_2499_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6169_ (.A1(_2699_),
    .A2(_2709_),
    .B(_2710_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6170_ (.I0(\registers[12][18] ),
    .I1(\registers[13][18] ),
    .I2(\registers[14][18] ),
    .I3(\registers[15][18] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6171_ (.I0(\registers[8][18] ),
    .I1(\registers[9][18] ),
    .I2(\registers[10][18] ),
    .I3(\registers[11][18] ),
    .S0(_2440_),
    .S1(_2532_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6172_ (.I0(_2711_),
    .I1(_2712_),
    .S(_2685_),
    .Z(_2713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6173_ (.I0(\registers[2][18] ),
    .I1(\registers[3][18] ),
    .S(_2451_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6174_ (.I(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6175_ (.I0(\registers[0][18] ),
    .I1(\registers[1][18] ),
    .S(_2689_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6176_ (.I0(\registers[6][18] ),
    .I1(\registers[7][18] ),
    .S(_2665_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6177_ (.A1(_2455_),
    .A2(_2716_),
    .B1(_2717_),
    .B2(_2459_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6178_ (.A1(_2449_),
    .A2(_2715_),
    .B(_2718_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6179_ (.I0(\registers[4][18] ),
    .I1(\registers[5][18] ),
    .S(_2694_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6180_ (.I(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6181_ (.A1(_2465_),
    .A2(_2721_),
    .B(_2697_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6182_ (.A1(_2432_),
    .A2(_2713_),
    .B1(_2719_),
    .B2(_2722_),
    .C(_2514_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6183_ (.I0(\registers[28][18] ),
    .I1(\registers[29][18] ),
    .I2(\registers[30][18] ),
    .I3(\registers[31][18] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6184_ (.I0(\registers[24][18] ),
    .I1(\registers[25][18] ),
    .I2(\registers[26][18] ),
    .I3(\registers[27][18] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6185_ (.I0(_2724_),
    .I1(_2725_),
    .S(_2482_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6186_ (.I0(\registers[16][18] ),
    .I1(\registers[17][18] ),
    .S(_2649_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6187_ (.I0(\registers[18][18] ),
    .I1(\registers[19][18] ),
    .S(_2651_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6188_ (.I0(\registers[20][18] ),
    .I1(\registers[21][18] ),
    .S(_2602_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6189_ (.I0(\registers[22][18] ),
    .I1(\registers[23][18] ),
    .S(_2654_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6190_ (.I0(_2727_),
    .I1(_2728_),
    .I2(_2729_),
    .I3(_2730_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6191_ (.A1(_2517_),
    .A2(_2726_),
    .B1(_2731_),
    .B2(_2522_),
    .C(_2495_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6192_ (.A1(net89),
    .A2(_2499_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6193_ (.A1(_2723_),
    .A2(_2732_),
    .B(_2733_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6194_ (.I(_2431_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6195_ (.I0(\registers[12][19] ),
    .I1(\registers[13][19] ),
    .I2(\registers[14][19] ),
    .I3(\registers[15][19] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6196_ (.I(_2439_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6197_ (.I0(\registers[8][19] ),
    .I1(\registers[9][19] ),
    .I2(\registers[10][19] ),
    .I3(\registers[11][19] ),
    .S0(_2736_),
    .S1(_2532_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6198_ (.I0(_2735_),
    .I1(_2737_),
    .S(_2685_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6199_ (.I(_2448_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6200_ (.I(_2450_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6201_ (.I0(\registers[2][19] ),
    .I1(\registers[3][19] ),
    .S(_2740_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6202_ (.I(_2741_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6203_ (.I(_2454_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6204_ (.I0(\registers[0][19] ),
    .I1(\registers[1][19] ),
    .S(_2689_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6205_ (.I0(\registers[6][19] ),
    .I1(\registers[7][19] ),
    .S(_2665_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6206_ (.I(_2458_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6207_ (.A1(_2743_),
    .A2(_2744_),
    .B1(_2745_),
    .B2(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6208_ (.A1(_2739_),
    .A2(_2742_),
    .B(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6209_ (.I(_2464_),
    .Z(_2749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6210_ (.I0(\registers[4][19] ),
    .I1(\registers[5][19] ),
    .S(_2694_),
    .Z(_2750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6211_ (.I(_2750_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6212_ (.A1(_2749_),
    .A2(_2751_),
    .B(_2697_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6213_ (.A1(_2734_),
    .A2(_2738_),
    .B1(_2748_),
    .B2(_2752_),
    .C(_2514_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6214_ (.I0(\registers[28][19] ),
    .I1(\registers[29][19] ),
    .I2(\registers[30][19] ),
    .I3(\registers[31][19] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6215_ (.I0(\registers[24][19] ),
    .I1(\registers[25][19] ),
    .I2(\registers[26][19] ),
    .I3(\registers[27][19] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6216_ (.I(_2444_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6217_ (.I0(_2754_),
    .I1(_2755_),
    .S(_2756_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6218_ (.I0(\registers[16][19] ),
    .I1(\registers[17][19] ),
    .S(_2649_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6219_ (.I0(\registers[18][19] ),
    .I1(\registers[19][19] ),
    .S(_2651_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6220_ (.I0(\registers[20][19] ),
    .I1(\registers[21][19] ),
    .S(_2602_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6221_ (.I0(\registers[22][19] ),
    .I1(\registers[23][19] ),
    .S(_2654_),
    .Z(_2761_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6222_ (.I0(_2758_),
    .I1(_2759_),
    .I2(_2760_),
    .I3(_2761_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6223_ (.I(_2494_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6224_ (.A1(_2517_),
    .A2(_2757_),
    .B1(_2762_),
    .B2(_2522_),
    .C(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6225_ (.I(_2498_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6226_ (.A1(net90),
    .A2(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6227_ (.A1(_2753_),
    .A2(_2764_),
    .B(_2766_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6228_ (.I0(\registers[28][1] ),
    .I1(\registers[29][1] ),
    .I2(\registers[30][1] ),
    .I3(\registers[31][1] ),
    .S0(_2530_),
    .S1(_2582_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6229_ (.I0(\registers[24][1] ),
    .I1(\registers[25][1] ),
    .I2(\registers[26][1] ),
    .I3(\registers[27][1] ),
    .S0(_2736_),
    .S1(_2532_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6230_ (.I0(_2767_),
    .I1(_2768_),
    .S(_2685_),
    .Z(_2769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6231_ (.I0(\registers[18][1] ),
    .I1(\registers[19][1] ),
    .S(_2740_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6232_ (.I(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6233_ (.I0(\registers[16][1] ),
    .I1(\registers[17][1] ),
    .S(_2689_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6234_ (.I0(\registers[22][1] ),
    .I1(\registers[23][1] ),
    .S(_2665_),
    .Z(_2773_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6235_ (.A1(_2743_),
    .A2(_2772_),
    .B1(_2773_),
    .B2(_2746_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6236_ (.A1(_2739_),
    .A2(_2771_),
    .B(_2774_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6237_ (.I0(\registers[20][1] ),
    .I1(\registers[21][1] ),
    .S(_2694_),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6238_ (.I(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6239_ (.A1(_2749_),
    .A2(_2777_),
    .B(_2697_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6240_ (.A1(_2734_),
    .A2(_2769_),
    .B1(_2775_),
    .B2(_2778_),
    .C(_2472_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6241_ (.I0(\registers[12][1] ),
    .I1(\registers[13][1] ),
    .I2(\registers[14][1] ),
    .I3(\registers[15][1] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6242_ (.I0(\registers[8][1] ),
    .I1(\registers[9][1] ),
    .I2(\registers[10][1] ),
    .I3(\registers[11][1] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6243_ (.I0(_2780_),
    .I1(_2781_),
    .S(_2756_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6244_ (.I0(\registers[0][1] ),
    .I1(\registers[1][1] ),
    .S(_2649_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6245_ (.I0(\registers[2][1] ),
    .I1(\registers[3][1] ),
    .S(_2651_),
    .Z(_2784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6246_ (.I0(\registers[4][1] ),
    .I1(\registers[5][1] ),
    .S(_2602_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6247_ (.I0(\registers[6][1] ),
    .I1(\registers[7][1] ),
    .S(_2654_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6248_ (.I0(_2783_),
    .I1(_2784_),
    .I2(_2785_),
    .I3(_2786_),
    .S0(_2554_),
    .S1(_2555_),
    .Z(_2787_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6249_ (.A1(_2475_),
    .A2(_2782_),
    .B1(_2787_),
    .B2(_2485_),
    .C(_2763_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6250_ (.A1(net91),
    .A2(_2765_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6251_ (.A1(_2779_),
    .A2(_2788_),
    .B(_2789_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6252_ (.I(_2434_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6253_ (.I0(\registers[12][20] ),
    .I1(\registers[13][20] ),
    .I2(\registers[14][20] ),
    .I3(\registers[15][20] ),
    .S0(_2790_),
    .S1(_2582_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6254_ (.I(_2436_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6255_ (.I0(\registers[8][20] ),
    .I1(\registers[9][20] ),
    .I2(\registers[10][20] ),
    .I3(\registers[11][20] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6256_ (.I0(_2791_),
    .I1(_2793_),
    .S(_2685_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6257_ (.I0(\registers[2][20] ),
    .I1(\registers[3][20] ),
    .S(_2740_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6258_ (.I(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6259_ (.I0(\registers[0][20] ),
    .I1(\registers[1][20] ),
    .S(_2689_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6260_ (.I0(\registers[6][20] ),
    .I1(\registers[7][20] ),
    .S(_2665_),
    .Z(_2798_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6261_ (.A1(_2743_),
    .A2(_2797_),
    .B1(_2798_),
    .B2(_2746_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6262_ (.A1(_2739_),
    .A2(_2796_),
    .B(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6263_ (.I0(\registers[4][20] ),
    .I1(\registers[5][20] ),
    .S(_2694_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6264_ (.I(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6265_ (.A1(_2749_),
    .A2(_2802_),
    .B(_2697_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6266_ (.A1(_2734_),
    .A2(_2794_),
    .B1(_2800_),
    .B2(_2803_),
    .C(_2514_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6267_ (.I0(\registers[28][20] ),
    .I1(\registers[29][20] ),
    .I2(\registers[30][20] ),
    .I3(\registers[31][20] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2805_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6268_ (.I0(\registers[24][20] ),
    .I1(\registers[25][20] ),
    .I2(\registers[26][20] ),
    .I3(\registers[27][20] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6269_ (.I0(_2805_),
    .I1(_2806_),
    .S(_2756_),
    .Z(_2807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6270_ (.I0(\registers[16][20] ),
    .I1(\registers[17][20] ),
    .S(_2649_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6271_ (.I0(\registers[18][20] ),
    .I1(\registers[19][20] ),
    .S(_2651_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6272_ (.I0(\registers[20][20] ),
    .I1(\registers[21][20] ),
    .S(_2602_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6273_ (.I0(\registers[22][20] ),
    .I1(\registers[23][20] ),
    .S(_2654_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6274_ (.I(_2447_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6275_ (.I(net4),
    .Z(_2813_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6276_ (.I0(_2808_),
    .I1(_2809_),
    .I2(_2810_),
    .I3(_2811_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6277_ (.A1(_2517_),
    .A2(_2807_),
    .B1(_2814_),
    .B2(_2522_),
    .C(_2763_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6278_ (.A1(net92),
    .A2(_2765_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6279_ (.A1(_2804_),
    .A2(_2815_),
    .B(_2816_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6280_ (.I0(\registers[12][21] ),
    .I1(\registers[13][21] ),
    .I2(\registers[14][21] ),
    .I3(\registers[15][21] ),
    .S0(_2790_),
    .S1(_2582_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6281_ (.I0(\registers[8][21] ),
    .I1(\registers[9][21] ),
    .I2(\registers[10][21] ),
    .I3(\registers[11][21] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6282_ (.I0(_2817_),
    .I1(_2818_),
    .S(_2685_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6283_ (.I0(\registers[2][21] ),
    .I1(\registers[3][21] ),
    .S(_2740_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6284_ (.I(_2820_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6285_ (.I0(\registers[0][21] ),
    .I1(\registers[1][21] ),
    .S(_2689_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6286_ (.I0(\registers[6][21] ),
    .I1(\registers[7][21] ),
    .S(_2665_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6287_ (.A1(_2743_),
    .A2(_2822_),
    .B1(_2823_),
    .B2(_2746_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6288_ (.A1(_2739_),
    .A2(_2821_),
    .B(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6289_ (.I0(\registers[4][21] ),
    .I1(\registers[5][21] ),
    .S(_2694_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6290_ (.I(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6291_ (.A1(_2749_),
    .A2(_2827_),
    .B(_2697_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6292_ (.I(net6),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6293_ (.A1(_2734_),
    .A2(_2819_),
    .B1(_2825_),
    .B2(_2828_),
    .C(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6294_ (.I(_2516_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6295_ (.I0(\registers[28][21] ),
    .I1(\registers[29][21] ),
    .I2(\registers[30][21] ),
    .I3(\registers[31][21] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6296_ (.I0(\registers[24][21] ),
    .I1(\registers[25][21] ),
    .I2(\registers[26][21] ),
    .I3(\registers[27][21] ),
    .S0(_2597_),
    .S1(_2646_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6297_ (.I0(_2832_),
    .I1(_2833_),
    .S(_2756_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6298_ (.I0(\registers[16][21] ),
    .I1(\registers[17][21] ),
    .S(_2649_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6299_ (.I0(\registers[18][21] ),
    .I1(\registers[19][21] ),
    .S(_2651_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6300_ (.I0(\registers[20][21] ),
    .I1(\registers[21][21] ),
    .S(_2602_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6301_ (.I0(\registers[22][21] ),
    .I1(\registers[23][21] ),
    .S(_2654_),
    .Z(_2838_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6302_ (.I0(_2835_),
    .I1(_2836_),
    .I2(_2837_),
    .I3(_2838_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6303_ (.I(_2521_),
    .Z(_2840_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6304_ (.A1(_2831_),
    .A2(_2834_),
    .B1(_2839_),
    .B2(_2840_),
    .C(_2763_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6305_ (.A1(net93),
    .A2(_2765_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6306_ (.A1(_2830_),
    .A2(_2841_),
    .B(_2842_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6307_ (.I(_2436_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6308_ (.I0(\registers[28][22] ),
    .I1(\registers[29][22] ),
    .I2(\registers[30][22] ),
    .I3(\registers[31][22] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6309_ (.I0(\registers[24][22] ),
    .I1(\registers[25][22] ),
    .I2(\registers[26][22] ),
    .I3(\registers[27][22] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6310_ (.I0(_2844_),
    .I1(_2845_),
    .S(_2685_),
    .Z(_2846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6311_ (.I0(\registers[18][22] ),
    .I1(\registers[19][22] ),
    .S(_2740_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6312_ (.I(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6313_ (.I0(\registers[16][22] ),
    .I1(\registers[17][22] ),
    .S(_2689_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6314_ (.I0(\registers[22][22] ),
    .I1(\registers[23][22] ),
    .S(_2665_),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6315_ (.A1(_2743_),
    .A2(_2849_),
    .B1(_2850_),
    .B2(_2746_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6316_ (.A1(_2739_),
    .A2(_2848_),
    .B(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6317_ (.I0(\registers[20][22] ),
    .I1(\registers[21][22] ),
    .S(_2694_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6318_ (.I(_2853_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6319_ (.A1(_2749_),
    .A2(_2854_),
    .B(_2697_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6320_ (.A1(_2734_),
    .A2(_2846_),
    .B1(_2852_),
    .B2(_2855_),
    .C(_2472_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6321_ (.I0(\registers[12][22] ),
    .I1(\registers[13][22] ),
    .I2(\registers[14][22] ),
    .I3(\registers[15][22] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6322_ (.I(_2434_),
    .Z(_2858_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6323_ (.I0(\registers[8][22] ),
    .I1(\registers[9][22] ),
    .I2(\registers[10][22] ),
    .I3(\registers[11][22] ),
    .S0(_2858_),
    .S1(_2646_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6324_ (.I0(_2857_),
    .I1(_2859_),
    .S(_2756_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6325_ (.I0(\registers[0][22] ),
    .I1(\registers[1][22] ),
    .S(_2649_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6326_ (.I0(\registers[2][22] ),
    .I1(\registers[3][22] ),
    .S(_2651_),
    .Z(_2862_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6327_ (.I(_2433_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6328_ (.I0(\registers[4][22] ),
    .I1(\registers[5][22] ),
    .S(_2863_),
    .Z(_2864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6329_ (.I0(\registers[6][22] ),
    .I1(\registers[7][22] ),
    .S(_2654_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6330_ (.I0(_2861_),
    .I1(_2862_),
    .I2(_2864_),
    .I3(_2865_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6331_ (.A1(_2475_),
    .A2(_2860_),
    .B1(_2866_),
    .B2(_2485_),
    .C(_2763_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6332_ (.A1(net94),
    .A2(_2765_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6333_ (.A1(_2856_),
    .A2(_2867_),
    .B(_2868_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6334_ (.I0(\registers[28][23] ),
    .I1(\registers[29][23] ),
    .I2(\registers[30][23] ),
    .I3(\registers[31][23] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6335_ (.I0(\registers[24][23] ),
    .I1(\registers[25][23] ),
    .I2(\registers[26][23] ),
    .I3(\registers[27][23] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6336_ (.I0(_2869_),
    .I1(_2870_),
    .S(_2685_),
    .Z(_2871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6337_ (.I0(\registers[18][23] ),
    .I1(\registers[19][23] ),
    .S(_2740_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6338_ (.I(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6339_ (.I0(\registers[16][23] ),
    .I1(\registers[17][23] ),
    .S(_2689_),
    .Z(_2874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6340_ (.I0(\registers[22][23] ),
    .I1(\registers[23][23] ),
    .S(_2665_),
    .Z(_2875_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6341_ (.A1(_2743_),
    .A2(_2874_),
    .B1(_2875_),
    .B2(_2746_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6342_ (.A1(_2739_),
    .A2(_2873_),
    .B(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6343_ (.I0(\registers[20][23] ),
    .I1(\registers[21][23] ),
    .S(_2694_),
    .Z(_2878_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6344_ (.I(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6345_ (.A1(_2749_),
    .A2(_2879_),
    .B(_2697_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6346_ (.A1(_2734_),
    .A2(_2871_),
    .B1(_2877_),
    .B2(_2880_),
    .C(_2472_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6347_ (.I0(\registers[12][23] ),
    .I1(\registers[13][23] ),
    .I2(\registers[14][23] ),
    .I3(\registers[15][23] ),
    .S0(_2644_),
    .S1(_2700_),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6348_ (.I0(\registers[8][23] ),
    .I1(\registers[9][23] ),
    .I2(\registers[10][23] ),
    .I3(\registers[11][23] ),
    .S0(_2858_),
    .S1(_2646_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6349_ (.I0(_2882_),
    .I1(_2883_),
    .S(_2756_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6350_ (.I0(\registers[0][23] ),
    .I1(\registers[1][23] ),
    .S(_2649_),
    .Z(_2885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6351_ (.I0(\registers[2][23] ),
    .I1(\registers[3][23] ),
    .S(_2651_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6352_ (.I0(\registers[4][23] ),
    .I1(\registers[5][23] ),
    .S(_2863_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6353_ (.I0(\registers[6][23] ),
    .I1(\registers[7][23] ),
    .S(_2654_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6354_ (.I0(_2885_),
    .I1(_2886_),
    .I2(_2887_),
    .I3(_2888_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6355_ (.A1(_2475_),
    .A2(_2884_),
    .B1(_2889_),
    .B2(_2485_),
    .C(_2763_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6356_ (.A1(net95),
    .A2(_2765_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6357_ (.A1(_2881_),
    .A2(_2890_),
    .B(_2891_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6358_ (.I0(\registers[28][24] ),
    .I1(\registers[29][24] ),
    .I2(\registers[30][24] ),
    .I3(\registers[31][24] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6359_ (.I0(\registers[24][24] ),
    .I1(\registers[25][24] ),
    .I2(\registers[26][24] ),
    .I3(\registers[27][24] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6360_ (.I0(_2892_),
    .I1(_2893_),
    .S(_2685_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6361_ (.I0(\registers[18][24] ),
    .I1(\registers[19][24] ),
    .S(_2740_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6362_ (.I(_2895_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6363_ (.I0(\registers[16][24] ),
    .I1(\registers[17][24] ),
    .S(_2689_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6364_ (.I0(\registers[22][24] ),
    .I1(\registers[23][24] ),
    .S(_2665_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6365_ (.A1(_2743_),
    .A2(_2897_),
    .B1(_2898_),
    .B2(_2746_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6366_ (.A1(_2739_),
    .A2(_2896_),
    .B(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6367_ (.I0(\registers[20][24] ),
    .I1(\registers[21][24] ),
    .S(_2694_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6368_ (.I(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6369_ (.A1(_2749_),
    .A2(_2902_),
    .B(_2697_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6370_ (.A1(_2734_),
    .A2(_2894_),
    .B1(_2900_),
    .B2(_2903_),
    .C(_2472_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6371_ (.I(_2434_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6372_ (.I0(\registers[12][24] ),
    .I1(\registers[13][24] ),
    .I2(\registers[14][24] ),
    .I3(\registers[15][24] ),
    .S0(_2905_),
    .S1(_2700_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6373_ (.I(_2436_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6374_ (.I0(\registers[8][24] ),
    .I1(\registers[9][24] ),
    .I2(\registers[10][24] ),
    .I3(\registers[11][24] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6375_ (.I0(_2906_),
    .I1(_2908_),
    .S(_2756_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6376_ (.I(_2488_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6377_ (.I0(\registers[0][24] ),
    .I1(\registers[1][24] ),
    .S(_2910_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6378_ (.I(_2488_),
    .Z(_2912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6379_ (.I0(\registers[2][24] ),
    .I1(\registers[3][24] ),
    .S(_2912_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6380_ (.I0(\registers[4][24] ),
    .I1(\registers[5][24] ),
    .S(_2863_),
    .Z(_2914_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6381_ (.I(_2488_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6382_ (.I0(\registers[6][24] ),
    .I1(\registers[7][24] ),
    .S(_2915_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6383_ (.I0(_2911_),
    .I1(_2913_),
    .I2(_2914_),
    .I3(_2916_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2917_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6384_ (.A1(_2475_),
    .A2(_2909_),
    .B1(_2917_),
    .B2(_2485_),
    .C(_2763_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6385_ (.A1(net96),
    .A2(_2765_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6386_ (.A1(_2904_),
    .A2(_2918_),
    .B(_2919_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6387_ (.I0(\registers[12][25] ),
    .I1(\registers[13][25] ),
    .I2(\registers[14][25] ),
    .I3(\registers[15][25] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6388_ (.I0(\registers[8][25] ),
    .I1(\registers[9][25] ),
    .I2(\registers[10][25] ),
    .I3(\registers[11][25] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6389_ (.I0(_2920_),
    .I1(_2921_),
    .S(_2685_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6390_ (.I0(\registers[2][25] ),
    .I1(\registers[3][25] ),
    .S(_2740_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6391_ (.I(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6392_ (.I0(\registers[0][25] ),
    .I1(\registers[1][25] ),
    .S(_2689_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6393_ (.I(_2439_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6394_ (.I0(\registers[6][25] ),
    .I1(\registers[7][25] ),
    .S(_2926_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6395_ (.A1(_2743_),
    .A2(_2925_),
    .B1(_2927_),
    .B2(_2746_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6396_ (.A1(_2739_),
    .A2(_2924_),
    .B(_2928_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6397_ (.I0(\registers[4][25] ),
    .I1(\registers[5][25] ),
    .S(_2694_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6398_ (.I(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6399_ (.A1(_2749_),
    .A2(_2931_),
    .B(_2697_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6400_ (.A1(_2734_),
    .A2(_2922_),
    .B1(_2929_),
    .B2(_2932_),
    .C(_2829_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6401_ (.I0(\registers[28][25] ),
    .I1(\registers[29][25] ),
    .I2(\registers[30][25] ),
    .I3(\registers[31][25] ),
    .S0(_2905_),
    .S1(_2700_),
    .Z(_2934_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6402_ (.I0(\registers[24][25] ),
    .I1(\registers[25][25] ),
    .I2(\registers[26][25] ),
    .I3(\registers[27][25] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6403_ (.I0(_2934_),
    .I1(_2935_),
    .S(_2756_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6404_ (.I0(\registers[16][25] ),
    .I1(\registers[17][25] ),
    .S(_2910_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6405_ (.I0(\registers[18][25] ),
    .I1(\registers[19][25] ),
    .S(_2912_),
    .Z(_2938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6406_ (.I0(\registers[20][25] ),
    .I1(\registers[21][25] ),
    .S(_2863_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6407_ (.I0(\registers[22][25] ),
    .I1(\registers[23][25] ),
    .S(_2915_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6408_ (.I0(_2937_),
    .I1(_2938_),
    .I2(_2939_),
    .I3(_2940_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6409_ (.A1(_2831_),
    .A2(_2936_),
    .B1(_2941_),
    .B2(_2840_),
    .C(_2763_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6410_ (.A1(net97),
    .A2(_2765_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6411_ (.A1(_2933_),
    .A2(_2942_),
    .B(_2943_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6412_ (.I0(\registers[28][26] ),
    .I1(\registers[29][26] ),
    .I2(\registers[30][26] ),
    .I3(\registers[31][26] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2944_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6413_ (.I0(\registers[24][26] ),
    .I1(\registers[25][26] ),
    .I2(\registers[26][26] ),
    .I3(\registers[27][26] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2945_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6414_ (.I(_2444_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6415_ (.I0(_2944_),
    .I1(_2945_),
    .S(_2946_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6416_ (.I0(\registers[18][26] ),
    .I1(\registers[19][26] ),
    .S(_2740_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6417_ (.I(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6418_ (.I(_2439_),
    .Z(_2950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6419_ (.I0(\registers[16][26] ),
    .I1(\registers[17][26] ),
    .S(_2950_),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6420_ (.I0(\registers[22][26] ),
    .I1(\registers[23][26] ),
    .S(_2926_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6421_ (.A1(_2743_),
    .A2(_2951_),
    .B1(_2952_),
    .B2(_2746_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6422_ (.A1(_2739_),
    .A2(_2949_),
    .B(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6423_ (.I(_2450_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6424_ (.I0(\registers[20][26] ),
    .I1(\registers[21][26] ),
    .S(_2955_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6425_ (.I(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6426_ (.I(net5),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6427_ (.A1(_2749_),
    .A2(_2957_),
    .B(_2958_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6428_ (.A1(_2734_),
    .A2(_2947_),
    .B1(_2954_),
    .B2(_2959_),
    .C(_2472_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6429_ (.I(_2447_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6430_ (.I0(\registers[12][26] ),
    .I1(\registers[13][26] ),
    .I2(\registers[14][26] ),
    .I3(\registers[15][26] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6431_ (.I0(\registers[8][26] ),
    .I1(\registers[9][26] ),
    .I2(\registers[10][26] ),
    .I3(\registers[11][26] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_2963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6432_ (.I0(_2962_),
    .I1(_2963_),
    .S(_2756_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6433_ (.I0(\registers[0][26] ),
    .I1(\registers[1][26] ),
    .S(_2910_),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6434_ (.I0(\registers[2][26] ),
    .I1(\registers[3][26] ),
    .S(_2912_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6435_ (.I0(\registers[4][26] ),
    .I1(\registers[5][26] ),
    .S(_2863_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6436_ (.I0(\registers[6][26] ),
    .I1(\registers[7][26] ),
    .S(_2915_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6437_ (.I0(_2965_),
    .I1(_2966_),
    .I2(_2967_),
    .I3(_2968_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6438_ (.A1(_2475_),
    .A2(_2964_),
    .B1(_2969_),
    .B2(_2485_),
    .C(_2763_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6439_ (.A1(net98),
    .A2(_2765_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6440_ (.A1(_2960_),
    .A2(_2970_),
    .B(_2971_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6441_ (.I0(\registers[12][27] ),
    .I1(\registers[13][27] ),
    .I2(\registers[14][27] ),
    .I3(\registers[15][27] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6442_ (.I0(\registers[8][27] ),
    .I1(\registers[9][27] ),
    .I2(\registers[10][27] ),
    .I3(\registers[11][27] ),
    .S0(_2736_),
    .S1(_2792_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6443_ (.I0(_2972_),
    .I1(_2973_),
    .S(_2946_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6444_ (.I0(\registers[2][27] ),
    .I1(\registers[3][27] ),
    .S(_2740_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6445_ (.I(_2975_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6446_ (.I0(\registers[0][27] ),
    .I1(\registers[1][27] ),
    .S(_2950_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6447_ (.I0(\registers[6][27] ),
    .I1(\registers[7][27] ),
    .S(_2926_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6448_ (.A1(_2743_),
    .A2(_2977_),
    .B1(_2978_),
    .B2(_2746_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6449_ (.A1(_2739_),
    .A2(_2976_),
    .B(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6450_ (.I0(\registers[4][27] ),
    .I1(\registers[5][27] ),
    .S(_2955_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6451_ (.I(_2981_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6452_ (.A1(_2749_),
    .A2(_2982_),
    .B(_2958_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6453_ (.A1(_2734_),
    .A2(_2974_),
    .B1(_2980_),
    .B2(_2983_),
    .C(_2829_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6454_ (.I0(\registers[28][27] ),
    .I1(\registers[29][27] ),
    .I2(\registers[30][27] ),
    .I3(\registers[31][27] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_2985_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6455_ (.I0(\registers[24][27] ),
    .I1(\registers[25][27] ),
    .I2(\registers[26][27] ),
    .I3(\registers[27][27] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6456_ (.I0(_2985_),
    .I1(_2986_),
    .S(_2756_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6457_ (.I0(\registers[16][27] ),
    .I1(\registers[17][27] ),
    .S(_2910_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6458_ (.I0(\registers[18][27] ),
    .I1(\registers[19][27] ),
    .S(_2912_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6459_ (.I0(\registers[20][27] ),
    .I1(\registers[21][27] ),
    .S(_2863_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6460_ (.I0(\registers[22][27] ),
    .I1(\registers[23][27] ),
    .S(_2915_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6461_ (.I0(_2988_),
    .I1(_2989_),
    .I2(_2990_),
    .I3(_2991_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6462_ (.A1(_2831_),
    .A2(_2987_),
    .B1(_2992_),
    .B2(_2840_),
    .C(_2763_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6463_ (.A1(net99),
    .A2(_2765_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6464_ (.A1(_2984_),
    .A2(_2993_),
    .B(_2994_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6465_ (.I(_2431_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6466_ (.I0(\registers[28][28] ),
    .I1(\registers[29][28] ),
    .I2(\registers[30][28] ),
    .I3(\registers[31][28] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6467_ (.I(_2439_),
    .Z(_2997_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6468_ (.I0(\registers[24][28] ),
    .I1(\registers[25][28] ),
    .I2(\registers[26][28] ),
    .I3(\registers[27][28] ),
    .S0(_2997_),
    .S1(_2792_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6469_ (.I0(_2996_),
    .I1(_2998_),
    .S(_2946_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6470_ (.I(_2448_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6471_ (.I(_2450_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6472_ (.I0(\registers[18][28] ),
    .I1(\registers[19][28] ),
    .S(_3001_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6473_ (.I(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6474_ (.I(_2454_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6475_ (.I0(\registers[16][28] ),
    .I1(\registers[17][28] ),
    .S(_2950_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6476_ (.I0(\registers[22][28] ),
    .I1(\registers[23][28] ),
    .S(_2926_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6477_ (.I(_2458_),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6478_ (.A1(_3004_),
    .A2(_3005_),
    .B1(_3006_),
    .B2(_3007_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6479_ (.A1(_3000_),
    .A2(_3003_),
    .B(_3008_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6480_ (.I(_2464_),
    .Z(_3010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6481_ (.I0(\registers[20][28] ),
    .I1(\registers[21][28] ),
    .S(_2955_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6482_ (.I(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6483_ (.A1(_3010_),
    .A2(_3012_),
    .B(_2958_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6484_ (.A1(_2995_),
    .A2(_2999_),
    .B1(_3009_),
    .B2(_3013_),
    .C(_2472_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6485_ (.I0(\registers[12][28] ),
    .I1(\registers[13][28] ),
    .I2(\registers[14][28] ),
    .I3(\registers[15][28] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6486_ (.I0(\registers[8][28] ),
    .I1(\registers[9][28] ),
    .I2(\registers[10][28] ),
    .I3(\registers[11][28] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6487_ (.I(_2444_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6488_ (.I0(_3015_),
    .I1(_3016_),
    .S(_3017_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6489_ (.I0(\registers[0][28] ),
    .I1(\registers[1][28] ),
    .S(_2910_),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6490_ (.I0(\registers[2][28] ),
    .I1(\registers[3][28] ),
    .S(_2912_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6491_ (.I0(\registers[4][28] ),
    .I1(\registers[5][28] ),
    .S(_2863_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6492_ (.I0(\registers[6][28] ),
    .I1(\registers[7][28] ),
    .S(_2915_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6493_ (.I0(_3019_),
    .I1(_3020_),
    .I2(_3021_),
    .I3(_3022_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6494_ (.I(_2494_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6495_ (.A1(_2475_),
    .A2(_3018_),
    .B1(_3023_),
    .B2(_2485_),
    .C(_3024_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6496_ (.I(_2498_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6497_ (.A1(net100),
    .A2(_3026_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6498_ (.A1(_3014_),
    .A2(_3025_),
    .B(_3027_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6499_ (.I0(\registers[12][29] ),
    .I1(\registers[13][29] ),
    .I2(\registers[14][29] ),
    .I3(\registers[15][29] ),
    .S0(_2790_),
    .S1(_2843_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6500_ (.I0(\registers[8][29] ),
    .I1(\registers[9][29] ),
    .I2(\registers[10][29] ),
    .I3(\registers[11][29] ),
    .S0(_2997_),
    .S1(_2792_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6501_ (.I0(_3028_),
    .I1(_3029_),
    .S(_2946_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6502_ (.I0(\registers[2][29] ),
    .I1(\registers[3][29] ),
    .S(_3001_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6503_ (.I(_3031_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6504_ (.I0(\registers[0][29] ),
    .I1(\registers[1][29] ),
    .S(_2950_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6505_ (.I0(\registers[6][29] ),
    .I1(\registers[7][29] ),
    .S(_2926_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6506_ (.A1(_3004_),
    .A2(_3033_),
    .B1(_3034_),
    .B2(_3007_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6507_ (.A1(_3000_),
    .A2(_3032_),
    .B(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6508_ (.I0(\registers[4][29] ),
    .I1(\registers[5][29] ),
    .S(_2955_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6509_ (.I(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6510_ (.A1(_3010_),
    .A2(_3038_),
    .B(_2958_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6511_ (.A1(_2995_),
    .A2(_3030_),
    .B1(_3036_),
    .B2(_3039_),
    .C(_2829_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6512_ (.I0(\registers[28][29] ),
    .I1(\registers[29][29] ),
    .I2(\registers[30][29] ),
    .I3(\registers[31][29] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6513_ (.I0(\registers[24][29] ),
    .I1(\registers[25][29] ),
    .I2(\registers[26][29] ),
    .I3(\registers[27][29] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6514_ (.I0(_3041_),
    .I1(_3042_),
    .S(_3017_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6515_ (.I0(\registers[16][29] ),
    .I1(\registers[17][29] ),
    .S(_2910_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6516_ (.I0(\registers[18][29] ),
    .I1(\registers[19][29] ),
    .S(_2912_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6517_ (.I0(\registers[20][29] ),
    .I1(\registers[21][29] ),
    .S(_2863_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6518_ (.I0(\registers[22][29] ),
    .I1(\registers[23][29] ),
    .S(_2915_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6519_ (.I0(_3044_),
    .I1(_3045_),
    .I2(_3046_),
    .I3(_3047_),
    .S0(_2812_),
    .S1(_2813_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6520_ (.A1(_2831_),
    .A2(_3043_),
    .B1(_3048_),
    .B2(_2840_),
    .C(_3024_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6521_ (.A1(net101),
    .A2(_3026_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6522_ (.A1(_3040_),
    .A2(_3049_),
    .B(_3050_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6523_ (.I(_2434_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6524_ (.I0(\registers[28][2] ),
    .I1(\registers[29][2] ),
    .I2(\registers[30][2] ),
    .I3(\registers[31][2] ),
    .S0(_3051_),
    .S1(_2843_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6525_ (.I(_2436_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6526_ (.I0(\registers[24][2] ),
    .I1(\registers[25][2] ),
    .I2(\registers[26][2] ),
    .I3(\registers[27][2] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6527_ (.I0(_3052_),
    .I1(_3054_),
    .S(_2946_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6528_ (.I0(\registers[18][2] ),
    .I1(\registers[19][2] ),
    .S(_3001_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6529_ (.I(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6530_ (.I0(\registers[16][2] ),
    .I1(\registers[17][2] ),
    .S(_2950_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6531_ (.I0(\registers[22][2] ),
    .I1(\registers[23][2] ),
    .S(_2926_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6532_ (.A1(_3004_),
    .A2(_3058_),
    .B1(_3059_),
    .B2(_3007_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6533_ (.A1(_3000_),
    .A2(_3057_),
    .B(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6534_ (.I0(\registers[20][2] ),
    .I1(\registers[21][2] ),
    .S(_2955_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6535_ (.I(_3062_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6536_ (.A1(_3010_),
    .A2(_3063_),
    .B(_2958_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6537_ (.A1(_2995_),
    .A2(_3055_),
    .B1(_3061_),
    .B2(_3064_),
    .C(_2472_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6538_ (.I0(\registers[12][2] ),
    .I1(\registers[13][2] ),
    .I2(\registers[14][2] ),
    .I3(\registers[15][2] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6539_ (.I0(\registers[8][2] ),
    .I1(\registers[9][2] ),
    .I2(\registers[10][2] ),
    .I3(\registers[11][2] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6540_ (.I0(_3066_),
    .I1(_3067_),
    .S(_3017_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6541_ (.I0(\registers[0][2] ),
    .I1(\registers[1][2] ),
    .S(_2910_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6542_ (.I0(\registers[2][2] ),
    .I1(\registers[3][2] ),
    .S(_2912_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6543_ (.I0(\registers[4][2] ),
    .I1(\registers[5][2] ),
    .S(_2863_),
    .Z(_3071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6544_ (.I0(\registers[6][2] ),
    .I1(\registers[7][2] ),
    .S(_2915_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _6545_ (.I(_2447_),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6546_ (.I(net4),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6547_ (.I0(_3069_),
    .I1(_3070_),
    .I2(_3071_),
    .I3(_3072_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6548_ (.A1(_2475_),
    .A2(_3068_),
    .B1(_3075_),
    .B2(_2485_),
    .C(_3024_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6549_ (.A1(net102),
    .A2(_3026_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6550_ (.A1(_3065_),
    .A2(_3076_),
    .B(_3077_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6551_ (.I0(\registers[12][30] ),
    .I1(\registers[13][30] ),
    .I2(\registers[14][30] ),
    .I3(\registers[15][30] ),
    .S0(_3051_),
    .S1(_2843_),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6552_ (.I0(\registers[8][30] ),
    .I1(\registers[9][30] ),
    .I2(\registers[10][30] ),
    .I3(\registers[11][30] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6553_ (.I0(_3078_),
    .I1(_3079_),
    .S(_2946_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6554_ (.I0(\registers[2][30] ),
    .I1(\registers[3][30] ),
    .S(_3001_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6555_ (.I(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6556_ (.I0(\registers[0][30] ),
    .I1(\registers[1][30] ),
    .S(_2950_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6557_ (.I0(\registers[6][30] ),
    .I1(\registers[7][30] ),
    .S(_2926_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6558_ (.A1(_3004_),
    .A2(_3083_),
    .B1(_3084_),
    .B2(_3007_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6559_ (.A1(_3000_),
    .A2(_3082_),
    .B(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6560_ (.I0(\registers[4][30] ),
    .I1(\registers[5][30] ),
    .S(_2955_),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6561_ (.I(_3087_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6562_ (.A1(_3010_),
    .A2(_3088_),
    .B(_2958_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6563_ (.A1(_2995_),
    .A2(_3080_),
    .B1(_3086_),
    .B2(_3089_),
    .C(_2829_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6564_ (.I0(\registers[28][30] ),
    .I1(\registers[29][30] ),
    .I2(\registers[30][30] ),
    .I3(\registers[31][30] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6565_ (.I0(\registers[24][30] ),
    .I1(\registers[25][30] ),
    .I2(\registers[26][30] ),
    .I3(\registers[27][30] ),
    .S0(_2858_),
    .S1(_2907_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6566_ (.I0(_3091_),
    .I1(_3092_),
    .S(_3017_),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6567_ (.I0(\registers[16][30] ),
    .I1(\registers[17][30] ),
    .S(_2910_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6568_ (.I0(\registers[18][30] ),
    .I1(\registers[19][30] ),
    .S(_2912_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6569_ (.I0(\registers[20][30] ),
    .I1(\registers[21][30] ),
    .S(_2863_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6570_ (.I0(\registers[22][30] ),
    .I1(\registers[23][30] ),
    .S(_2915_),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6571_ (.I0(_3094_),
    .I1(_3095_),
    .I2(_3096_),
    .I3(_3097_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6572_ (.A1(_2831_),
    .A2(_3093_),
    .B1(_3098_),
    .B2(_2840_),
    .C(_3024_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6573_ (.A1(net103),
    .A2(_3026_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6574_ (.A1(_3090_),
    .A2(_3099_),
    .B(_3100_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6575_ (.I0(\registers[28][31] ),
    .I1(\registers[29][31] ),
    .I2(\registers[30][31] ),
    .I3(\registers[31][31] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6576_ (.I0(\registers[24][31] ),
    .I1(\registers[25][31] ),
    .I2(\registers[26][31] ),
    .I3(\registers[27][31] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6577_ (.I0(_3101_),
    .I1(_3102_),
    .S(_2946_),
    .Z(_3103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6578_ (.I0(\registers[18][31] ),
    .I1(\registers[19][31] ),
    .S(_3001_),
    .Z(_3104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6579_ (.I(_3104_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6580_ (.I0(\registers[16][31] ),
    .I1(\registers[17][31] ),
    .S(_2950_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6581_ (.I0(\registers[22][31] ),
    .I1(\registers[23][31] ),
    .S(_2926_),
    .Z(_3107_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6582_ (.A1(_3004_),
    .A2(_3106_),
    .B1(_3107_),
    .B2(_3007_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6583_ (.A1(_3000_),
    .A2(_3105_),
    .B(_3108_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6584_ (.I0(\registers[20][31] ),
    .I1(\registers[21][31] ),
    .S(_2955_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6585_ (.I(_3110_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6586_ (.A1(_3010_),
    .A2(_3111_),
    .B(_2958_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6587_ (.A1(_2995_),
    .A2(_3103_),
    .B1(_3109_),
    .B2(_3112_),
    .C(_2472_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6588_ (.I0(\registers[12][31] ),
    .I1(\registers[13][31] ),
    .I2(\registers[14][31] ),
    .I3(\registers[15][31] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6589_ (.I0(\registers[8][31] ),
    .I1(\registers[9][31] ),
    .I2(\registers[10][31] ),
    .I3(\registers[11][31] ),
    .S0(_2435_),
    .S1(_2907_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6590_ (.I0(_3114_),
    .I1(_3115_),
    .S(_3017_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6591_ (.I0(\registers[0][31] ),
    .I1(\registers[1][31] ),
    .S(_2910_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6592_ (.I0(\registers[2][31] ),
    .I1(\registers[3][31] ),
    .S(_2912_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6593_ (.I0(\registers[4][31] ),
    .I1(\registers[5][31] ),
    .S(_2486_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6594_ (.I0(\registers[6][31] ),
    .I1(\registers[7][31] ),
    .S(_2915_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6595_ (.I0(_3117_),
    .I1(_3118_),
    .I2(_3119_),
    .I3(_3120_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3121_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6596_ (.A1(_2475_),
    .A2(_3116_),
    .B1(_3121_),
    .B2(_2485_),
    .C(_3024_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6597_ (.A1(net104),
    .A2(_3026_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6598_ (.A1(_3113_),
    .A2(_3122_),
    .B(_3123_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6599_ (.I0(\registers[12][3] ),
    .I1(\registers[13][3] ),
    .I2(\registers[14][3] ),
    .I3(\registers[15][3] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6600_ (.I0(\registers[8][3] ),
    .I1(\registers[9][3] ),
    .I2(\registers[10][3] ),
    .I3(\registers[11][3] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6601_ (.I0(_3124_),
    .I1(_3125_),
    .S(_2946_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6602_ (.I0(\registers[2][3] ),
    .I1(\registers[3][3] ),
    .S(_3001_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6603_ (.I(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6604_ (.I0(\registers[0][3] ),
    .I1(\registers[1][3] ),
    .S(_2950_),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6605_ (.I0(\registers[6][3] ),
    .I1(\registers[7][3] ),
    .S(_2926_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6606_ (.A1(_3004_),
    .A2(_3129_),
    .B1(_3130_),
    .B2(_3007_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6607_ (.A1(_3000_),
    .A2(_3128_),
    .B(_3131_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6608_ (.I0(\registers[4][3] ),
    .I1(\registers[5][3] ),
    .S(_2955_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6609_ (.I(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6610_ (.A1(_3010_),
    .A2(_3134_),
    .B(_2958_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6611_ (.A1(_2995_),
    .A2(_3126_),
    .B1(_3132_),
    .B2(_3135_),
    .C(_2829_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6612_ (.I0(\registers[28][3] ),
    .I1(\registers[29][3] ),
    .I2(\registers[30][3] ),
    .I3(\registers[31][3] ),
    .S0(_2905_),
    .S1(_2961_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6613_ (.I0(\registers[24][3] ),
    .I1(\registers[25][3] ),
    .I2(\registers[26][3] ),
    .I3(\registers[27][3] ),
    .S0(_2435_),
    .S1(_2907_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6614_ (.I0(_3137_),
    .I1(_3138_),
    .S(_3017_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6615_ (.I0(\registers[16][3] ),
    .I1(\registers[17][3] ),
    .S(_2910_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6616_ (.I0(\registers[18][3] ),
    .I1(\registers[19][3] ),
    .S(_2912_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6617_ (.I0(\registers[20][3] ),
    .I1(\registers[21][3] ),
    .S(_2486_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6618_ (.I0(\registers[22][3] ),
    .I1(\registers[23][3] ),
    .S(_2915_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6619_ (.I0(_3140_),
    .I1(_3141_),
    .I2(_3142_),
    .I3(_3143_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6620_ (.A1(_2831_),
    .A2(_3139_),
    .B1(_3144_),
    .B2(_2840_),
    .C(_3024_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6621_ (.A1(net105),
    .A2(_3026_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6622_ (.A1(_3136_),
    .A2(_3145_),
    .B(_3146_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6623_ (.I0(\registers[28][4] ),
    .I1(\registers[29][4] ),
    .I2(\registers[30][4] ),
    .I3(\registers[31][4] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6624_ (.I0(\registers[24][4] ),
    .I1(\registers[25][4] ),
    .I2(\registers[26][4] ),
    .I3(\registers[27][4] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6625_ (.I0(_3147_),
    .I1(_3148_),
    .S(_2946_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6626_ (.I0(\registers[18][4] ),
    .I1(\registers[19][4] ),
    .S(_3001_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6627_ (.I(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6628_ (.I0(\registers[16][4] ),
    .I1(\registers[17][4] ),
    .S(_2950_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6629_ (.I0(\registers[22][4] ),
    .I1(\registers[23][4] ),
    .S(_2926_),
    .Z(_3153_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6630_ (.A1(_3004_),
    .A2(_3152_),
    .B1(_3153_),
    .B2(_3007_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6631_ (.A1(_3000_),
    .A2(_3151_),
    .B(_3154_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6632_ (.I0(\registers[20][4] ),
    .I1(\registers[21][4] ),
    .S(_2955_),
    .Z(_3156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6633_ (.I(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6634_ (.A1(_3010_),
    .A2(_3157_),
    .B(_2958_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6635_ (.A1(_2995_),
    .A2(_3149_),
    .B1(_3155_),
    .B2(_3158_),
    .C(_2471_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6636_ (.I0(\registers[12][4] ),
    .I1(\registers[13][4] ),
    .I2(\registers[14][4] ),
    .I3(\registers[15][4] ),
    .S0(_2479_),
    .S1(_2961_),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6637_ (.I0(\registers[8][4] ),
    .I1(\registers[9][4] ),
    .I2(\registers[10][4] ),
    .I3(\registers[11][4] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6638_ (.I0(_3160_),
    .I1(_3161_),
    .S(_3017_),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6639_ (.I0(\registers[0][4] ),
    .I1(\registers[1][4] ),
    .S(_2552_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6640_ (.I0(\registers[2][4] ),
    .I1(\registers[3][4] ),
    .S(_2548_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6641_ (.I0(\registers[4][4] ),
    .I1(\registers[5][4] ),
    .S(_2486_),
    .Z(_3165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6642_ (.I0(\registers[6][4] ),
    .I1(\registers[7][4] ),
    .S(_2489_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6643_ (.I0(_3163_),
    .I1(_3164_),
    .I2(_3165_),
    .I3(_3166_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6644_ (.A1(_2474_),
    .A2(_3162_),
    .B1(_3167_),
    .B2(_2484_),
    .C(_3024_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6645_ (.A1(net106),
    .A2(_3026_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6646_ (.A1(_3159_),
    .A2(_3168_),
    .B(_3169_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6647_ (.I0(\registers[12][5] ),
    .I1(\registers[13][5] ),
    .I2(\registers[14][5] ),
    .I3(\registers[15][5] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6648_ (.I0(\registers[8][5] ),
    .I1(\registers[9][5] ),
    .I2(\registers[10][5] ),
    .I3(\registers[11][5] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6649_ (.I0(_3170_),
    .I1(_3171_),
    .S(_2946_),
    .Z(_3172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6650_ (.I0(\registers[2][5] ),
    .I1(\registers[3][5] ),
    .S(_3001_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6651_ (.I(_3173_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6652_ (.I0(\registers[0][5] ),
    .I1(\registers[1][5] ),
    .S(_2950_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6653_ (.I0(\registers[6][5] ),
    .I1(\registers[7][5] ),
    .S(_2460_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6654_ (.A1(_3004_),
    .A2(_3175_),
    .B1(_3176_),
    .B2(_3007_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6655_ (.A1(_3000_),
    .A2(_3174_),
    .B(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6656_ (.I0(\registers[4][5] ),
    .I1(\registers[5][5] ),
    .S(_2955_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6657_ (.I(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6658_ (.A1(_3010_),
    .A2(_3180_),
    .B(_2958_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _6659_ (.A1(_2995_),
    .A2(_3172_),
    .B1(_3178_),
    .B2(_3181_),
    .C(_2829_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6660_ (.I0(\registers[28][5] ),
    .I1(\registers[29][5] ),
    .I2(\registers[30][5] ),
    .I3(\registers[31][5] ),
    .S0(_2479_),
    .S1(_2961_),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6661_ (.I0(\registers[24][5] ),
    .I1(\registers[25][5] ),
    .I2(\registers[26][5] ),
    .I3(\registers[27][5] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6662_ (.I0(_3183_),
    .I1(_3184_),
    .S(_3017_),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6663_ (.I0(\registers[16][5] ),
    .I1(\registers[17][5] ),
    .S(_2552_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6664_ (.I0(\registers[18][5] ),
    .I1(\registers[19][5] ),
    .S(_2548_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6665_ (.I0(\registers[20][5] ),
    .I1(\registers[21][5] ),
    .S(_2486_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6666_ (.I0(\registers[22][5] ),
    .I1(\registers[23][5] ),
    .S(_2489_),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6667_ (.I0(_3186_),
    .I1(_3187_),
    .I2(_3188_),
    .I3(_3189_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6668_ (.A1(_2831_),
    .A2(_3185_),
    .B1(_3190_),
    .B2(_2840_),
    .C(_3024_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6669_ (.A1(net107),
    .A2(_3026_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6670_ (.A1(_3182_),
    .A2(_3191_),
    .B(_3192_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6671_ (.I0(\registers[28][6] ),
    .I1(\registers[29][6] ),
    .I2(\registers[30][6] ),
    .I3(\registers[31][6] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6672_ (.I0(\registers[24][6] ),
    .I1(\registers[25][6] ),
    .I2(\registers[26][6] ),
    .I3(\registers[27][6] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6673_ (.I0(_3193_),
    .I1(_3194_),
    .S(_2444_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6674_ (.I0(\registers[18][6] ),
    .I1(\registers[19][6] ),
    .S(_3001_),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6675_ (.I(_3196_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6676_ (.I0(\registers[16][6] ),
    .I1(\registers[17][6] ),
    .S(_2507_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6677_ (.I0(\registers[22][6] ),
    .I1(\registers[23][6] ),
    .S(_2460_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6678_ (.A1(_3004_),
    .A2(_3198_),
    .B1(_3199_),
    .B2(_3007_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6679_ (.A1(_3000_),
    .A2(_3197_),
    .B(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6680_ (.I0(\registers[20][6] ),
    .I1(\registers[21][6] ),
    .S(_2476_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6681_ (.I(_3202_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6682_ (.A1(_3010_),
    .A2(_3203_),
    .B(_2431_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _6683_ (.A1(_2995_),
    .A2(_3195_),
    .B1(_3201_),
    .B2(_3204_),
    .C(_2471_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6684_ (.I0(\registers[12][6] ),
    .I1(\registers[13][6] ),
    .I2(\registers[14][6] ),
    .I3(\registers[15][6] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6685_ (.I0(\registers[8][6] ),
    .I1(\registers[9][6] ),
    .I2(\registers[10][6] ),
    .I3(\registers[11][6] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6686_ (.I0(_3206_),
    .I1(_3207_),
    .S(_3017_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6687_ (.I0(\registers[0][6] ),
    .I1(\registers[1][6] ),
    .S(_2552_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6688_ (.I0(\registers[2][6] ),
    .I1(\registers[3][6] ),
    .S(_2548_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6689_ (.I0(\registers[4][6] ),
    .I1(\registers[5][6] ),
    .S(_2486_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6690_ (.I0(\registers[6][6] ),
    .I1(\registers[7][6] ),
    .S(_2489_),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6691_ (.I0(_3209_),
    .I1(_3210_),
    .I2(_3211_),
    .I3(_3212_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6692_ (.A1(_2474_),
    .A2(_3208_),
    .B1(_3213_),
    .B2(_2484_),
    .C(_3024_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6693_ (.A1(net108),
    .A2(_3026_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6694_ (.A1(_3205_),
    .A2(_3214_),
    .B(_3215_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6695_ (.I0(\registers[12][7] ),
    .I1(\registers[13][7] ),
    .I2(\registers[14][7] ),
    .I3(\registers[15][7] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6696_ (.I0(\registers[8][7] ),
    .I1(\registers[9][7] ),
    .I2(\registers[10][7] ),
    .I3(\registers[11][7] ),
    .S0(_2997_),
    .S1(_3053_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6697_ (.I0(_3216_),
    .I1(_3217_),
    .S(_2444_),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6698_ (.I0(\registers[2][7] ),
    .I1(\registers[3][7] ),
    .S(_3001_),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6699_ (.I(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6700_ (.I0(\registers[0][7] ),
    .I1(\registers[1][7] ),
    .S(_2507_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6701_ (.I0(\registers[6][7] ),
    .I1(\registers[7][7] ),
    .S(_2460_),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6702_ (.A1(_3004_),
    .A2(_3221_),
    .B1(_3222_),
    .B2(_3007_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6703_ (.A1(_3000_),
    .A2(_3220_),
    .B(_3223_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6704_ (.I0(\registers[4][7] ),
    .I1(\registers[5][7] ),
    .S(_2476_),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6705_ (.I(_3225_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6706_ (.A1(_3010_),
    .A2(_3226_),
    .B(_2431_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _6707_ (.A1(_2995_),
    .A2(_3218_),
    .B1(_3224_),
    .B2(_3227_),
    .C(_2829_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6708_ (.I0(\registers[28][7] ),
    .I1(\registers[29][7] ),
    .I2(\registers[30][7] ),
    .I3(\registers[31][7] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6709_ (.I0(\registers[24][7] ),
    .I1(\registers[25][7] ),
    .I2(\registers[26][7] ),
    .I3(\registers[27][7] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6710_ (.I0(_3229_),
    .I1(_3230_),
    .S(_3017_),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6711_ (.I0(\registers[16][7] ),
    .I1(\registers[17][7] ),
    .S(_2552_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6712_ (.I0(\registers[18][7] ),
    .I1(\registers[19][7] ),
    .S(_2548_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6713_ (.I0(\registers[20][7] ),
    .I1(\registers[21][7] ),
    .S(_2486_),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6714_ (.I0(\registers[22][7] ),
    .I1(\registers[23][7] ),
    .S(_2489_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6715_ (.I0(_3232_),
    .I1(_3233_),
    .I2(_3234_),
    .I3(_3235_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6716_ (.A1(_2831_),
    .A2(_3231_),
    .B1(_3236_),
    .B2(_2840_),
    .C(_3024_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6717_ (.A1(net109),
    .A2(_3026_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6718_ (.A1(_3228_),
    .A2(_3237_),
    .B(_3238_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6719_ (.I0(\registers[12][8] ),
    .I1(\registers[13][8] ),
    .I2(\registers[14][8] ),
    .I3(\registers[15][8] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6720_ (.I0(\registers[8][8] ),
    .I1(\registers[9][8] ),
    .I2(\registers[10][8] ),
    .I3(\registers[11][8] ),
    .S0(_2456_),
    .S1(_3053_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6721_ (.I0(_3239_),
    .I1(_3240_),
    .S(_2444_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6722_ (.I0(\registers[2][8] ),
    .I1(\registers[3][8] ),
    .S(_2466_),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6723_ (.I(_3242_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6724_ (.I0(\registers[0][8] ),
    .I1(\registers[1][8] ),
    .S(_2507_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6725_ (.I0(\registers[6][8] ),
    .I1(\registers[7][8] ),
    .S(_2460_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6726_ (.A1(_2454_),
    .A2(_3244_),
    .B1(_3245_),
    .B2(_2458_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6727_ (.A1(_2448_),
    .A2(_3243_),
    .B(_3246_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6728_ (.I0(\registers[4][8] ),
    .I1(\registers[5][8] ),
    .S(_2476_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6729_ (.I(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6730_ (.A1(_2464_),
    .A2(_3249_),
    .B(_2431_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _6731_ (.A1(_2469_),
    .A2(_3241_),
    .B1(_3247_),
    .B2(_3250_),
    .C(_2829_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6732_ (.I0(\registers[28][8] ),
    .I1(\registers[29][8] ),
    .I2(\registers[30][8] ),
    .I3(\registers[31][8] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6733_ (.I0(\registers[24][8] ),
    .I1(\registers[25][8] ),
    .I2(\registers[26][8] ),
    .I3(\registers[27][8] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6734_ (.I0(_3252_),
    .I1(_3253_),
    .S(_2445_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6735_ (.I0(\registers[16][8] ),
    .I1(\registers[17][8] ),
    .S(_2552_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6736_ (.I0(\registers[18][8] ),
    .I1(\registers[19][8] ),
    .S(_2548_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6737_ (.I0(\registers[20][8] ),
    .I1(\registers[21][8] ),
    .S(_2486_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6738_ (.I0(\registers[22][8] ),
    .I1(\registers[23][8] ),
    .S(_2489_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6739_ (.I0(_3255_),
    .I1(_3256_),
    .I2(_3257_),
    .I3(_3258_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6740_ (.A1(_2831_),
    .A2(_3254_),
    .B1(_3259_),
    .B2(_2840_),
    .C(_2494_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6741_ (.A1(net110),
    .A2(_2498_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6742_ (.A1(_3251_),
    .A2(_3260_),
    .B(_3261_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6743_ (.I0(\registers[12][9] ),
    .I1(\registers[13][9] ),
    .I2(\registers[14][9] ),
    .I3(\registers[15][9] ),
    .S0(_3051_),
    .S1(_2441_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6744_ (.I0(\registers[8][9] ),
    .I1(\registers[9][9] ),
    .I2(\registers[10][9] ),
    .I3(\registers[11][9] ),
    .S0(_2456_),
    .S1(_3053_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6745_ (.I0(_3262_),
    .I1(_3263_),
    .S(_2444_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6746_ (.I0(\registers[2][9] ),
    .I1(\registers[3][9] ),
    .S(_2466_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6747_ (.I(_3265_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6748_ (.I0(\registers[0][9] ),
    .I1(\registers[1][9] ),
    .S(_2507_),
    .Z(_3267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6749_ (.I0(\registers[6][9] ),
    .I1(\registers[7][9] ),
    .S(_2460_),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _6750_ (.A1(_2454_),
    .A2(_3267_),
    .B1(_3268_),
    .B2(_2458_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6751_ (.A1(_2448_),
    .A2(_3266_),
    .B(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6752_ (.I0(\registers[4][9] ),
    .I1(\registers[5][9] ),
    .S(_2476_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _6753_ (.I(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6754_ (.A1(_2464_),
    .A2(_3272_),
    .B(_2431_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _6755_ (.A1(_2469_),
    .A2(_3264_),
    .B1(_3270_),
    .B2(_3273_),
    .C(_2829_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6756_ (.I0(\registers[28][9] ),
    .I1(\registers[29][9] ),
    .I2(\registers[30][9] ),
    .I3(\registers[31][9] ),
    .S0(_2479_),
    .S1(_2480_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6757_ (.I0(\registers[24][9] ),
    .I1(\registers[25][9] ),
    .I2(\registers[26][9] ),
    .I3(\registers[27][9] ),
    .S0(_2435_),
    .S1(_2437_),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6758_ (.I0(_3275_),
    .I1(_3276_),
    .S(_2445_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6759_ (.I0(\registers[16][9] ),
    .I1(\registers[17][9] ),
    .S(_2552_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6760_ (.I0(\registers[18][9] ),
    .I1(\registers[19][9] ),
    .S(_2548_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6761_ (.I0(\registers[20][9] ),
    .I1(\registers[21][9] ),
    .S(_2486_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6762_ (.I0(\registers[22][9] ),
    .I1(\registers[23][9] ),
    .S(_2489_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _6763_ (.I0(_3278_),
    .I1(_3279_),
    .I2(_3280_),
    .I3(_3281_),
    .S0(_3073_),
    .S1(_3074_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _6764_ (.A1(_2831_),
    .A2(_3277_),
    .B1(_3282_),
    .B2(_2840_),
    .C(_2494_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6765_ (.A1(net111),
    .A2(_2498_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _6766_ (.A1(_3274_),
    .A2(_3283_),
    .B(_3284_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6767_ (.A1(_1532_),
    .A2(\registers[0][0] ),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _6768_ (.A1(_1116_),
    .A2(_1338_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6769_ (.I(_3286_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6770_ (.I0(_1229_),
    .I1(_3285_),
    .S(_3287_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6771_ (.A1(_1532_),
    .A2(\registers[0][10] ),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6772_ (.I0(_1235_),
    .I1(_3288_),
    .S(_3287_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6773_ (.A1(_1532_),
    .A2(\registers[0][11] ),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6774_ (.I0(_1237_),
    .I1(_3289_),
    .S(_3287_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6775_ (.A1(_1532_),
    .A2(\registers[0][12] ),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6776_ (.I0(_1239_),
    .I1(_3290_),
    .S(_3287_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6777_ (.A1(_1532_),
    .A2(\registers[0][13] ),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6778_ (.I0(_1241_),
    .I1(_3291_),
    .S(_3287_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6779_ (.A1(_1532_),
    .A2(\registers[0][14] ),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6780_ (.I0(_1243_),
    .I1(_3292_),
    .S(_3287_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6781_ (.I(_1455_),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6782_ (.A1(_3293_),
    .A2(\registers[0][15] ),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6783_ (.I0(_1245_),
    .I1(_3294_),
    .S(_3287_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6784_ (.A1(_3293_),
    .A2(\registers[0][16] ),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6785_ (.I0(_1247_),
    .I1(_3295_),
    .S(_3287_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6786_ (.A1(_3293_),
    .A2(\registers[0][17] ),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6787_ (.I0(_1249_),
    .I1(_3296_),
    .S(_3287_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6788_ (.A1(_3293_),
    .A2(\registers[0][18] ),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6789_ (.I0(_1251_),
    .I1(_3297_),
    .S(_3287_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6790_ (.A1(_3293_),
    .A2(\registers[0][19] ),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6791_ (.I(_3286_),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6792_ (.I0(_1253_),
    .I1(_3298_),
    .S(_3299_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6793_ (.A1(_3293_),
    .A2(\registers[0][1] ),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6794_ (.I0(_1257_),
    .I1(_3300_),
    .S(_3299_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6795_ (.A1(_3293_),
    .A2(\registers[0][20] ),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6796_ (.I0(_1259_),
    .I1(_3301_),
    .S(_3299_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6797_ (.A1(_3293_),
    .A2(\registers[0][21] ),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6798_ (.I0(_1261_),
    .I1(_3302_),
    .S(_3299_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6799_ (.A1(_3293_),
    .A2(\registers[0][22] ),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6800_ (.I0(_1263_),
    .I1(_3303_),
    .S(_3299_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6801_ (.A1(_3293_),
    .A2(\registers[0][23] ),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6802_ (.I0(_1265_),
    .I1(_3304_),
    .S(_3299_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6803_ (.I(_1455_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6804_ (.A1(_3305_),
    .A2(\registers[0][24] ),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6805_ (.I0(_1267_),
    .I1(_3306_),
    .S(_3299_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6806_ (.A1(_3305_),
    .A2(\registers[0][25] ),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6807_ (.I0(_1269_),
    .I1(_3307_),
    .S(_3299_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6808_ (.A1(_3305_),
    .A2(\registers[0][26] ),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6809_ (.I0(_1271_),
    .I1(_3308_),
    .S(_3299_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6810_ (.A1(_3305_),
    .A2(\registers[0][27] ),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6811_ (.I0(_1273_),
    .I1(_3309_),
    .S(_3299_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6812_ (.A1(_3305_),
    .A2(\registers[0][28] ),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6813_ (.I(_3286_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6814_ (.I0(_1275_),
    .I1(_3310_),
    .S(_3311_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6815_ (.A1(_3305_),
    .A2(\registers[0][29] ),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6816_ (.I0(_1279_),
    .I1(_3312_),
    .S(_3311_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6817_ (.A1(_3305_),
    .A2(\registers[0][2] ),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6818_ (.I0(_1281_),
    .I1(_3313_),
    .S(_3311_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6819_ (.A1(_3305_),
    .A2(\registers[0][30] ),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6820_ (.I0(_1283_),
    .I1(_3314_),
    .S(_3311_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6821_ (.A1(_3305_),
    .A2(\registers[0][31] ),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6822_ (.I0(_1088_),
    .I1(_3315_),
    .S(_3311_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6823_ (.A1(_3305_),
    .A2(\registers[0][3] ),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6824_ (.I0(_1098_),
    .I1(_3316_),
    .S(_3311_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6825_ (.I(_1455_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6826_ (.A1(_3317_),
    .A2(\registers[0][4] ),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6827_ (.I0(_1100_),
    .I1(_3318_),
    .S(_3311_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6828_ (.A1(_3317_),
    .A2(\registers[0][5] ),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6829_ (.I0(_1102_),
    .I1(_3319_),
    .S(_3311_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6830_ (.A1(_3317_),
    .A2(\registers[0][6] ),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6831_ (.I0(_1104_),
    .I1(_3320_),
    .S(_3311_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6832_ (.A1(_3317_),
    .A2(\registers[0][7] ),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6833_ (.I0(_1106_),
    .I1(_3321_),
    .S(_3311_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6834_ (.A1(_3317_),
    .A2(\registers[0][8] ),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6835_ (.I0(_1108_),
    .I1(_3322_),
    .S(_3286_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6836_ (.A1(_3317_),
    .A2(\registers[0][9] ),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6837_ (.I0(_1110_),
    .I1(_3323_),
    .S(_3286_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6838_ (.A1(_3317_),
    .A2(\registers[10][0] ),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _6839_ (.A1(_1119_),
    .A2(_1498_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6840_ (.I(_3325_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6841_ (.I0(_1229_),
    .I1(_3324_),
    .S(_3326_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6842_ (.A1(_3317_),
    .A2(\registers[10][10] ),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6843_ (.I0(_1235_),
    .I1(_3327_),
    .S(_3326_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6844_ (.A1(_3317_),
    .A2(\registers[10][11] ),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6845_ (.I0(_1237_),
    .I1(_3328_),
    .S(_3326_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6846_ (.A1(_3317_),
    .A2(\registers[10][12] ),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6847_ (.I0(_1239_),
    .I1(_3329_),
    .S(_3326_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6848_ (.I(_1089_),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6849_ (.I(_3330_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6850_ (.A1(_3331_),
    .A2(\registers[10][13] ),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6851_ (.I0(_1241_),
    .I1(_3332_),
    .S(_3326_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6852_ (.A1(_3331_),
    .A2(\registers[10][14] ),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6853_ (.I0(_1243_),
    .I1(_3333_),
    .S(_3326_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6854_ (.A1(_3331_),
    .A2(\registers[10][15] ),
    .Z(_3334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6855_ (.I0(_1245_),
    .I1(_3334_),
    .S(_3326_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6856_ (.A1(_3331_),
    .A2(\registers[10][16] ),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6857_ (.I0(_1247_),
    .I1(_3335_),
    .S(_3326_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6858_ (.A1(_3331_),
    .A2(\registers[10][17] ),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6859_ (.I0(_1249_),
    .I1(_3336_),
    .S(_3326_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6860_ (.A1(_3331_),
    .A2(\registers[10][18] ),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6861_ (.I0(_1251_),
    .I1(_3337_),
    .S(_3326_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6862_ (.A1(_3331_),
    .A2(\registers[10][19] ),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6863_ (.I(_3325_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6864_ (.I0(_1253_),
    .I1(_3338_),
    .S(_3339_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6865_ (.A1(_3331_),
    .A2(\registers[10][1] ),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6866_ (.I0(_1257_),
    .I1(_3340_),
    .S(_3339_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6867_ (.A1(_3331_),
    .A2(\registers[10][20] ),
    .Z(_3341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6868_ (.I0(_1259_),
    .I1(_3341_),
    .S(_3339_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6869_ (.A1(_3331_),
    .A2(\registers[10][21] ),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6870_ (.I0(_1261_),
    .I1(_3342_),
    .S(_3339_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6871_ (.I(_3330_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6872_ (.A1(_3343_),
    .A2(\registers[10][22] ),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6873_ (.I0(_1263_),
    .I1(_3344_),
    .S(_3339_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6874_ (.A1(_3343_),
    .A2(\registers[10][23] ),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6875_ (.I0(_1265_),
    .I1(_3345_),
    .S(_3339_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6876_ (.A1(_3343_),
    .A2(\registers[10][24] ),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6877_ (.I0(_1267_),
    .I1(_3346_),
    .S(_3339_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6878_ (.A1(_3343_),
    .A2(\registers[10][25] ),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6879_ (.I0(_1269_),
    .I1(_3347_),
    .S(_3339_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6880_ (.A1(_3343_),
    .A2(\registers[10][26] ),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6881_ (.I0(_1271_),
    .I1(_3348_),
    .S(_3339_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6882_ (.A1(_3343_),
    .A2(\registers[10][27] ),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6883_ (.I0(_1273_),
    .I1(_3349_),
    .S(_3339_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6884_ (.A1(_3343_),
    .A2(\registers[10][28] ),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6885_ (.I(_3325_),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6886_ (.I0(_1275_),
    .I1(_3350_),
    .S(_3351_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6887_ (.A1(_3343_),
    .A2(\registers[10][29] ),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6888_ (.I0(_1279_),
    .I1(_3352_),
    .S(_3351_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6889_ (.A1(_3343_),
    .A2(\registers[10][2] ),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6890_ (.I0(_1281_),
    .I1(_3353_),
    .S(_3351_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6891_ (.A1(_3343_),
    .A2(\registers[10][30] ),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6892_ (.I0(_1283_),
    .I1(_3354_),
    .S(_3351_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6893_ (.I(_3330_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6894_ (.A1(_3355_),
    .A2(\registers[10][31] ),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6895_ (.I0(_1088_),
    .I1(_3356_),
    .S(_3351_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6896_ (.A1(_3355_),
    .A2(\registers[10][3] ),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6897_ (.I0(_1098_),
    .I1(_3357_),
    .S(_3351_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6898_ (.A1(_3355_),
    .A2(\registers[10][4] ),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6899_ (.I0(_1100_),
    .I1(_3358_),
    .S(_3351_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6900_ (.A1(_3355_),
    .A2(\registers[10][5] ),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6901_ (.I0(_1102_),
    .I1(_3359_),
    .S(_3351_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6902_ (.A1(_3355_),
    .A2(\registers[10][6] ),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6903_ (.I0(_1104_),
    .I1(_3360_),
    .S(_3351_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6904_ (.A1(_3355_),
    .A2(\registers[10][7] ),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6905_ (.I0(_1106_),
    .I1(_3361_),
    .S(_3351_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6906_ (.A1(_3355_),
    .A2(\registers[10][8] ),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6907_ (.I0(_1108_),
    .I1(_3362_),
    .S(_3325_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6908_ (.A1(_3355_),
    .A2(\registers[10][9] ),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6909_ (.I0(_1110_),
    .I1(_3363_),
    .S(_3325_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6910_ (.A1(_1569_),
    .A2(\registers[11][0] ),
    .Z(_3364_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _6911_ (.A1(_1232_),
    .A2(_1498_),
    .Z(_3365_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6912_ (.I(_3365_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6913_ (.I0(_3364_),
    .I1(_1115_),
    .S(_3366_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6914_ (.A1(_1569_),
    .A2(\registers[11][10] ),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6915_ (.I0(_3367_),
    .I1(_1123_),
    .S(_3366_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6916_ (.A1(_1569_),
    .A2(\registers[11][11] ),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6917_ (.I0(_3368_),
    .I1(_1125_),
    .S(_3366_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6918_ (.A1(_1569_),
    .A2(\registers[11][12] ),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6919_ (.I0(_3369_),
    .I1(_1127_),
    .S(_3366_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6920_ (.I(_1223_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6921_ (.A1(_3370_),
    .A2(\registers[11][13] ),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6922_ (.I0(_3371_),
    .I1(_1129_),
    .S(_3366_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6923_ (.A1(_3370_),
    .A2(\registers[11][14] ),
    .Z(_3372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6924_ (.I0(_3372_),
    .I1(_1131_),
    .S(_3366_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6925_ (.A1(_3370_),
    .A2(\registers[11][15] ),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6926_ (.I0(_3373_),
    .I1(_1133_),
    .S(_3366_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6927_ (.A1(_3370_),
    .A2(\registers[11][16] ),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6928_ (.I0(_3374_),
    .I1(_1135_),
    .S(_3366_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6929_ (.A1(_3370_),
    .A2(\registers[11][17] ),
    .Z(_3375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6930_ (.I0(_3375_),
    .I1(_1137_),
    .S(_3366_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6931_ (.A1(_3370_),
    .A2(\registers[11][18] ),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6932_ (.I0(_3376_),
    .I1(_1139_),
    .S(_3366_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6933_ (.A1(_3370_),
    .A2(\registers[11][19] ),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6934_ (.I(_3365_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6935_ (.I0(_3377_),
    .I1(_1142_),
    .S(_3378_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6936_ (.A1(_3370_),
    .A2(\registers[11][1] ),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6937_ (.I0(_3379_),
    .I1(_1145_),
    .S(_3378_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6938_ (.A1(_3370_),
    .A2(\registers[11][20] ),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6939_ (.I0(_3380_),
    .I1(_1147_),
    .S(_3378_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6940_ (.A1(_3370_),
    .A2(\registers[11][21] ),
    .Z(_3381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6941_ (.I0(_3381_),
    .I1(_1149_),
    .S(_3378_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6942_ (.I(_1223_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6943_ (.A1(_3382_),
    .A2(\registers[11][22] ),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6944_ (.I0(_3383_),
    .I1(_1151_),
    .S(_3378_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6945_ (.A1(_3382_),
    .A2(\registers[11][23] ),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6946_ (.I0(_3384_),
    .I1(_1153_),
    .S(_3378_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6947_ (.A1(_3382_),
    .A2(\registers[11][24] ),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6948_ (.I0(_3385_),
    .I1(_1155_),
    .S(_3378_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6949_ (.A1(_3382_),
    .A2(\registers[11][25] ),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6950_ (.I0(_3386_),
    .I1(_1157_),
    .S(_3378_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6951_ (.A1(_3382_),
    .A2(\registers[11][26] ),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6952_ (.I0(_3387_),
    .I1(_1159_),
    .S(_3378_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6953_ (.A1(_3382_),
    .A2(\registers[11][27] ),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6954_ (.I0(_3388_),
    .I1(_1161_),
    .S(_3378_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6955_ (.A1(_3382_),
    .A2(\registers[11][28] ),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6956_ (.I(_3365_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6957_ (.I0(_3389_),
    .I1(_1164_),
    .S(_3390_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6958_ (.A1(_3382_),
    .A2(\registers[11][29] ),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6959_ (.I0(_3391_),
    .I1(_1167_),
    .S(_3390_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6960_ (.A1(_3382_),
    .A2(\registers[11][2] ),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6961_ (.I0(_3392_),
    .I1(_1169_),
    .S(_3390_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6962_ (.A1(_3382_),
    .A2(\registers[11][30] ),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6963_ (.I0(_3393_),
    .I1(_1171_),
    .S(_3390_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _6964_ (.I(_1223_),
    .Z(_3394_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6965_ (.A1(_3394_),
    .A2(\registers[11][31] ),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6966_ (.I0(_3395_),
    .I1(_1173_),
    .S(_3390_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6967_ (.A1(_3394_),
    .A2(\registers[11][3] ),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6968_ (.I0(_3396_),
    .I1(_1175_),
    .S(_3390_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6969_ (.A1(_3394_),
    .A2(\registers[11][4] ),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6970_ (.I0(_3397_),
    .I1(_1177_),
    .S(_3390_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6971_ (.A1(_3394_),
    .A2(\registers[11][5] ),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6972_ (.I0(_3398_),
    .I1(_1179_),
    .S(_3390_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6973_ (.A1(_3394_),
    .A2(\registers[11][6] ),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6974_ (.I0(_3399_),
    .I1(_1181_),
    .S(_3390_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6975_ (.A1(_3394_),
    .A2(\registers[11][7] ),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6976_ (.I0(_3400_),
    .I1(_1183_),
    .S(_3390_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6977_ (.A1(_3394_),
    .A2(\registers[11][8] ),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6978_ (.I0(_3401_),
    .I1(_1186_),
    .S(_3365_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6979_ (.A1(_3394_),
    .A2(\registers[11][9] ),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6980_ (.I0(_3402_),
    .I1(_1188_),
    .S(_3365_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6981_ (.A1(_3355_),
    .A2(\registers[12][0] ),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _6982_ (.A1(net13),
    .A2(_1497_),
    .A3(net12),
    .Z(_3404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _6983_ (.A1(_1338_),
    .A2(_3404_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _6984_ (.I(_3405_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6985_ (.I0(_1229_),
    .I1(_3403_),
    .S(_3406_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6986_ (.A1(_3355_),
    .A2(\registers[12][10] ),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6987_ (.I0(_1235_),
    .I1(_3407_),
    .S(_3406_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _6988_ (.I(_3330_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6989_ (.A1(_3408_),
    .A2(\registers[12][11] ),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6990_ (.I0(_1237_),
    .I1(_3409_),
    .S(_3406_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6991_ (.A1(_3408_),
    .A2(\registers[12][12] ),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6992_ (.I0(_1239_),
    .I1(_3410_),
    .S(_3406_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6993_ (.A1(_3408_),
    .A2(\registers[12][13] ),
    .Z(_3411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6994_ (.I0(_1241_),
    .I1(_3411_),
    .S(_3406_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6995_ (.A1(_3408_),
    .A2(\registers[12][14] ),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6996_ (.I0(_1243_),
    .I1(_3412_),
    .S(_3406_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6997_ (.A1(_3408_),
    .A2(\registers[12][15] ),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _6998_ (.I0(_1245_),
    .I1(_3413_),
    .S(_3406_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _6999_ (.A1(_3408_),
    .A2(\registers[12][16] ),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7000_ (.I0(_1247_),
    .I1(_3414_),
    .S(_3406_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7001_ (.A1(_3408_),
    .A2(\registers[12][17] ),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7002_ (.I0(_1249_),
    .I1(_3415_),
    .S(_3406_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7003_ (.A1(_3408_),
    .A2(\registers[12][18] ),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7004_ (.I0(_1251_),
    .I1(_3416_),
    .S(_3406_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7005_ (.A1(_3408_),
    .A2(\registers[12][19] ),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7006_ (.I(_3405_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7007_ (.I0(_1253_),
    .I1(_3417_),
    .S(_3418_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7008_ (.A1(_3408_),
    .A2(\registers[12][1] ),
    .Z(_3419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7009_ (.I0(_1257_),
    .I1(_3419_),
    .S(_3418_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7010_ (.I(_3330_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7011_ (.A1(_3420_),
    .A2(\registers[12][20] ),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7012_ (.I0(_1259_),
    .I1(_3421_),
    .S(_3418_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7013_ (.A1(_3420_),
    .A2(\registers[12][21] ),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7014_ (.I0(_1261_),
    .I1(_3422_),
    .S(_3418_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7015_ (.A1(_3420_),
    .A2(\registers[12][22] ),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7016_ (.I0(_1263_),
    .I1(_3423_),
    .S(_3418_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7017_ (.A1(_3420_),
    .A2(\registers[12][23] ),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7018_ (.I0(_1265_),
    .I1(_3424_),
    .S(_3418_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7019_ (.A1(_3420_),
    .A2(\registers[12][24] ),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7020_ (.I0(_1267_),
    .I1(_3425_),
    .S(_3418_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7021_ (.A1(_3420_),
    .A2(\registers[12][25] ),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7022_ (.I0(_1269_),
    .I1(_3426_),
    .S(_3418_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7023_ (.A1(_3420_),
    .A2(\registers[12][26] ),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7024_ (.I0(_1271_),
    .I1(_3427_),
    .S(_3418_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7025_ (.A1(_3420_),
    .A2(\registers[12][27] ),
    .Z(_3428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7026_ (.I0(_1273_),
    .I1(_3428_),
    .S(_3418_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7027_ (.A1(_3420_),
    .A2(\registers[12][28] ),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7028_ (.I(_3405_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7029_ (.I0(_1275_),
    .I1(_3429_),
    .S(_3430_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7030_ (.A1(_3420_),
    .A2(\registers[12][29] ),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7031_ (.I0(_1279_),
    .I1(_3431_),
    .S(_3430_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7032_ (.I(_3330_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7033_ (.A1(_3432_),
    .A2(\registers[12][2] ),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7034_ (.I0(_1281_),
    .I1(_3433_),
    .S(_3430_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7035_ (.A1(_3432_),
    .A2(\registers[12][30] ),
    .Z(_3434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7036_ (.I0(_1283_),
    .I1(_3434_),
    .S(_3430_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7037_ (.I(net39),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7038_ (.A1(_3432_),
    .A2(\registers[12][31] ),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7039_ (.I0(_3435_),
    .I1(_3436_),
    .S(_3430_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _7040_ (.I(net40),
    .Z(_3437_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7041_ (.A1(_3432_),
    .A2(\registers[12][3] ),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7042_ (.I0(_3437_),
    .I1(_3438_),
    .S(_3430_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7043_ (.I(net41),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7044_ (.A1(_3432_),
    .A2(\registers[12][4] ),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7045_ (.I0(_3439_),
    .I1(_3440_),
    .S(_3430_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7046_ (.I(net42),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7047_ (.A1(_3432_),
    .A2(\registers[12][5] ),
    .Z(_3442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7048_ (.I0(_3441_),
    .I1(_3442_),
    .S(_3430_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7049_ (.I(net43),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7050_ (.A1(_3432_),
    .A2(\registers[12][6] ),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7051_ (.I0(_3443_),
    .I1(_3444_),
    .S(_3430_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7052_ (.I(net44),
    .Z(_3445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7053_ (.A1(_3432_),
    .A2(\registers[12][7] ),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7054_ (.I0(_3445_),
    .I1(_3446_),
    .S(_3430_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7055_ (.I(net45),
    .Z(_3447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7056_ (.A1(_3432_),
    .A2(\registers[12][8] ),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7057_ (.I0(_3447_),
    .I1(_3448_),
    .S(_3405_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7058_ (.I(net46),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7059_ (.A1(_3432_),
    .A2(\registers[12][9] ),
    .Z(_3450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7060_ (.I0(_3449_),
    .I1(_3450_),
    .S(_3405_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _7061_ (.I(net15),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7062_ (.I(_3330_),
    .Z(_3452_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7063_ (.A1(_3452_),
    .A2(\registers[13][0] ),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7064_ (.A1(_1095_),
    .A2(_3404_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7065_ (.I(_3454_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7066_ (.I0(_3451_),
    .I1(_3453_),
    .S(_3455_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7067_ (.I(net16),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7068_ (.A1(_3452_),
    .A2(\registers[13][10] ),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7069_ (.I0(_3456_),
    .I1(_3457_),
    .S(_3455_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _7070_ (.I(net17),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7071_ (.A1(_3452_),
    .A2(\registers[13][11] ),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7072_ (.I0(_3458_),
    .I1(_3459_),
    .S(_3455_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7073_ (.I(net18),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7074_ (.A1(_3452_),
    .A2(\registers[13][12] ),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7075_ (.I0(_3460_),
    .I1(_3461_),
    .S(_3455_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7076_ (.I(net19),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7077_ (.A1(_3452_),
    .A2(\registers[13][13] ),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7078_ (.I0(_3462_),
    .I1(_3463_),
    .S(_3455_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7079_ (.I(net20),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7080_ (.A1(_3452_),
    .A2(\registers[13][14] ),
    .Z(_3465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7081_ (.I0(_3464_),
    .I1(_3465_),
    .S(_3455_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7082_ (.I(net21),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7083_ (.A1(_3452_),
    .A2(\registers[13][15] ),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7084_ (.I0(_3466_),
    .I1(_3467_),
    .S(_3455_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7085_ (.I(net22),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7086_ (.A1(_3452_),
    .A2(\registers[13][16] ),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7087_ (.I0(_3468_),
    .I1(_3469_),
    .S(_3455_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7088_ (.I(net23),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7089_ (.A1(_3452_),
    .A2(\registers[13][17] ),
    .Z(_3471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7090_ (.I0(_3470_),
    .I1(_3471_),
    .S(_3455_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7091_ (.I(net24),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7092_ (.A1(_3452_),
    .A2(\registers[13][18] ),
    .Z(_3473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7093_ (.I0(_3472_),
    .I1(_3473_),
    .S(_3455_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7094_ (.I(net25),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7095_ (.I(_3330_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7096_ (.A1(_3475_),
    .A2(\registers[13][19] ),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7097_ (.I(_3454_),
    .Z(_3477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7098_ (.I0(_3474_),
    .I1(_3476_),
    .S(_3477_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7099_ (.I(net26),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7100_ (.A1(_3475_),
    .A2(\registers[13][1] ),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7101_ (.I0(_3478_),
    .I1(_3479_),
    .S(_3477_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _7102_ (.I(net27),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7103_ (.A1(_3475_),
    .A2(\registers[13][20] ),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7104_ (.I0(_3480_),
    .I1(_3481_),
    .S(_3477_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _7105_ (.I(net28),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7106_ (.A1(_3475_),
    .A2(\registers[13][21] ),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7107_ (.I0(_3482_),
    .I1(_3483_),
    .S(_3477_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7108_ (.I(net29),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7109_ (.A1(_3475_),
    .A2(\registers[13][22] ),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7110_ (.I0(_3484_),
    .I1(_3485_),
    .S(_3477_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7111_ (.I(net30),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7112_ (.A1(_3475_),
    .A2(\registers[13][23] ),
    .Z(_3487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7113_ (.I0(_3486_),
    .I1(_3487_),
    .S(_3477_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7114_ (.I(net31),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7115_ (.A1(_3475_),
    .A2(\registers[13][24] ),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7116_ (.I0(_3488_),
    .I1(_3489_),
    .S(_3477_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7117_ (.I(net32),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7118_ (.A1(_3475_),
    .A2(\registers[13][25] ),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7119_ (.I0(_3490_),
    .I1(_3491_),
    .S(_3477_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7120_ (.I(net33),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7121_ (.A1(_3475_),
    .A2(\registers[13][26] ),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7122_ (.I0(_3492_),
    .I1(_3493_),
    .S(_3477_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _7123_ (.I(net34),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7124_ (.A1(_3475_),
    .A2(\registers[13][27] ),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7125_ (.I0(_3494_),
    .I1(_3495_),
    .S(_3477_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7126_ (.I(net35),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7127_ (.I(_3330_),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7128_ (.A1(_3497_),
    .A2(\registers[13][28] ),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7129_ (.I(_3454_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7130_ (.I0(_3496_),
    .I1(_3498_),
    .S(_3499_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7131_ (.I(net36),
    .Z(_3500_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7132_ (.A1(_3497_),
    .A2(\registers[13][29] ),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7133_ (.I0(_3500_),
    .I1(_3501_),
    .S(_3499_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7134_ (.I(net37),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7135_ (.A1(_3497_),
    .A2(\registers[13][2] ),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7136_ (.I0(_3502_),
    .I1(_3503_),
    .S(_3499_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7137_ (.I(net38),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7138_ (.A1(_3497_),
    .A2(\registers[13][30] ),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7139_ (.I0(_3504_),
    .I1(_3505_),
    .S(_3499_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7140_ (.A1(_3497_),
    .A2(\registers[13][31] ),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7141_ (.I0(_3435_),
    .I1(_3506_),
    .S(_3499_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7142_ (.A1(_3497_),
    .A2(\registers[13][3] ),
    .Z(_3507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7143_ (.I0(_3437_),
    .I1(_3507_),
    .S(_3499_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7144_ (.A1(_3497_),
    .A2(\registers[13][4] ),
    .Z(_3508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7145_ (.I0(_3439_),
    .I1(_3508_),
    .S(_3499_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7146_ (.A1(_3497_),
    .A2(\registers[13][5] ),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7147_ (.I0(_3441_),
    .I1(_3509_),
    .S(_3499_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7148_ (.A1(_3497_),
    .A2(\registers[13][6] ),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7149_ (.I0(_3443_),
    .I1(_3510_),
    .S(_3499_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7150_ (.A1(_3497_),
    .A2(\registers[13][7] ),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7151_ (.I0(_3445_),
    .I1(_3511_),
    .S(_3499_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7152_ (.I(_3330_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7153_ (.A1(_3512_),
    .A2(\registers[13][8] ),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7154_ (.I0(_3447_),
    .I1(_3513_),
    .S(_3454_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7155_ (.A1(_3512_),
    .A2(\registers[13][9] ),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7156_ (.I0(_3449_),
    .I1(_3514_),
    .S(_3454_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7157_ (.A1(_3512_),
    .A2(\registers[14][0] ),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7158_ (.A1(_1119_),
    .A2(_3404_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7159_ (.I(_3516_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7160_ (.I0(_3451_),
    .I1(_3515_),
    .S(_3517_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7161_ (.A1(_3512_),
    .A2(\registers[14][10] ),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7162_ (.I0(_3456_),
    .I1(_3518_),
    .S(_3517_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7163_ (.A1(_3512_),
    .A2(\registers[14][11] ),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7164_ (.I0(_3458_),
    .I1(_3519_),
    .S(_3517_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7165_ (.A1(_3512_),
    .A2(\registers[14][12] ),
    .Z(_3520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7166_ (.I0(_3460_),
    .I1(_3520_),
    .S(_3517_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7167_ (.A1(_3512_),
    .A2(\registers[14][13] ),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7168_ (.I0(_3462_),
    .I1(_3521_),
    .S(_3517_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7169_ (.A1(_3512_),
    .A2(\registers[14][14] ),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7170_ (.I0(_3464_),
    .I1(_3522_),
    .S(_3517_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7171_ (.A1(_3512_),
    .A2(\registers[14][15] ),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7172_ (.I0(_3466_),
    .I1(_3523_),
    .S(_3517_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7173_ (.A1(_3512_),
    .A2(\registers[14][16] ),
    .Z(_3524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7174_ (.I0(_3468_),
    .I1(_3524_),
    .S(_3517_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7175_ (.I(_1089_),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7176_ (.I(_3525_),
    .Z(_3526_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7177_ (.A1(_3526_),
    .A2(\registers[14][17] ),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7178_ (.I0(_3470_),
    .I1(_3527_),
    .S(_3517_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7179_ (.A1(_3526_),
    .A2(\registers[14][18] ),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7180_ (.I0(_3472_),
    .I1(_3528_),
    .S(_3517_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7181_ (.A1(_3526_),
    .A2(\registers[14][19] ),
    .Z(_3529_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7182_ (.I(_3516_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7183_ (.I0(_3474_),
    .I1(_3529_),
    .S(_3530_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7184_ (.A1(_3526_),
    .A2(\registers[14][1] ),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7185_ (.I0(_3478_),
    .I1(_3531_),
    .S(_3530_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7186_ (.A1(_3526_),
    .A2(\registers[14][20] ),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7187_ (.I0(_3480_),
    .I1(_3532_),
    .S(_3530_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7188_ (.A1(_3526_),
    .A2(\registers[14][21] ),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7189_ (.I0(_3482_),
    .I1(_3533_),
    .S(_3530_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7190_ (.A1(_3526_),
    .A2(\registers[14][22] ),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7191_ (.I0(_3484_),
    .I1(_3534_),
    .S(_3530_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7192_ (.A1(_3526_),
    .A2(\registers[14][23] ),
    .Z(_3535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7193_ (.I0(_3486_),
    .I1(_3535_),
    .S(_3530_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7194_ (.A1(_3526_),
    .A2(\registers[14][24] ),
    .Z(_3536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7195_ (.I0(_3488_),
    .I1(_3536_),
    .S(_3530_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7196_ (.A1(_3526_),
    .A2(\registers[14][25] ),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7197_ (.I0(_3490_),
    .I1(_3537_),
    .S(_3530_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7198_ (.I(_3525_),
    .Z(_3538_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7199_ (.A1(_3538_),
    .A2(\registers[14][26] ),
    .Z(_3539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7200_ (.I0(_3492_),
    .I1(_3539_),
    .S(_3530_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7201_ (.A1(_3538_),
    .A2(\registers[14][27] ),
    .Z(_3540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7202_ (.I0(_3494_),
    .I1(_3540_),
    .S(_3530_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7203_ (.A1(_3538_),
    .A2(\registers[14][28] ),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7204_ (.I(_3516_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7205_ (.I0(_3496_),
    .I1(_3541_),
    .S(_3542_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7206_ (.A1(_3538_),
    .A2(\registers[14][29] ),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7207_ (.I0(_3500_),
    .I1(_3543_),
    .S(_3542_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7208_ (.A1(_3538_),
    .A2(\registers[14][2] ),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7209_ (.I0(_3502_),
    .I1(_3544_),
    .S(_3542_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7210_ (.A1(_3538_),
    .A2(\registers[14][30] ),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7211_ (.I0(_3504_),
    .I1(_3545_),
    .S(_3542_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7212_ (.A1(_3538_),
    .A2(\registers[14][31] ),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7213_ (.I0(_3435_),
    .I1(_3546_),
    .S(_3542_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7214_ (.A1(_3538_),
    .A2(\registers[14][3] ),
    .Z(_3547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7215_ (.I0(_3437_),
    .I1(_3547_),
    .S(_3542_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7216_ (.A1(_3538_),
    .A2(\registers[14][4] ),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7217_ (.I0(_3439_),
    .I1(_3548_),
    .S(_3542_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7218_ (.A1(_3538_),
    .A2(\registers[14][5] ),
    .Z(_3549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7219_ (.I0(_3441_),
    .I1(_3549_),
    .S(_3542_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7220_ (.I(_3525_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7221_ (.A1(_3550_),
    .A2(\registers[14][6] ),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7222_ (.I0(_3443_),
    .I1(_3551_),
    .S(_3542_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7223_ (.A1(_3550_),
    .A2(\registers[14][7] ),
    .Z(_3552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7224_ (.I0(_3445_),
    .I1(_3552_),
    .S(_3542_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7225_ (.A1(_3550_),
    .A2(\registers[14][8] ),
    .Z(_3553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7226_ (.I0(_3447_),
    .I1(_3553_),
    .S(_3516_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7227_ (.A1(_3550_),
    .A2(\registers[14][9] ),
    .Z(_3554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7228_ (.I0(_3449_),
    .I1(_3554_),
    .S(_3516_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7229_ (.A1(_3550_),
    .A2(\registers[15][0] ),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7230_ (.A1(_1232_),
    .A2(_3404_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7231_ (.I(_3556_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7232_ (.I0(_3451_),
    .I1(_3555_),
    .S(_3557_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7233_ (.A1(_3550_),
    .A2(\registers[15][10] ),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7234_ (.I0(_3456_),
    .I1(_3558_),
    .S(_3557_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7235_ (.A1(_3550_),
    .A2(\registers[15][11] ),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7236_ (.I0(_3458_),
    .I1(_3559_),
    .S(_3557_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7237_ (.A1(_3550_),
    .A2(\registers[15][12] ),
    .Z(_3560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7238_ (.I0(_3460_),
    .I1(_3560_),
    .S(_3557_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7239_ (.A1(_3550_),
    .A2(\registers[15][13] ),
    .Z(_3561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7240_ (.I0(_3462_),
    .I1(_3561_),
    .S(_3557_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7241_ (.A1(_3550_),
    .A2(\registers[15][14] ),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7242_ (.I0(_3464_),
    .I1(_3562_),
    .S(_3557_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7243_ (.I(_3525_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7244_ (.A1(_3563_),
    .A2(\registers[15][15] ),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7245_ (.I0(_3466_),
    .I1(_3564_),
    .S(_3557_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7246_ (.A1(_3563_),
    .A2(\registers[15][16] ),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7247_ (.I0(_3468_),
    .I1(_3565_),
    .S(_3557_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7248_ (.A1(_3563_),
    .A2(\registers[15][17] ),
    .Z(_3566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7249_ (.I0(_3470_),
    .I1(_3566_),
    .S(_3557_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7250_ (.A1(_3563_),
    .A2(\registers[15][18] ),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7251_ (.I0(_3472_),
    .I1(_3567_),
    .S(_3557_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7252_ (.A1(_3563_),
    .A2(\registers[15][19] ),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7253_ (.I(_3556_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7254_ (.I0(_3474_),
    .I1(_3568_),
    .S(_3569_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7255_ (.A1(_3563_),
    .A2(\registers[15][1] ),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7256_ (.I0(_3478_),
    .I1(_3570_),
    .S(_3569_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7257_ (.A1(_3563_),
    .A2(\registers[15][20] ),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7258_ (.I0(_3480_),
    .I1(_3571_),
    .S(_3569_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7259_ (.A1(_3563_),
    .A2(\registers[15][21] ),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7260_ (.I0(_3482_),
    .I1(_3572_),
    .S(_3569_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7261_ (.A1(_3563_),
    .A2(\registers[15][22] ),
    .Z(_3573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7262_ (.I0(_3484_),
    .I1(_3573_),
    .S(_3569_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7263_ (.A1(_3563_),
    .A2(\registers[15][23] ),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7264_ (.I0(_3486_),
    .I1(_3574_),
    .S(_3569_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7265_ (.I(_3525_),
    .Z(_3575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7266_ (.A1(_3575_),
    .A2(\registers[15][24] ),
    .Z(_3576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7267_ (.I0(_3488_),
    .I1(_3576_),
    .S(_3569_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7268_ (.A1(_3575_),
    .A2(\registers[15][25] ),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7269_ (.I0(_3490_),
    .I1(_3577_),
    .S(_3569_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7270_ (.A1(_3575_),
    .A2(\registers[15][26] ),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7271_ (.I0(_3492_),
    .I1(_3578_),
    .S(_3569_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7272_ (.A1(_3575_),
    .A2(\registers[15][27] ),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7273_ (.I0(_3494_),
    .I1(_3579_),
    .S(_3569_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7274_ (.A1(_3575_),
    .A2(\registers[15][28] ),
    .Z(_3580_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7275_ (.I(_3556_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7276_ (.I0(_3496_),
    .I1(_3580_),
    .S(_3581_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7277_ (.A1(_3575_),
    .A2(\registers[15][29] ),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7278_ (.I0(_3500_),
    .I1(_3582_),
    .S(_3581_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7279_ (.A1(_3575_),
    .A2(\registers[15][2] ),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7280_ (.I0(_3502_),
    .I1(_3583_),
    .S(_3581_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7281_ (.A1(_3575_),
    .A2(\registers[15][30] ),
    .Z(_3584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7282_ (.I0(_3504_),
    .I1(_3584_),
    .S(_3581_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7283_ (.A1(_3575_),
    .A2(\registers[15][31] ),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7284_ (.I0(_3435_),
    .I1(_3585_),
    .S(_3581_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7285_ (.A1(_3575_),
    .A2(\registers[15][3] ),
    .Z(_3586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7286_ (.I0(_3437_),
    .I1(_3586_),
    .S(_3581_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7287_ (.I(_3525_),
    .Z(_3587_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7288_ (.A1(_3587_),
    .A2(\registers[15][4] ),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7289_ (.I0(_3439_),
    .I1(_3588_),
    .S(_3581_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7290_ (.A1(_3587_),
    .A2(\registers[15][5] ),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7291_ (.I0(_3441_),
    .I1(_3589_),
    .S(_3581_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7292_ (.A1(_3587_),
    .A2(\registers[15][6] ),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7293_ (.I0(_3443_),
    .I1(_3590_),
    .S(_3581_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7294_ (.A1(_3587_),
    .A2(\registers[15][7] ),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7295_ (.I0(_3445_),
    .I1(_3591_),
    .S(_3581_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7296_ (.A1(_3587_),
    .A2(\registers[15][8] ),
    .Z(_3592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7297_ (.I0(_3447_),
    .I1(_3592_),
    .S(_3556_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7298_ (.A1(_3587_),
    .A2(\registers[15][9] ),
    .Z(_3593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7299_ (.I0(_3449_),
    .I1(_3593_),
    .S(_3556_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7300_ (.A1(_3587_),
    .A2(\registers[16][0] ),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _7301_ (.A1(net13),
    .A2(_1497_),
    .A3(net12),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _7302_ (.A1(net10),
    .A2(net11),
    .A3(_1117_),
    .A4(_3595_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7303_ (.I(_3596_),
    .Z(_3597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7304_ (.I0(_3451_),
    .I1(_3594_),
    .S(_3597_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7305_ (.A1(_3587_),
    .A2(\registers[16][10] ),
    .Z(_3598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7306_ (.I0(_3456_),
    .I1(_3598_),
    .S(_3597_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7307_ (.A1(_3587_),
    .A2(\registers[16][11] ),
    .Z(_3599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7308_ (.I0(_3458_),
    .I1(_3599_),
    .S(_3597_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7309_ (.A1(_3587_),
    .A2(\registers[16][12] ),
    .Z(_3600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7310_ (.I0(_3460_),
    .I1(_3600_),
    .S(_3597_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7311_ (.I(_3525_),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7312_ (.A1(_3601_),
    .A2(\registers[16][13] ),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7313_ (.I0(_3462_),
    .I1(_3602_),
    .S(_3597_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7314_ (.A1(_3601_),
    .A2(\registers[16][14] ),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7315_ (.I0(_3464_),
    .I1(_3603_),
    .S(_3597_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7316_ (.A1(_3601_),
    .A2(\registers[16][15] ),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7317_ (.I0(_3466_),
    .I1(_3604_),
    .S(_3597_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7318_ (.A1(_3601_),
    .A2(\registers[16][16] ),
    .Z(_3605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7319_ (.I0(_3468_),
    .I1(_3605_),
    .S(_3597_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7320_ (.A1(_3601_),
    .A2(\registers[16][17] ),
    .Z(_3606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7321_ (.I0(_3470_),
    .I1(_3606_),
    .S(_3597_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7322_ (.A1(_3601_),
    .A2(\registers[16][18] ),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7323_ (.I0(_3472_),
    .I1(_3607_),
    .S(_3597_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7324_ (.A1(_3601_),
    .A2(\registers[16][19] ),
    .Z(_3608_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7325_ (.I(_3596_),
    .Z(_3609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7326_ (.I0(_3474_),
    .I1(_3608_),
    .S(_3609_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7327_ (.A1(_3601_),
    .A2(\registers[16][1] ),
    .Z(_3610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7328_ (.I0(_3478_),
    .I1(_3610_),
    .S(_3609_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7329_ (.A1(_3601_),
    .A2(\registers[16][20] ),
    .Z(_3611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7330_ (.I0(_3480_),
    .I1(_3611_),
    .S(_3609_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7331_ (.A1(_3601_),
    .A2(\registers[16][21] ),
    .Z(_3612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7332_ (.I0(_3482_),
    .I1(_3612_),
    .S(_3609_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7333_ (.I(_3525_),
    .Z(_3613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7334_ (.A1(_3613_),
    .A2(\registers[16][22] ),
    .Z(_3614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7335_ (.I0(_3484_),
    .I1(_3614_),
    .S(_3609_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7336_ (.A1(_3613_),
    .A2(\registers[16][23] ),
    .Z(_3615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7337_ (.I0(_3486_),
    .I1(_3615_),
    .S(_3609_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7338_ (.A1(_3613_),
    .A2(\registers[16][24] ),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7339_ (.I0(_3488_),
    .I1(_3616_),
    .S(_3609_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7340_ (.A1(_3613_),
    .A2(\registers[16][25] ),
    .Z(_3617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7341_ (.I0(_3490_),
    .I1(_3617_),
    .S(_3609_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7342_ (.A1(_3613_),
    .A2(\registers[16][26] ),
    .Z(_3618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7343_ (.I0(_3492_),
    .I1(_3618_),
    .S(_3609_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7344_ (.A1(_3613_),
    .A2(\registers[16][27] ),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7345_ (.I0(_3494_),
    .I1(_3619_),
    .S(_3609_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7346_ (.A1(_3613_),
    .A2(\registers[16][28] ),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7347_ (.I(_3596_),
    .Z(_3621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7348_ (.I0(_3496_),
    .I1(_3620_),
    .S(_3621_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7349_ (.A1(_3613_),
    .A2(\registers[16][29] ),
    .Z(_3622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7350_ (.I0(_3500_),
    .I1(_3622_),
    .S(_3621_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7351_ (.A1(_3613_),
    .A2(\registers[16][2] ),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7352_ (.I0(_3502_),
    .I1(_3623_),
    .S(_3621_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7353_ (.A1(_3613_),
    .A2(\registers[16][30] ),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7354_ (.I0(_3504_),
    .I1(_3624_),
    .S(_3621_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7355_ (.I(_3525_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7356_ (.A1(_3625_),
    .A2(\registers[16][31] ),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7357_ (.I0(_3435_),
    .I1(_3626_),
    .S(_3621_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7358_ (.A1(_3625_),
    .A2(\registers[16][3] ),
    .Z(_3627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7359_ (.I0(_3437_),
    .I1(_3627_),
    .S(_3621_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7360_ (.A1(_3625_),
    .A2(\registers[16][4] ),
    .Z(_3628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7361_ (.I0(_3439_),
    .I1(_3628_),
    .S(_3621_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7362_ (.A1(_3625_),
    .A2(\registers[16][5] ),
    .Z(_3629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7363_ (.I0(_3441_),
    .I1(_3629_),
    .S(_3621_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7364_ (.A1(_3625_),
    .A2(\registers[16][6] ),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7365_ (.I0(_3443_),
    .I1(_3630_),
    .S(_3621_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7366_ (.A1(_3625_),
    .A2(\registers[16][7] ),
    .Z(_3631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7367_ (.I0(_3445_),
    .I1(_3631_),
    .S(_3621_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7368_ (.A1(_3625_),
    .A2(\registers[16][8] ),
    .Z(_3632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7369_ (.I0(_3447_),
    .I1(_3632_),
    .S(_3596_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7370_ (.A1(_3625_),
    .A2(\registers[16][9] ),
    .Z(_3633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7371_ (.I0(_3449_),
    .I1(_3633_),
    .S(_3596_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7372_ (.A1(_3625_),
    .A2(\registers[17][0] ),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _7373_ (.A1(net11),
    .A2(_1094_),
    .A3(_3595_),
    .Z(_3635_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7374_ (.I(_3635_),
    .Z(_3636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7375_ (.I0(_3451_),
    .I1(_3634_),
    .S(_3636_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7376_ (.A1(_3625_),
    .A2(\registers[17][10] ),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7377_ (.I0(_3456_),
    .I1(_3637_),
    .S(_3636_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7378_ (.I(_3525_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7379_ (.A1(_3638_),
    .A2(\registers[17][11] ),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7380_ (.I0(_3458_),
    .I1(_3639_),
    .S(_3636_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7381_ (.A1(_3638_),
    .A2(\registers[17][12] ),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7382_ (.I0(_3460_),
    .I1(_3640_),
    .S(_3636_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7383_ (.A1(_3638_),
    .A2(\registers[17][13] ),
    .Z(_3641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7384_ (.I0(_3462_),
    .I1(_3641_),
    .S(_3636_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7385_ (.A1(_3638_),
    .A2(\registers[17][14] ),
    .Z(_3642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7386_ (.I0(_3464_),
    .I1(_3642_),
    .S(_3636_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7387_ (.A1(_3638_),
    .A2(\registers[17][15] ),
    .Z(_3643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7388_ (.I0(_3466_),
    .I1(_3643_),
    .S(_3636_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7389_ (.A1(_3638_),
    .A2(\registers[17][16] ),
    .Z(_3644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7390_ (.I0(_3468_),
    .I1(_3644_),
    .S(_3636_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7391_ (.A1(_3638_),
    .A2(\registers[17][17] ),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7392_ (.I0(_3470_),
    .I1(_3645_),
    .S(_3636_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7393_ (.A1(_3638_),
    .A2(\registers[17][18] ),
    .Z(_3646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7394_ (.I0(_3472_),
    .I1(_3646_),
    .S(_3636_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7395_ (.A1(_3638_),
    .A2(\registers[17][19] ),
    .Z(_3647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7396_ (.I(_3635_),
    .Z(_3648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7397_ (.I0(_3474_),
    .I1(_3647_),
    .S(_3648_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7398_ (.A1(_3638_),
    .A2(\registers[17][1] ),
    .Z(_3649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7399_ (.I0(_3478_),
    .I1(_3649_),
    .S(_3648_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7400_ (.I(_1089_),
    .Z(_3650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7401_ (.I(_3650_),
    .Z(_3651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7402_ (.A1(_3651_),
    .A2(\registers[17][20] ),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7403_ (.I0(_3480_),
    .I1(_3652_),
    .S(_3648_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7404_ (.A1(_3651_),
    .A2(\registers[17][21] ),
    .Z(_3653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7405_ (.I0(_3482_),
    .I1(_3653_),
    .S(_3648_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7406_ (.A1(_3651_),
    .A2(\registers[17][22] ),
    .Z(_3654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7407_ (.I0(_3484_),
    .I1(_3654_),
    .S(_3648_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7408_ (.A1(_3651_),
    .A2(\registers[17][23] ),
    .Z(_3655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7409_ (.I0(_3486_),
    .I1(_3655_),
    .S(_3648_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7410_ (.A1(_3651_),
    .A2(\registers[17][24] ),
    .Z(_3656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7411_ (.I0(_3488_),
    .I1(_3656_),
    .S(_3648_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7412_ (.A1(_3651_),
    .A2(\registers[17][25] ),
    .Z(_3657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7413_ (.I0(_3490_),
    .I1(_3657_),
    .S(_3648_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7414_ (.A1(_3651_),
    .A2(\registers[17][26] ),
    .Z(_3658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7415_ (.I0(_3492_),
    .I1(_3658_),
    .S(_3648_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7416_ (.A1(_3651_),
    .A2(\registers[17][27] ),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7417_ (.I0(_3494_),
    .I1(_3659_),
    .S(_3648_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7418_ (.A1(_3651_),
    .A2(\registers[17][28] ),
    .Z(_3660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7419_ (.I(_3635_),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7420_ (.I0(_3496_),
    .I1(_3660_),
    .S(_3661_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7421_ (.A1(_3651_),
    .A2(\registers[17][29] ),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7422_ (.I0(_3500_),
    .I1(_3662_),
    .S(_3661_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7423_ (.I(_3650_),
    .Z(_3663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7424_ (.A1(_3663_),
    .A2(\registers[17][2] ),
    .Z(_3664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7425_ (.I0(_3502_),
    .I1(_3664_),
    .S(_3661_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7426_ (.A1(_3663_),
    .A2(\registers[17][30] ),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7427_ (.I0(_3504_),
    .I1(_3665_),
    .S(_3661_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7428_ (.A1(_3663_),
    .A2(\registers[17][31] ),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7429_ (.I0(_3435_),
    .I1(_3666_),
    .S(_3661_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7430_ (.A1(_3663_),
    .A2(\registers[17][3] ),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7431_ (.I0(_3437_),
    .I1(_3667_),
    .S(_3661_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7432_ (.A1(_3663_),
    .A2(\registers[17][4] ),
    .Z(_3668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7433_ (.I0(_3439_),
    .I1(_3668_),
    .S(_3661_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7434_ (.A1(_3663_),
    .A2(\registers[17][5] ),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7435_ (.I0(_3441_),
    .I1(_3669_),
    .S(_3661_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7436_ (.A1(_3663_),
    .A2(\registers[17][6] ),
    .Z(_3670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7437_ (.I0(_3443_),
    .I1(_3670_),
    .S(_3661_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7438_ (.A1(_3663_),
    .A2(\registers[17][7] ),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7439_ (.I0(_3445_),
    .I1(_3671_),
    .S(_3661_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7440_ (.A1(_3663_),
    .A2(\registers[17][8] ),
    .Z(_3672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7441_ (.I0(_3447_),
    .I1(_3672_),
    .S(_3635_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7442_ (.A1(_3663_),
    .A2(\registers[17][9] ),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7443_ (.I0(_3449_),
    .I1(_3673_),
    .S(_3635_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7444_ (.I(_3650_),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7445_ (.A1(_3674_),
    .A2(\registers[18][0] ),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _7446_ (.A1(net11),
    .A2(_1118_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _7447_ (.A1(_3676_),
    .A2(_3595_),
    .Z(_3677_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7448_ (.I(_3677_),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7449_ (.I0(_3451_),
    .I1(_3675_),
    .S(_3678_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7450_ (.A1(_3674_),
    .A2(\registers[18][10] ),
    .Z(_3679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7451_ (.I0(_3456_),
    .I1(_3679_),
    .S(_3678_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7452_ (.A1(_3674_),
    .A2(\registers[18][11] ),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7453_ (.I0(_3458_),
    .I1(_3680_),
    .S(_3678_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7454_ (.A1(_3674_),
    .A2(\registers[18][12] ),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7455_ (.I0(_3460_),
    .I1(_3681_),
    .S(_3678_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7456_ (.A1(_3674_),
    .A2(\registers[18][13] ),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7457_ (.I0(_3462_),
    .I1(_3682_),
    .S(_3678_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7458_ (.A1(_3674_),
    .A2(\registers[18][14] ),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7459_ (.I0(_3464_),
    .I1(_3683_),
    .S(_3678_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7460_ (.A1(_3674_),
    .A2(\registers[18][15] ),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7461_ (.I0(_3466_),
    .I1(_3684_),
    .S(_3678_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7462_ (.A1(_3674_),
    .A2(\registers[18][16] ),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7463_ (.I0(_3468_),
    .I1(_3685_),
    .S(_3678_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7464_ (.A1(_3674_),
    .A2(\registers[18][17] ),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7465_ (.I0(_3470_),
    .I1(_3686_),
    .S(_3678_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7466_ (.A1(_3674_),
    .A2(\registers[18][18] ),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7467_ (.I0(_3472_),
    .I1(_3687_),
    .S(_3678_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7468_ (.I(_3650_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7469_ (.A1(_3688_),
    .A2(\registers[18][19] ),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7470_ (.I(_3677_),
    .Z(_3690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7471_ (.I0(_3474_),
    .I1(_3689_),
    .S(_3690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7472_ (.A1(_3688_),
    .A2(\registers[18][1] ),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7473_ (.I0(_3478_),
    .I1(_3691_),
    .S(_3690_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7474_ (.A1(_3688_),
    .A2(\registers[18][20] ),
    .Z(_3692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7475_ (.I0(_3480_),
    .I1(_3692_),
    .S(_3690_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7476_ (.A1(_3688_),
    .A2(\registers[18][21] ),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7477_ (.I0(_3482_),
    .I1(_3693_),
    .S(_3690_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7478_ (.A1(_3688_),
    .A2(\registers[18][22] ),
    .Z(_3694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7479_ (.I0(_3484_),
    .I1(_3694_),
    .S(_3690_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7480_ (.A1(_3688_),
    .A2(\registers[18][23] ),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7481_ (.I0(_3486_),
    .I1(_3695_),
    .S(_3690_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7482_ (.A1(_3688_),
    .A2(\registers[18][24] ),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7483_ (.I0(_3488_),
    .I1(_3696_),
    .S(_3690_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7484_ (.A1(_3688_),
    .A2(\registers[18][25] ),
    .Z(_3697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7485_ (.I0(_3490_),
    .I1(_3697_),
    .S(_3690_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7486_ (.A1(_3688_),
    .A2(\registers[18][26] ),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7487_ (.I0(_3492_),
    .I1(_3698_),
    .S(_3690_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7488_ (.A1(_3688_),
    .A2(\registers[18][27] ),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7489_ (.I0(_3494_),
    .I1(_3699_),
    .S(_3690_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7490_ (.I(_3650_),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7491_ (.A1(_3700_),
    .A2(\registers[18][28] ),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7492_ (.I(_3677_),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7493_ (.I0(_3496_),
    .I1(_3701_),
    .S(_3702_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7494_ (.A1(_3700_),
    .A2(\registers[18][29] ),
    .Z(_3703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7495_ (.I0(_3500_),
    .I1(_3703_),
    .S(_3702_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7496_ (.A1(_3700_),
    .A2(\registers[18][2] ),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7497_ (.I0(_3502_),
    .I1(_3704_),
    .S(_3702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7498_ (.A1(_3700_),
    .A2(\registers[18][30] ),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7499_ (.I0(_3504_),
    .I1(_3705_),
    .S(_3702_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7500_ (.A1(_3700_),
    .A2(\registers[18][31] ),
    .Z(_3706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7501_ (.I0(_3435_),
    .I1(_3706_),
    .S(_3702_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7502_ (.A1(_3700_),
    .A2(\registers[18][3] ),
    .Z(_3707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7503_ (.I0(_3437_),
    .I1(_3707_),
    .S(_3702_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7504_ (.A1(_3700_),
    .A2(\registers[18][4] ),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7505_ (.I0(_3439_),
    .I1(_3708_),
    .S(_3702_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7506_ (.A1(_3700_),
    .A2(\registers[18][5] ),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7507_ (.I0(_3441_),
    .I1(_3709_),
    .S(_3702_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7508_ (.A1(_3700_),
    .A2(\registers[18][6] ),
    .Z(_3710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7509_ (.I0(_3443_),
    .I1(_3710_),
    .S(_3702_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7510_ (.A1(_3700_),
    .A2(\registers[18][7] ),
    .Z(_3711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7511_ (.I0(_3445_),
    .I1(_3711_),
    .S(_3702_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7512_ (.I(_3650_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7513_ (.A1(_3712_),
    .A2(\registers[18][8] ),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7514_ (.I0(_3447_),
    .I1(_3713_),
    .S(_3677_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7515_ (.A1(_3712_),
    .A2(\registers[18][9] ),
    .Z(_3714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7516_ (.I0(_3449_),
    .I1(_3714_),
    .S(_3677_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7517_ (.A1(_3712_),
    .A2(\registers[19][0] ),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _7518_ (.I(_1232_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _7519_ (.A1(_3716_),
    .A2(_3595_),
    .Z(_3717_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7520_ (.I(_3717_),
    .Z(_3718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7521_ (.I0(_3451_),
    .I1(_3715_),
    .S(_3718_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7522_ (.A1(_3712_),
    .A2(\registers[19][10] ),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7523_ (.I0(_3456_),
    .I1(_3719_),
    .S(_3718_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7524_ (.A1(_3712_),
    .A2(\registers[19][11] ),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7525_ (.I0(_3458_),
    .I1(_3720_),
    .S(_3718_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7526_ (.A1(_3712_),
    .A2(\registers[19][12] ),
    .Z(_3721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7527_ (.I0(_3460_),
    .I1(_3721_),
    .S(_3718_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7528_ (.A1(_3712_),
    .A2(\registers[19][13] ),
    .Z(_3722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7529_ (.I0(_3462_),
    .I1(_3722_),
    .S(_3718_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7530_ (.A1(_3712_),
    .A2(\registers[19][14] ),
    .Z(_3723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7531_ (.I0(_3464_),
    .I1(_3723_),
    .S(_3718_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7532_ (.A1(_3712_),
    .A2(\registers[19][15] ),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7533_ (.I0(_3466_),
    .I1(_3724_),
    .S(_3718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7534_ (.A1(_3712_),
    .A2(\registers[19][16] ),
    .Z(_3725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7535_ (.I0(_3468_),
    .I1(_3725_),
    .S(_3718_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7536_ (.I(_3650_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7537_ (.A1(_3726_),
    .A2(\registers[19][17] ),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7538_ (.I0(_3470_),
    .I1(_3727_),
    .S(_3718_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7539_ (.A1(_3726_),
    .A2(\registers[19][18] ),
    .Z(_3728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7540_ (.I0(_3472_),
    .I1(_3728_),
    .S(_3718_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7541_ (.A1(_3726_),
    .A2(\registers[19][19] ),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7542_ (.I(_3717_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7543_ (.I0(_3474_),
    .I1(_3729_),
    .S(_3730_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7544_ (.A1(_3726_),
    .A2(\registers[19][1] ),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7545_ (.I0(_3478_),
    .I1(_3731_),
    .S(_3730_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7546_ (.A1(_3726_),
    .A2(\registers[19][20] ),
    .Z(_3732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7547_ (.I0(_3480_),
    .I1(_3732_),
    .S(_3730_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7548_ (.A1(_3726_),
    .A2(\registers[19][21] ),
    .Z(_3733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7549_ (.I0(_3482_),
    .I1(_3733_),
    .S(_3730_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7550_ (.A1(_3726_),
    .A2(\registers[19][22] ),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7551_ (.I0(_3484_),
    .I1(_3734_),
    .S(_3730_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7552_ (.A1(_3726_),
    .A2(\registers[19][23] ),
    .Z(_3735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7553_ (.I0(_3486_),
    .I1(_3735_),
    .S(_3730_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7554_ (.A1(_3726_),
    .A2(\registers[19][24] ),
    .Z(_3736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7555_ (.I0(_3488_),
    .I1(_3736_),
    .S(_3730_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7556_ (.A1(_3726_),
    .A2(\registers[19][25] ),
    .Z(_3737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7557_ (.I0(_3490_),
    .I1(_3737_),
    .S(_3730_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7558_ (.I(_3650_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7559_ (.A1(_3738_),
    .A2(\registers[19][26] ),
    .Z(_3739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7560_ (.I0(_3492_),
    .I1(_3739_),
    .S(_3730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7561_ (.A1(_3738_),
    .A2(\registers[19][27] ),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7562_ (.I0(_3494_),
    .I1(_3740_),
    .S(_3730_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7563_ (.A1(_3738_),
    .A2(\registers[19][28] ),
    .Z(_3741_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7564_ (.I(_3717_),
    .Z(_3742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7565_ (.I0(_3496_),
    .I1(_3741_),
    .S(_3742_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7566_ (.A1(_3738_),
    .A2(\registers[19][29] ),
    .Z(_3743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7567_ (.I0(_3500_),
    .I1(_3743_),
    .S(_3742_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7568_ (.A1(_3738_),
    .A2(\registers[19][2] ),
    .Z(_3744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7569_ (.I0(_3502_),
    .I1(_3744_),
    .S(_3742_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7570_ (.A1(_3738_),
    .A2(\registers[19][30] ),
    .Z(_3745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7571_ (.I0(_3504_),
    .I1(_3745_),
    .S(_3742_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7572_ (.A1(_3738_),
    .A2(\registers[19][31] ),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7573_ (.I0(_3435_),
    .I1(_3746_),
    .S(_3742_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7574_ (.A1(_3738_),
    .A2(\registers[19][3] ),
    .Z(_3747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7575_ (.I0(_3437_),
    .I1(_3747_),
    .S(_3742_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7576_ (.A1(_3738_),
    .A2(\registers[19][4] ),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7577_ (.I0(_3439_),
    .I1(_3748_),
    .S(_3742_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7578_ (.A1(_3738_),
    .A2(\registers[19][5] ),
    .Z(_3749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7579_ (.I0(_3441_),
    .I1(_3749_),
    .S(_3742_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7580_ (.I(_3650_),
    .Z(_3750_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7581_ (.A1(_3750_),
    .A2(\registers[19][6] ),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7582_ (.I0(_3443_),
    .I1(_3751_),
    .S(_3742_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7583_ (.A1(_3750_),
    .A2(\registers[19][7] ),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7584_ (.I0(_3445_),
    .I1(_3752_),
    .S(_3742_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7585_ (.A1(_3750_),
    .A2(\registers[19][8] ),
    .Z(_3753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7586_ (.I0(_3447_),
    .I1(_3753_),
    .S(_3717_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7587_ (.A1(_3750_),
    .A2(\registers[19][9] ),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7588_ (.I0(_3449_),
    .I1(_3754_),
    .S(_3717_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7589_ (.A1(_3750_),
    .A2(\registers[1][0] ),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7590_ (.A1(_1095_),
    .A2(_1116_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7591_ (.I(_3756_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7592_ (.I0(_3451_),
    .I1(_3755_),
    .S(_3757_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7593_ (.A1(_3750_),
    .A2(\registers[1][10] ),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7594_ (.I0(_3456_),
    .I1(_3758_),
    .S(_3757_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7595_ (.A1(_3750_),
    .A2(\registers[1][11] ),
    .Z(_3759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7596_ (.I0(_3458_),
    .I1(_3759_),
    .S(_3757_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7597_ (.A1(_3750_),
    .A2(\registers[1][12] ),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7598_ (.I0(_3460_),
    .I1(_3760_),
    .S(_3757_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7599_ (.A1(_3750_),
    .A2(\registers[1][13] ),
    .Z(_3761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7600_ (.I0(_3462_),
    .I1(_3761_),
    .S(_3757_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7601_ (.A1(_3750_),
    .A2(\registers[1][14] ),
    .Z(_3762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7602_ (.I0(_3464_),
    .I1(_3762_),
    .S(_3757_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7603_ (.I(_3650_),
    .Z(_3763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7604_ (.A1(_3763_),
    .A2(\registers[1][15] ),
    .Z(_3764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7605_ (.I0(_3466_),
    .I1(_3764_),
    .S(_3757_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7606_ (.A1(_3763_),
    .A2(\registers[1][16] ),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7607_ (.I0(_3468_),
    .I1(_3765_),
    .S(_3757_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7608_ (.A1(_3763_),
    .A2(\registers[1][17] ),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7609_ (.I0(_3470_),
    .I1(_3766_),
    .S(_3757_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7610_ (.A1(_3763_),
    .A2(\registers[1][18] ),
    .Z(_3767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7611_ (.I0(_3472_),
    .I1(_3767_),
    .S(_3757_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7612_ (.A1(_3763_),
    .A2(\registers[1][19] ),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7613_ (.I(_3756_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7614_ (.I0(_3474_),
    .I1(_3768_),
    .S(_3769_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7615_ (.A1(_3763_),
    .A2(\registers[1][1] ),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7616_ (.I0(_3478_),
    .I1(_3770_),
    .S(_3769_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7617_ (.A1(_3763_),
    .A2(\registers[1][20] ),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7618_ (.I0(_3480_),
    .I1(_3771_),
    .S(_3769_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7619_ (.A1(_3763_),
    .A2(\registers[1][21] ),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7620_ (.I0(_3482_),
    .I1(_3772_),
    .S(_3769_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7621_ (.A1(_3763_),
    .A2(\registers[1][22] ),
    .Z(_3773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7622_ (.I0(_3484_),
    .I1(_3773_),
    .S(_3769_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7623_ (.A1(_3763_),
    .A2(\registers[1][23] ),
    .Z(_3774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7624_ (.I0(_3486_),
    .I1(_3774_),
    .S(_3769_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7625_ (.I(_1089_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7626_ (.I(_3775_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7627_ (.A1(_3776_),
    .A2(\registers[1][24] ),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7628_ (.I0(_3488_),
    .I1(_3777_),
    .S(_3769_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7629_ (.A1(_3776_),
    .A2(\registers[1][25] ),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7630_ (.I0(_3490_),
    .I1(_3778_),
    .S(_3769_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7631_ (.A1(_3776_),
    .A2(\registers[1][26] ),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7632_ (.I0(_3492_),
    .I1(_3779_),
    .S(_3769_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7633_ (.A1(_3776_),
    .A2(\registers[1][27] ),
    .Z(_3780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7634_ (.I0(_3494_),
    .I1(_3780_),
    .S(_3769_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7635_ (.A1(_3776_),
    .A2(\registers[1][28] ),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7636_ (.I(_3756_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7637_ (.I0(_3496_),
    .I1(_3781_),
    .S(_3782_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7638_ (.A1(_3776_),
    .A2(\registers[1][29] ),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7639_ (.I0(_3500_),
    .I1(_3783_),
    .S(_3782_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7640_ (.A1(_3776_),
    .A2(\registers[1][2] ),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7641_ (.I0(_3502_),
    .I1(_3784_),
    .S(_3782_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7642_ (.A1(_3776_),
    .A2(\registers[1][30] ),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7643_ (.I0(_3504_),
    .I1(_3785_),
    .S(_3782_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7644_ (.A1(_3776_),
    .A2(\registers[1][31] ),
    .Z(_3786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7645_ (.I0(_3435_),
    .I1(_3786_),
    .S(_3782_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7646_ (.A1(_3776_),
    .A2(\registers[1][3] ),
    .Z(_3787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7647_ (.I0(_3437_),
    .I1(_3787_),
    .S(_3782_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7648_ (.I(_3775_),
    .Z(_3788_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7649_ (.A1(_3788_),
    .A2(\registers[1][4] ),
    .Z(_3789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7650_ (.I0(_3439_),
    .I1(_3789_),
    .S(_3782_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7651_ (.A1(_3788_),
    .A2(\registers[1][5] ),
    .Z(_3790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7652_ (.I0(_3441_),
    .I1(_3790_),
    .S(_3782_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7653_ (.A1(_3788_),
    .A2(\registers[1][6] ),
    .Z(_3791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7654_ (.I0(_3443_),
    .I1(_3791_),
    .S(_3782_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7655_ (.A1(_3788_),
    .A2(\registers[1][7] ),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7656_ (.I0(_3445_),
    .I1(_3792_),
    .S(_3782_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7657_ (.A1(_3788_),
    .A2(\registers[1][8] ),
    .Z(_3793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7658_ (.I0(_3447_),
    .I1(_3793_),
    .S(_3756_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7659_ (.A1(_3788_),
    .A2(\registers[1][9] ),
    .Z(_3794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7660_ (.I0(_3449_),
    .I1(_3794_),
    .S(_3756_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7661_ (.A1(_3788_),
    .A2(\registers[20][0] ),
    .Z(_3795_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _7662_ (.A1(net13),
    .A2(_1497_),
    .A3(_1335_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7663_ (.A1(_1338_),
    .A2(_3796_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7664_ (.I(_3797_),
    .Z(_3798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7665_ (.I0(_3451_),
    .I1(_3795_),
    .S(_3798_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7666_ (.A1(_3788_),
    .A2(\registers[20][10] ),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7667_ (.I0(_3456_),
    .I1(_3799_),
    .S(_3798_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7668_ (.A1(_3788_),
    .A2(\registers[20][11] ),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7669_ (.I0(_3458_),
    .I1(_3800_),
    .S(_3798_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7670_ (.A1(_3788_),
    .A2(\registers[20][12] ),
    .Z(_3801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7671_ (.I0(_3460_),
    .I1(_3801_),
    .S(_3798_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7672_ (.I(_3775_),
    .Z(_3802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7673_ (.A1(_3802_),
    .A2(\registers[20][13] ),
    .Z(_3803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7674_ (.I0(_3462_),
    .I1(_3803_),
    .S(_3798_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7675_ (.A1(_3802_),
    .A2(\registers[20][14] ),
    .Z(_3804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7676_ (.I0(_3464_),
    .I1(_3804_),
    .S(_3798_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7677_ (.A1(_3802_),
    .A2(\registers[20][15] ),
    .Z(_3805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7678_ (.I0(_3466_),
    .I1(_3805_),
    .S(_3798_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7679_ (.A1(_3802_),
    .A2(\registers[20][16] ),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7680_ (.I0(_3468_),
    .I1(_3806_),
    .S(_3798_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7681_ (.A1(_3802_),
    .A2(\registers[20][17] ),
    .Z(_3807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7682_ (.I0(_3470_),
    .I1(_3807_),
    .S(_3798_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7683_ (.A1(_3802_),
    .A2(\registers[20][18] ),
    .Z(_3808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7684_ (.I0(_3472_),
    .I1(_3808_),
    .S(_3798_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7685_ (.A1(_3802_),
    .A2(\registers[20][19] ),
    .Z(_3809_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7686_ (.I(_3797_),
    .Z(_3810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7687_ (.I0(_3474_),
    .I1(_3809_),
    .S(_3810_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7688_ (.A1(_3802_),
    .A2(\registers[20][1] ),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7689_ (.I0(_3478_),
    .I1(_3811_),
    .S(_3810_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7690_ (.A1(_3802_),
    .A2(\registers[20][20] ),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7691_ (.I0(_3480_),
    .I1(_3812_),
    .S(_3810_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7692_ (.A1(_3802_),
    .A2(\registers[20][21] ),
    .Z(_3813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7693_ (.I0(_3482_),
    .I1(_3813_),
    .S(_3810_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7694_ (.I(_3775_),
    .Z(_3814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7695_ (.A1(_3814_),
    .A2(\registers[20][22] ),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7696_ (.I0(_3484_),
    .I1(_3815_),
    .S(_3810_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7697_ (.A1(_3814_),
    .A2(\registers[20][23] ),
    .Z(_3816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7698_ (.I0(_3486_),
    .I1(_3816_),
    .S(_3810_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7699_ (.A1(_3814_),
    .A2(\registers[20][24] ),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7700_ (.I0(_3488_),
    .I1(_3817_),
    .S(_3810_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7701_ (.A1(_3814_),
    .A2(\registers[20][25] ),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7702_ (.I0(_3490_),
    .I1(_3818_),
    .S(_3810_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7703_ (.A1(_3814_),
    .A2(\registers[20][26] ),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7704_ (.I0(_3492_),
    .I1(_3819_),
    .S(_3810_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7705_ (.A1(_3814_),
    .A2(\registers[20][27] ),
    .Z(_3820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7706_ (.I0(_3494_),
    .I1(_3820_),
    .S(_3810_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7707_ (.A1(_3814_),
    .A2(\registers[20][28] ),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7708_ (.I(_3797_),
    .Z(_3822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7709_ (.I0(_3496_),
    .I1(_3821_),
    .S(_3822_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7710_ (.A1(_3814_),
    .A2(\registers[20][29] ),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7711_ (.I0(_3500_),
    .I1(_3823_),
    .S(_3822_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7712_ (.A1(_3814_),
    .A2(\registers[20][2] ),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7713_ (.I0(_3502_),
    .I1(_3824_),
    .S(_3822_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7714_ (.A1(_3814_),
    .A2(\registers[20][30] ),
    .Z(_3825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7715_ (.I0(_3504_),
    .I1(_3825_),
    .S(_3822_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7716_ (.I(_3775_),
    .Z(_3826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7717_ (.A1(_3826_),
    .A2(\registers[20][31] ),
    .Z(_3827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7718_ (.I0(_3435_),
    .I1(_3827_),
    .S(_3822_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7719_ (.A1(_3826_),
    .A2(\registers[20][3] ),
    .Z(_3828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7720_ (.I0(_3437_),
    .I1(_3828_),
    .S(_3822_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7721_ (.A1(_3826_),
    .A2(\registers[20][4] ),
    .Z(_3829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7722_ (.I0(_3439_),
    .I1(_3829_),
    .S(_3822_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7723_ (.A1(_3826_),
    .A2(\registers[20][5] ),
    .Z(_3830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7724_ (.I0(_3441_),
    .I1(_3830_),
    .S(_3822_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7725_ (.A1(_3826_),
    .A2(\registers[20][6] ),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7726_ (.I0(_3443_),
    .I1(_3831_),
    .S(_3822_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7727_ (.A1(_3826_),
    .A2(\registers[20][7] ),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7728_ (.I0(_3445_),
    .I1(_3832_),
    .S(_3822_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7729_ (.A1(_3826_),
    .A2(\registers[20][8] ),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7730_ (.I0(_3447_),
    .I1(_3833_),
    .S(_3797_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7731_ (.A1(_3826_),
    .A2(\registers[20][9] ),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7732_ (.I0(_3449_),
    .I1(_3834_),
    .S(_3797_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7733_ (.A1(_3826_),
    .A2(\registers[21][0] ),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7734_ (.A1(_1095_),
    .A2(_3796_),
    .ZN(_3836_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7735_ (.I(_3836_),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7736_ (.I0(_3451_),
    .I1(_3835_),
    .S(_3837_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7737_ (.A1(_3826_),
    .A2(\registers[21][10] ),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7738_ (.I0(_3456_),
    .I1(_3838_),
    .S(_3837_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7739_ (.I(_3775_),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7740_ (.A1(_3839_),
    .A2(\registers[21][11] ),
    .Z(_3840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7741_ (.I0(_3458_),
    .I1(_3840_),
    .S(_3837_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7742_ (.A1(_3839_),
    .A2(\registers[21][12] ),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7743_ (.I0(_3460_),
    .I1(_3841_),
    .S(_3837_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7744_ (.A1(_3839_),
    .A2(\registers[21][13] ),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7745_ (.I0(_3462_),
    .I1(_3842_),
    .S(_3837_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7746_ (.A1(_3839_),
    .A2(\registers[21][14] ),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7747_ (.I0(_3464_),
    .I1(_3843_),
    .S(_3837_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7748_ (.A1(_3839_),
    .A2(\registers[21][15] ),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7749_ (.I0(_3466_),
    .I1(_3844_),
    .S(_3837_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7750_ (.A1(_3839_),
    .A2(\registers[21][16] ),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7751_ (.I0(_3468_),
    .I1(_3845_),
    .S(_3837_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7752_ (.A1(_3839_),
    .A2(\registers[21][17] ),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7753_ (.I0(_3470_),
    .I1(_3846_),
    .S(_3837_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7754_ (.A1(_3839_),
    .A2(\registers[21][18] ),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7755_ (.I0(_3472_),
    .I1(_3847_),
    .S(_3837_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7756_ (.A1(_3839_),
    .A2(\registers[21][19] ),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7757_ (.I(_3836_),
    .Z(_3849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7758_ (.I0(_3474_),
    .I1(_3848_),
    .S(_3849_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7759_ (.A1(_3839_),
    .A2(\registers[21][1] ),
    .Z(_3850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7760_ (.I0(_3478_),
    .I1(_3850_),
    .S(_3849_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7761_ (.I(_3775_),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7762_ (.A1(_3851_),
    .A2(\registers[21][20] ),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7763_ (.I0(_3480_),
    .I1(_3852_),
    .S(_3849_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7764_ (.A1(_3851_),
    .A2(\registers[21][21] ),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7765_ (.I0(_3482_),
    .I1(_3853_),
    .S(_3849_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7766_ (.A1(_3851_),
    .A2(\registers[21][22] ),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7767_ (.I0(_3484_),
    .I1(_3854_),
    .S(_3849_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7768_ (.A1(_3851_),
    .A2(\registers[21][23] ),
    .Z(_3855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7769_ (.I0(_3486_),
    .I1(_3855_),
    .S(_3849_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7770_ (.A1(_3851_),
    .A2(\registers[21][24] ),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7771_ (.I0(_3488_),
    .I1(_3856_),
    .S(_3849_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7772_ (.A1(_3851_),
    .A2(\registers[21][25] ),
    .Z(_3857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7773_ (.I0(_3490_),
    .I1(_3857_),
    .S(_3849_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7774_ (.A1(_3851_),
    .A2(\registers[21][26] ),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7775_ (.I0(_3492_),
    .I1(_3858_),
    .S(_3849_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7776_ (.A1(_3851_),
    .A2(\registers[21][27] ),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7777_ (.I0(_3494_),
    .I1(_3859_),
    .S(_3849_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7778_ (.A1(_3851_),
    .A2(\registers[21][28] ),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7779_ (.I(_3836_),
    .Z(_3861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7780_ (.I0(_3496_),
    .I1(_3860_),
    .S(_3861_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7781_ (.A1(_3851_),
    .A2(\registers[21][29] ),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7782_ (.I0(_3500_),
    .I1(_3862_),
    .S(_3861_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7783_ (.I(_3775_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7784_ (.A1(_3863_),
    .A2(\registers[21][2] ),
    .Z(_3864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7785_ (.I0(_3502_),
    .I1(_3864_),
    .S(_3861_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7786_ (.A1(_3863_),
    .A2(\registers[21][30] ),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7787_ (.I0(_3504_),
    .I1(_3865_),
    .S(_3861_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7788_ (.A1(_3863_),
    .A2(\registers[21][31] ),
    .Z(_3866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7789_ (.I0(_1173_),
    .I1(_3866_),
    .S(_3861_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7790_ (.A1(_3863_),
    .A2(\registers[21][3] ),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7791_ (.I0(_1175_),
    .I1(_3867_),
    .S(_3861_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7792_ (.A1(_3863_),
    .A2(\registers[21][4] ),
    .Z(_3868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7793_ (.I0(_1177_),
    .I1(_3868_),
    .S(_3861_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7794_ (.A1(_3863_),
    .A2(\registers[21][5] ),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7795_ (.I0(_1179_),
    .I1(_3869_),
    .S(_3861_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7796_ (.A1(_3863_),
    .A2(\registers[21][6] ),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7797_ (.I0(_1181_),
    .I1(_3870_),
    .S(_3861_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7798_ (.A1(_3863_),
    .A2(\registers[21][7] ),
    .Z(_3871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7799_ (.I0(_1183_),
    .I1(_3871_),
    .S(_3861_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7800_ (.A1(_3863_),
    .A2(\registers[21][8] ),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7801_ (.I0(_1186_),
    .I1(_3872_),
    .S(_3836_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7802_ (.A1(_3863_),
    .A2(\registers[21][9] ),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7803_ (.I0(_1188_),
    .I1(_3873_),
    .S(_3836_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7804_ (.I(_3775_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7805_ (.A1(_3874_),
    .A2(\registers[22][0] ),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7806_ (.A1(_1119_),
    .A2(_3796_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7807_ (.I(_3876_),
    .Z(_3877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7808_ (.I0(_1115_),
    .I1(_3875_),
    .S(_3877_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7809_ (.A1(_3874_),
    .A2(\registers[22][10] ),
    .Z(_3878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7810_ (.I0(_1123_),
    .I1(_3878_),
    .S(_3877_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7811_ (.A1(_3874_),
    .A2(\registers[22][11] ),
    .Z(_3879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7812_ (.I0(_1125_),
    .I1(_3879_),
    .S(_3877_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7813_ (.A1(_3874_),
    .A2(\registers[22][12] ),
    .Z(_3880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7814_ (.I0(_1127_),
    .I1(_3880_),
    .S(_3877_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7815_ (.A1(_3874_),
    .A2(\registers[22][13] ),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7816_ (.I0(_1129_),
    .I1(_3881_),
    .S(_3877_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7817_ (.A1(_3874_),
    .A2(\registers[22][14] ),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7818_ (.I0(_1131_),
    .I1(_3882_),
    .S(_3877_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7819_ (.A1(_3874_),
    .A2(\registers[22][15] ),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7820_ (.I0(_1133_),
    .I1(_3883_),
    .S(_3877_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7821_ (.A1(_3874_),
    .A2(\registers[22][16] ),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7822_ (.I0(_1135_),
    .I1(_3884_),
    .S(_3877_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7823_ (.A1(_3874_),
    .A2(\registers[22][17] ),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7824_ (.I0(_1137_),
    .I1(_3885_),
    .S(_3877_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7825_ (.A1(_3874_),
    .A2(\registers[22][18] ),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7826_ (.I0(_1139_),
    .I1(_3886_),
    .S(_3877_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7827_ (.I(_3775_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7828_ (.A1(_3887_),
    .A2(\registers[22][19] ),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7829_ (.I(_3876_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7830_ (.I0(_1142_),
    .I1(_3888_),
    .S(_3889_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7831_ (.A1(_3887_),
    .A2(\registers[22][1] ),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7832_ (.I0(_1145_),
    .I1(_3890_),
    .S(_3889_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7833_ (.A1(_3887_),
    .A2(\registers[22][20] ),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7834_ (.I0(_1147_),
    .I1(_3891_),
    .S(_3889_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7835_ (.A1(_3887_),
    .A2(\registers[22][21] ),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7836_ (.I0(_1149_),
    .I1(_3892_),
    .S(_3889_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7837_ (.A1(_3887_),
    .A2(\registers[22][22] ),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7838_ (.I0(_1151_),
    .I1(_3893_),
    .S(_3889_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7839_ (.A1(_3887_),
    .A2(\registers[22][23] ),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7840_ (.I0(_1153_),
    .I1(_3894_),
    .S(_3889_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7841_ (.A1(_3887_),
    .A2(\registers[22][24] ),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7842_ (.I0(_1155_),
    .I1(_3895_),
    .S(_3889_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7843_ (.A1(_3887_),
    .A2(\registers[22][25] ),
    .Z(_3896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7844_ (.I0(_1157_),
    .I1(_3896_),
    .S(_3889_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7845_ (.A1(_3887_),
    .A2(\registers[22][26] ),
    .Z(_3897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7846_ (.I0(_1159_),
    .I1(_3897_),
    .S(_3889_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7847_ (.A1(_3887_),
    .A2(\registers[22][27] ),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7848_ (.I0(_1161_),
    .I1(_3898_),
    .S(_3889_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _7849_ (.I(_1089_),
    .Z(_3899_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7850_ (.I(_3899_),
    .Z(_3900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7851_ (.A1(_3900_),
    .A2(\registers[22][28] ),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7852_ (.I(_3876_),
    .Z(_3902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7853_ (.I0(_1164_),
    .I1(_3901_),
    .S(_3902_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7854_ (.A1(_3900_),
    .A2(\registers[22][29] ),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7855_ (.I0(_1167_),
    .I1(_3903_),
    .S(_3902_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7856_ (.A1(_3900_),
    .A2(\registers[22][2] ),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7857_ (.I0(_1169_),
    .I1(_3904_),
    .S(_3902_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7858_ (.A1(_3900_),
    .A2(\registers[22][30] ),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7859_ (.I0(_1171_),
    .I1(_3905_),
    .S(_3902_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7860_ (.A1(_3900_),
    .A2(\registers[22][31] ),
    .Z(_3906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7861_ (.I0(_1173_),
    .I1(_3906_),
    .S(_3902_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7862_ (.A1(_3900_),
    .A2(\registers[22][3] ),
    .Z(_3907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7863_ (.I0(_1175_),
    .I1(_3907_),
    .S(_3902_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7864_ (.A1(_3900_),
    .A2(\registers[22][4] ),
    .Z(_3908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7865_ (.I0(_1177_),
    .I1(_3908_),
    .S(_3902_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7866_ (.A1(_3900_),
    .A2(\registers[22][5] ),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7867_ (.I0(_1179_),
    .I1(_3909_),
    .S(_3902_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7868_ (.A1(_3900_),
    .A2(\registers[22][6] ),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7869_ (.I0(_1181_),
    .I1(_3910_),
    .S(_3902_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7870_ (.A1(_3900_),
    .A2(\registers[22][7] ),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7871_ (.I0(_1183_),
    .I1(_3911_),
    .S(_3902_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7872_ (.I(_3899_),
    .Z(_3912_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7873_ (.A1(_3912_),
    .A2(\registers[22][8] ),
    .Z(_3913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7874_ (.I0(_1186_),
    .I1(_3913_),
    .S(_3876_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7875_ (.A1(_3912_),
    .A2(\registers[22][9] ),
    .Z(_3914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7876_ (.I0(_1188_),
    .I1(_3914_),
    .S(_3876_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7877_ (.A1(_3394_),
    .A2(\registers[23][0] ),
    .Z(_3915_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _7878_ (.A1(_1232_),
    .A2(_3796_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7879_ (.I(_3916_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7880_ (.I0(_3915_),
    .I1(net15),
    .S(_3917_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7881_ (.A1(_3394_),
    .A2(\registers[23][10] ),
    .Z(_3918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7882_ (.I0(_3918_),
    .I1(net16),
    .S(_3917_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7883_ (.I(_1223_),
    .Z(_3919_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7884_ (.A1(_3919_),
    .A2(\registers[23][11] ),
    .Z(_3920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7885_ (.I0(_3920_),
    .I1(net17),
    .S(_3917_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7886_ (.A1(_3919_),
    .A2(\registers[23][12] ),
    .Z(_3921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7887_ (.I0(_3921_),
    .I1(net18),
    .S(_3917_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7888_ (.A1(_3919_),
    .A2(\registers[23][13] ),
    .Z(_3922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7889_ (.I0(_3922_),
    .I1(net19),
    .S(_3917_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7890_ (.A1(_3919_),
    .A2(\registers[23][14] ),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7891_ (.I0(_3923_),
    .I1(net20),
    .S(_3917_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7892_ (.A1(_3919_),
    .A2(\registers[23][15] ),
    .Z(_3924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7893_ (.I0(_3924_),
    .I1(net21),
    .S(_3917_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7894_ (.A1(_3919_),
    .A2(\registers[23][16] ),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7895_ (.I0(_3925_),
    .I1(net22),
    .S(_3917_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7896_ (.A1(_3919_),
    .A2(\registers[23][17] ),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7897_ (.I0(_3926_),
    .I1(net23),
    .S(_3917_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7898_ (.A1(_3919_),
    .A2(\registers[23][18] ),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7899_ (.I0(_3927_),
    .I1(net24),
    .S(_3917_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7900_ (.A1(_3919_),
    .A2(\registers[23][19] ),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7901_ (.I(_3916_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7902_ (.I0(_3928_),
    .I1(net25),
    .S(_3929_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7903_ (.A1(_3919_),
    .A2(\registers[23][1] ),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7904_ (.I0(_3930_),
    .I1(net26),
    .S(_3929_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7905_ (.I(_1223_),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7906_ (.A1(_3931_),
    .A2(\registers[23][20] ),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7907_ (.I0(_3932_),
    .I1(net27),
    .S(_3929_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7908_ (.A1(_3931_),
    .A2(\registers[23][21] ),
    .Z(_3933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7909_ (.I0(_3933_),
    .I1(net28),
    .S(_3929_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7910_ (.A1(_3931_),
    .A2(\registers[23][22] ),
    .Z(_3934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7911_ (.I0(_3934_),
    .I1(net29),
    .S(_3929_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7912_ (.A1(_3931_),
    .A2(\registers[23][23] ),
    .Z(_3935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7913_ (.I0(_3935_),
    .I1(net30),
    .S(_3929_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7914_ (.A1(_3931_),
    .A2(\registers[23][24] ),
    .Z(_3936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7915_ (.I0(_3936_),
    .I1(net31),
    .S(_3929_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7916_ (.A1(_3931_),
    .A2(\registers[23][25] ),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7917_ (.I0(_3937_),
    .I1(net32),
    .S(_3929_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7918_ (.A1(_3931_),
    .A2(\registers[23][26] ),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7919_ (.I0(_3938_),
    .I1(net33),
    .S(_3929_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7920_ (.A1(_3931_),
    .A2(\registers[23][27] ),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7921_ (.I0(_3939_),
    .I1(net34),
    .S(_3929_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7922_ (.A1(_3931_),
    .A2(\registers[23][28] ),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7923_ (.I(_3916_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7924_ (.I0(_3940_),
    .I1(net35),
    .S(_3941_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7925_ (.A1(_3931_),
    .A2(\registers[23][29] ),
    .Z(_3942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7926_ (.I0(_3942_),
    .I1(net36),
    .S(_3941_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _7927_ (.I(_1223_),
    .Z(_3943_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7928_ (.A1(_3943_),
    .A2(\registers[23][2] ),
    .Z(_3944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7929_ (.I0(_3944_),
    .I1(net37),
    .S(_3941_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7930_ (.A1(_3943_),
    .A2(\registers[23][30] ),
    .Z(_3945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7931_ (.I0(_3945_),
    .I1(net38),
    .S(_3941_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7932_ (.A1(_3943_),
    .A2(\registers[23][31] ),
    .Z(_3946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7933_ (.I0(_3946_),
    .I1(net39),
    .S(_3941_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7934_ (.A1(_3943_),
    .A2(\registers[23][3] ),
    .Z(_3947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7935_ (.I0(_3947_),
    .I1(net40),
    .S(_3941_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7936_ (.A1(_3943_),
    .A2(\registers[23][4] ),
    .Z(_3948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7937_ (.I0(_3948_),
    .I1(net41),
    .S(_3941_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7938_ (.A1(_3943_),
    .A2(\registers[23][5] ),
    .Z(_3949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7939_ (.I0(_3949_),
    .I1(net42),
    .S(_3941_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7940_ (.A1(_3943_),
    .A2(\registers[23][6] ),
    .Z(_3950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7941_ (.I0(_3950_),
    .I1(net43),
    .S(_3941_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7942_ (.A1(_3943_),
    .A2(\registers[23][7] ),
    .Z(_3951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7943_ (.I0(_3951_),
    .I1(net44),
    .S(_3941_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7944_ (.A1(_3943_),
    .A2(\registers[23][8] ),
    .Z(_3952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7945_ (.I0(_3952_),
    .I1(net45),
    .S(_3916_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7946_ (.A1(_3943_),
    .A2(\registers[23][9] ),
    .Z(_3953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7947_ (.I0(_3953_),
    .I1(net46),
    .S(_3916_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7948_ (.A1(_3912_),
    .A2(\registers[24][0] ),
    .Z(_3954_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _7949_ (.A1(net13),
    .A2(net14),
    .A3(_1335_),
    .Z(_3955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _7950_ (.A1(_1338_),
    .A2(_3955_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7951_ (.I(_3956_),
    .Z(_3957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7952_ (.I0(_1115_),
    .I1(_3954_),
    .S(_3957_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7953_ (.A1(_3912_),
    .A2(\registers[24][10] ),
    .Z(_3958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7954_ (.I0(_1123_),
    .I1(_3958_),
    .S(_3957_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7955_ (.A1(_3912_),
    .A2(\registers[24][11] ),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7956_ (.I0(_1125_),
    .I1(_3959_),
    .S(_3957_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7957_ (.A1(_3912_),
    .A2(\registers[24][12] ),
    .Z(_3960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7958_ (.I0(_1127_),
    .I1(_3960_),
    .S(_3957_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7959_ (.A1(_3912_),
    .A2(\registers[24][13] ),
    .Z(_3961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7960_ (.I0(_1129_),
    .I1(_3961_),
    .S(_3957_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7961_ (.A1(_3912_),
    .A2(\registers[24][14] ),
    .Z(_3962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7962_ (.I0(_1131_),
    .I1(_3962_),
    .S(_3957_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7963_ (.A1(_3912_),
    .A2(\registers[24][15] ),
    .Z(_3963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7964_ (.I0(_1133_),
    .I1(_3963_),
    .S(_3957_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7965_ (.A1(_3912_),
    .A2(\registers[24][16] ),
    .Z(_3964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7966_ (.I0(_1135_),
    .I1(_3964_),
    .S(_3957_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7967_ (.I(_3899_),
    .Z(_3965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7968_ (.A1(_3965_),
    .A2(\registers[24][17] ),
    .Z(_3966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7969_ (.I0(_1137_),
    .I1(_3966_),
    .S(_3957_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7970_ (.A1(_3965_),
    .A2(\registers[24][18] ),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7971_ (.I0(_1139_),
    .I1(_3967_),
    .S(_3957_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7972_ (.A1(_3965_),
    .A2(\registers[24][19] ),
    .Z(_3968_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _7973_ (.I(_3956_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7974_ (.I0(_1142_),
    .I1(_3968_),
    .S(_3969_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7975_ (.A1(_3965_),
    .A2(\registers[24][1] ),
    .Z(_3970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7976_ (.I0(_1145_),
    .I1(_3970_),
    .S(_3969_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7977_ (.A1(_3965_),
    .A2(\registers[24][20] ),
    .Z(_3971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7978_ (.I0(_1147_),
    .I1(_3971_),
    .S(_3969_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7979_ (.A1(_3965_),
    .A2(\registers[24][21] ),
    .Z(_3972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7980_ (.I0(_1149_),
    .I1(_3972_),
    .S(_3969_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7981_ (.A1(_3965_),
    .A2(\registers[24][22] ),
    .Z(_3973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7982_ (.I0(_1151_),
    .I1(_3973_),
    .S(_3969_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7983_ (.A1(_3965_),
    .A2(\registers[24][23] ),
    .Z(_3974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7984_ (.I0(_1153_),
    .I1(_3974_),
    .S(_3969_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7985_ (.A1(_3965_),
    .A2(\registers[24][24] ),
    .Z(_3975_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7986_ (.I0(_1155_),
    .I1(_3975_),
    .S(_3969_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7987_ (.A1(_3965_),
    .A2(\registers[24][25] ),
    .Z(_3976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7988_ (.I0(_1157_),
    .I1(_3976_),
    .S(_3969_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7989_ (.I(_3899_),
    .Z(_3977_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7990_ (.A1(_3977_),
    .A2(\registers[24][26] ),
    .Z(_3978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7991_ (.I0(_1159_),
    .I1(_3978_),
    .S(_3969_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7992_ (.A1(_3977_),
    .A2(\registers[24][27] ),
    .Z(_3979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7993_ (.I0(_1161_),
    .I1(_3979_),
    .S(_3969_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7994_ (.A1(_3977_),
    .A2(\registers[24][28] ),
    .Z(_3980_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _7995_ (.I(_3956_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7996_ (.I0(_1164_),
    .I1(_3980_),
    .S(_3981_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7997_ (.A1(_3977_),
    .A2(\registers[24][29] ),
    .Z(_3982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _7998_ (.I0(_1167_),
    .I1(_3982_),
    .S(_3981_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _7999_ (.A1(_3977_),
    .A2(\registers[24][2] ),
    .Z(_3983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8000_ (.I0(_1169_),
    .I1(_3983_),
    .S(_3981_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8001_ (.A1(_3977_),
    .A2(\registers[24][30] ),
    .Z(_3984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8002_ (.I0(_1171_),
    .I1(_3984_),
    .S(_3981_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8003_ (.A1(_3977_),
    .A2(\registers[24][31] ),
    .Z(_3985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8004_ (.I0(_1173_),
    .I1(_3985_),
    .S(_3981_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8005_ (.A1(_3977_),
    .A2(\registers[24][3] ),
    .Z(_3986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8006_ (.I0(_1175_),
    .I1(_3986_),
    .S(_3981_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8007_ (.A1(_3977_),
    .A2(\registers[24][4] ),
    .Z(_3987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8008_ (.I0(_1177_),
    .I1(_3987_),
    .S(_3981_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8009_ (.A1(_3977_),
    .A2(\registers[24][5] ),
    .Z(_3988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8010_ (.I0(_1179_),
    .I1(_3988_),
    .S(_3981_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8011_ (.I(_3899_),
    .Z(_3989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8012_ (.A1(_3989_),
    .A2(\registers[24][6] ),
    .Z(_3990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8013_ (.I0(_1181_),
    .I1(_3990_),
    .S(_3981_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8014_ (.A1(_3989_),
    .A2(\registers[24][7] ),
    .Z(_3991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8015_ (.I0(_1183_),
    .I1(_3991_),
    .S(_3981_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8016_ (.A1(_3989_),
    .A2(\registers[24][8] ),
    .Z(_3992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8017_ (.I0(_1186_),
    .I1(_3992_),
    .S(_3956_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8018_ (.A1(_3989_),
    .A2(\registers[24][9] ),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8019_ (.I0(_1188_),
    .I1(_3993_),
    .S(_3956_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8020_ (.A1(_3989_),
    .A2(\registers[25][0] ),
    .Z(_3994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _8021_ (.A1(_1095_),
    .A2(_3955_),
    .ZN(_3995_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8022_ (.I(_3995_),
    .Z(_3996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8023_ (.I0(_1115_),
    .I1(_3994_),
    .S(_3996_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8024_ (.A1(_3989_),
    .A2(\registers[25][10] ),
    .Z(_3997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8025_ (.I0(_1123_),
    .I1(_3997_),
    .S(_3996_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8026_ (.A1(_3989_),
    .A2(\registers[25][11] ),
    .Z(_3998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8027_ (.I0(_1125_),
    .I1(_3998_),
    .S(_3996_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8028_ (.A1(_3989_),
    .A2(\registers[25][12] ),
    .Z(_3999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8029_ (.I0(_1127_),
    .I1(_3999_),
    .S(_3996_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8030_ (.A1(_3989_),
    .A2(\registers[25][13] ),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8031_ (.I0(_1129_),
    .I1(_4000_),
    .S(_3996_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8032_ (.A1(_3989_),
    .A2(\registers[25][14] ),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8033_ (.I0(_1131_),
    .I1(_4001_),
    .S(_3996_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8034_ (.I(_3899_),
    .Z(_4002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8035_ (.A1(_4002_),
    .A2(\registers[25][15] ),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8036_ (.I0(_1133_),
    .I1(_4003_),
    .S(_3996_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8037_ (.A1(_4002_),
    .A2(\registers[25][16] ),
    .Z(_4004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8038_ (.I0(_1135_),
    .I1(_4004_),
    .S(_3996_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8039_ (.A1(_4002_),
    .A2(\registers[25][17] ),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8040_ (.I0(_1137_),
    .I1(_4005_),
    .S(_3996_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8041_ (.A1(_4002_),
    .A2(\registers[25][18] ),
    .Z(_4006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8042_ (.I0(_1139_),
    .I1(_4006_),
    .S(_3996_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8043_ (.A1(_4002_),
    .A2(\registers[25][19] ),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8044_ (.I(_3995_),
    .Z(_4008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8045_ (.I0(_1142_),
    .I1(_4007_),
    .S(_4008_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8046_ (.A1(_4002_),
    .A2(\registers[25][1] ),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8047_ (.I0(_1145_),
    .I1(_4009_),
    .S(_4008_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8048_ (.A1(_4002_),
    .A2(\registers[25][20] ),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8049_ (.I0(_1147_),
    .I1(_4010_),
    .S(_4008_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8050_ (.A1(_4002_),
    .A2(\registers[25][21] ),
    .Z(_4011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8051_ (.I0(_1149_),
    .I1(_4011_),
    .S(_4008_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8052_ (.A1(_4002_),
    .A2(\registers[25][22] ),
    .Z(_4012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8053_ (.I0(_1151_),
    .I1(_4012_),
    .S(_4008_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8054_ (.A1(_4002_),
    .A2(\registers[25][23] ),
    .Z(_4013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8055_ (.I0(_1153_),
    .I1(_4013_),
    .S(_4008_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8056_ (.I(_3899_),
    .Z(_4014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8057_ (.A1(_4014_),
    .A2(\registers[25][24] ),
    .Z(_4015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8058_ (.I0(_1155_),
    .I1(_4015_),
    .S(_4008_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8059_ (.A1(_4014_),
    .A2(\registers[25][25] ),
    .Z(_4016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8060_ (.I0(_1157_),
    .I1(_4016_),
    .S(_4008_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8061_ (.A1(_4014_),
    .A2(\registers[25][26] ),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8062_ (.I0(_1159_),
    .I1(_4017_),
    .S(_4008_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8063_ (.A1(_4014_),
    .A2(\registers[25][27] ),
    .Z(_4018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8064_ (.I0(_1161_),
    .I1(_4018_),
    .S(_4008_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8065_ (.A1(_4014_),
    .A2(\registers[25][28] ),
    .Z(_4019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8066_ (.I(_3995_),
    .Z(_4020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8067_ (.I0(_1164_),
    .I1(_4019_),
    .S(_4020_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8068_ (.A1(_4014_),
    .A2(\registers[25][29] ),
    .Z(_4021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8069_ (.I0(_1167_),
    .I1(_4021_),
    .S(_4020_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8070_ (.A1(_4014_),
    .A2(\registers[25][2] ),
    .Z(_4022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8071_ (.I0(_1169_),
    .I1(_4022_),
    .S(_4020_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8072_ (.A1(_4014_),
    .A2(\registers[25][30] ),
    .Z(_4023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8073_ (.I0(_1171_),
    .I1(_4023_),
    .S(_4020_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8074_ (.A1(_4014_),
    .A2(\registers[25][31] ),
    .Z(_4024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8075_ (.I0(_1173_),
    .I1(_4024_),
    .S(_4020_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8076_ (.A1(_4014_),
    .A2(\registers[25][3] ),
    .Z(_4025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8077_ (.I0(_1175_),
    .I1(_4025_),
    .S(_4020_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8078_ (.I(_3899_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8079_ (.A1(_4026_),
    .A2(\registers[25][4] ),
    .Z(_4027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8080_ (.I0(_1177_),
    .I1(_4027_),
    .S(_4020_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8081_ (.A1(_4026_),
    .A2(\registers[25][5] ),
    .Z(_4028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8082_ (.I0(_1179_),
    .I1(_4028_),
    .S(_4020_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8083_ (.A1(_4026_),
    .A2(\registers[25][6] ),
    .Z(_4029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8084_ (.I0(_1181_),
    .I1(_4029_),
    .S(_4020_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8085_ (.A1(_4026_),
    .A2(\registers[25][7] ),
    .Z(_4030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8086_ (.I0(_1183_),
    .I1(_4030_),
    .S(_4020_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8087_ (.A1(_4026_),
    .A2(\registers[25][8] ),
    .Z(_4031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8088_ (.I0(_1186_),
    .I1(_4031_),
    .S(_3995_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8089_ (.A1(_4026_),
    .A2(\registers[25][9] ),
    .Z(_4032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8090_ (.I0(_1188_),
    .I1(_4032_),
    .S(_3995_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8091_ (.A1(_4026_),
    .A2(\registers[26][0] ),
    .Z(_4033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _8092_ (.A1(_1119_),
    .A2(_3955_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8093_ (.I(_4034_),
    .Z(_4035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8094_ (.I0(_1115_),
    .I1(_4033_),
    .S(_4035_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8095_ (.A1(_4026_),
    .A2(\registers[26][10] ),
    .Z(_4036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8096_ (.I0(_1123_),
    .I1(_4036_),
    .S(_4035_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8097_ (.A1(_4026_),
    .A2(\registers[26][11] ),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8098_ (.I0(_1125_),
    .I1(_4037_),
    .S(_4035_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8099_ (.A1(_4026_),
    .A2(\registers[26][12] ),
    .Z(_4038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8100_ (.I0(_1127_),
    .I1(_4038_),
    .S(_4035_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8101_ (.I(_3899_),
    .Z(_4039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8102_ (.A1(_4039_),
    .A2(\registers[26][13] ),
    .Z(_4040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8103_ (.I0(_1129_),
    .I1(_4040_),
    .S(_4035_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8104_ (.A1(_4039_),
    .A2(\registers[26][14] ),
    .Z(_4041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8105_ (.I0(_1131_),
    .I1(_4041_),
    .S(_4035_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8106_ (.A1(_4039_),
    .A2(\registers[26][15] ),
    .Z(_4042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8107_ (.I0(_1133_),
    .I1(_4042_),
    .S(_4035_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8108_ (.A1(_4039_),
    .A2(\registers[26][16] ),
    .Z(_4043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8109_ (.I0(_1135_),
    .I1(_4043_),
    .S(_4035_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8110_ (.A1(_4039_),
    .A2(\registers[26][17] ),
    .Z(_4044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8111_ (.I0(_1137_),
    .I1(_4044_),
    .S(_4035_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8112_ (.A1(_4039_),
    .A2(\registers[26][18] ),
    .Z(_4045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8113_ (.I0(_1139_),
    .I1(_4045_),
    .S(_4035_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8114_ (.A1(_4039_),
    .A2(\registers[26][19] ),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8115_ (.I(_4034_),
    .Z(_4047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8116_ (.I0(_1142_),
    .I1(_4046_),
    .S(_4047_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8117_ (.A1(_4039_),
    .A2(\registers[26][1] ),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8118_ (.I0(_1145_),
    .I1(_4048_),
    .S(_4047_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8119_ (.A1(_4039_),
    .A2(\registers[26][20] ),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8120_ (.I0(_1147_),
    .I1(_4049_),
    .S(_4047_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8121_ (.A1(_4039_),
    .A2(\registers[26][21] ),
    .Z(_4050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8122_ (.I0(_1149_),
    .I1(_4050_),
    .S(_4047_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8123_ (.I(_3899_),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8124_ (.A1(_4051_),
    .A2(\registers[26][22] ),
    .Z(_4052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8125_ (.I0(_1151_),
    .I1(_4052_),
    .S(_4047_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8126_ (.A1(_4051_),
    .A2(\registers[26][23] ),
    .Z(_4053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8127_ (.I0(_1153_),
    .I1(_4053_),
    .S(_4047_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8128_ (.A1(_4051_),
    .A2(\registers[26][24] ),
    .Z(_4054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8129_ (.I0(_1155_),
    .I1(_4054_),
    .S(_4047_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8130_ (.A1(_4051_),
    .A2(\registers[26][25] ),
    .Z(_4055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8131_ (.I0(_1157_),
    .I1(_4055_),
    .S(_4047_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8132_ (.A1(_4051_),
    .A2(\registers[26][26] ),
    .Z(_4056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8133_ (.I0(_1159_),
    .I1(_4056_),
    .S(_4047_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8134_ (.A1(_4051_),
    .A2(\registers[26][27] ),
    .Z(_4057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8135_ (.I0(_1161_),
    .I1(_4057_),
    .S(_4047_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8136_ (.A1(_4051_),
    .A2(\registers[26][28] ),
    .Z(_4058_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8137_ (.I(_4034_),
    .Z(_4059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8138_ (.I0(_1164_),
    .I1(_4058_),
    .S(_4059_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8139_ (.A1(_4051_),
    .A2(\registers[26][29] ),
    .Z(_4060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8140_ (.I0(_1167_),
    .I1(_4060_),
    .S(_4059_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8141_ (.A1(_4051_),
    .A2(\registers[26][2] ),
    .Z(_4061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8142_ (.I0(_1169_),
    .I1(_4061_),
    .S(_4059_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8143_ (.A1(_4051_),
    .A2(\registers[26][30] ),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8144_ (.I0(_1171_),
    .I1(_4062_),
    .S(_4059_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8145_ (.I(_1639_),
    .Z(_4063_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8146_ (.A1(_4063_),
    .A2(\registers[26][31] ),
    .Z(_4064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8147_ (.I0(_1173_),
    .I1(_4064_),
    .S(_4059_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8148_ (.A1(_4063_),
    .A2(\registers[26][3] ),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8149_ (.I0(_1175_),
    .I1(_4065_),
    .S(_4059_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8150_ (.A1(_4063_),
    .A2(\registers[26][4] ),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8151_ (.I0(_1177_),
    .I1(_4066_),
    .S(_4059_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8152_ (.A1(_4063_),
    .A2(\registers[26][5] ),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8153_ (.I0(_1179_),
    .I1(_4067_),
    .S(_4059_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8154_ (.A1(_4063_),
    .A2(\registers[26][6] ),
    .Z(_4068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8155_ (.I0(_1181_),
    .I1(_4068_),
    .S(_4059_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8156_ (.A1(_4063_),
    .A2(\registers[26][7] ),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8157_ (.I0(_1183_),
    .I1(_4069_),
    .S(_4059_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8158_ (.A1(_4063_),
    .A2(\registers[26][8] ),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8159_ (.I0(_1186_),
    .I1(_4070_),
    .S(_4034_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8160_ (.A1(_4063_),
    .A2(\registers[26][9] ),
    .Z(_4071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8161_ (.I0(_1188_),
    .I1(_4071_),
    .S(_4034_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8162_ (.I(_1090_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8163_ (.A1(_4072_),
    .A2(\registers[27][0] ),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _8164_ (.A1(_1232_),
    .A2(_3955_),
    .Z(_4074_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8165_ (.I(_4074_),
    .Z(_4075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8166_ (.I0(_4073_),
    .I1(net15),
    .S(_4075_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8167_ (.A1(_4072_),
    .A2(\registers[27][10] ),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8168_ (.I0(_4076_),
    .I1(net16),
    .S(_4075_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8169_ (.A1(_4072_),
    .A2(\registers[27][11] ),
    .Z(_4077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8170_ (.I0(_4077_),
    .I1(net17),
    .S(_4075_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8171_ (.A1(_4072_),
    .A2(\registers[27][12] ),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8172_ (.I0(_4078_),
    .I1(net18),
    .S(_4075_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8173_ (.A1(_4072_),
    .A2(\registers[27][13] ),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8174_ (.I0(_4079_),
    .I1(net19),
    .S(_4075_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8175_ (.A1(_4072_),
    .A2(\registers[27][14] ),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8176_ (.I0(_4080_),
    .I1(net20),
    .S(_4075_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8177_ (.A1(_4072_),
    .A2(\registers[27][15] ),
    .Z(_4081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8178_ (.I0(_4081_),
    .I1(net21),
    .S(_4075_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8179_ (.A1(_4072_),
    .A2(\registers[27][16] ),
    .Z(_4082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8180_ (.I0(_4082_),
    .I1(net22),
    .S(_4075_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8181_ (.A1(_4072_),
    .A2(\registers[27][17] ),
    .Z(_4083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8182_ (.I0(_4083_),
    .I1(net23),
    .S(_4075_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8183_ (.A1(_4072_),
    .A2(\registers[27][18] ),
    .Z(_4084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8184_ (.I0(_4084_),
    .I1(net24),
    .S(_4075_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8185_ (.I(_1090_),
    .Z(_4085_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8186_ (.A1(_4085_),
    .A2(\registers[27][19] ),
    .Z(_4086_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8187_ (.I(_4074_),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8188_ (.I0(_4086_),
    .I1(net25),
    .S(_4087_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8189_ (.A1(_4085_),
    .A2(\registers[27][1] ),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8190_ (.I0(_4088_),
    .I1(net26),
    .S(_4087_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8191_ (.A1(_4085_),
    .A2(\registers[27][20] ),
    .Z(_4089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8192_ (.I0(_4089_),
    .I1(net27),
    .S(_4087_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8193_ (.A1(_4085_),
    .A2(\registers[27][21] ),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8194_ (.I0(_4090_),
    .I1(net28),
    .S(_4087_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8195_ (.A1(_4085_),
    .A2(\registers[27][22] ),
    .Z(_4091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8196_ (.I0(_4091_),
    .I1(net29),
    .S(_4087_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8197_ (.A1(_4085_),
    .A2(\registers[27][23] ),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8198_ (.I0(_4092_),
    .I1(net30),
    .S(_4087_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8199_ (.A1(_4085_),
    .A2(\registers[27][24] ),
    .Z(_4093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8200_ (.I0(_4093_),
    .I1(net31),
    .S(_4087_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8201_ (.A1(_4085_),
    .A2(\registers[27][25] ),
    .Z(_4094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8202_ (.I0(_4094_),
    .I1(net32),
    .S(_4087_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8203_ (.A1(_4085_),
    .A2(\registers[27][26] ),
    .Z(_4095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8204_ (.I0(_4095_),
    .I1(net33),
    .S(_4087_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8205_ (.A1(_4085_),
    .A2(\registers[27][27] ),
    .Z(_4096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8206_ (.I0(_4096_),
    .I1(net34),
    .S(_4087_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8207_ (.I(_1090_),
    .Z(_4097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8208_ (.A1(_4097_),
    .A2(\registers[27][28] ),
    .Z(_4098_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8209_ (.I(_4074_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8210_ (.I0(_4098_),
    .I1(net35),
    .S(_4099_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8211_ (.A1(_4097_),
    .A2(\registers[27][29] ),
    .Z(_4100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8212_ (.I0(_4100_),
    .I1(net36),
    .S(_4099_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8213_ (.A1(_4097_),
    .A2(\registers[27][2] ),
    .Z(_4101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8214_ (.I0(_4101_),
    .I1(net37),
    .S(_4099_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8215_ (.A1(_4097_),
    .A2(\registers[27][30] ),
    .Z(_4102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8216_ (.I0(_4102_),
    .I1(net38),
    .S(_4099_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8217_ (.A1(_4097_),
    .A2(\registers[27][31] ),
    .Z(_4103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8218_ (.I0(_4103_),
    .I1(net39),
    .S(_4099_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8219_ (.A1(_4097_),
    .A2(\registers[27][3] ),
    .Z(_4104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8220_ (.I0(_4104_),
    .I1(net40),
    .S(_4099_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8221_ (.A1(_4097_),
    .A2(\registers[27][4] ),
    .Z(_4105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8222_ (.I0(_4105_),
    .I1(net41),
    .S(_4099_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8223_ (.A1(_4097_),
    .A2(\registers[27][5] ),
    .Z(_4106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8224_ (.I0(_4106_),
    .I1(net42),
    .S(_4099_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8225_ (.A1(_4097_),
    .A2(\registers[27][6] ),
    .Z(_4107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8226_ (.I0(_4107_),
    .I1(net43),
    .S(_4099_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8227_ (.A1(_4097_),
    .A2(\registers[27][7] ),
    .Z(_4108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8228_ (.I0(_4108_),
    .I1(net44),
    .S(_4099_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8229_ (.A1(_1091_),
    .A2(\registers[27][8] ),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8230_ (.I0(_4109_),
    .I1(net45),
    .S(_4074_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8231_ (.A1(_1091_),
    .A2(\registers[27][9] ),
    .Z(_4110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8232_ (.I0(_4110_),
    .I1(net46),
    .S(_4074_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8233_ (.A1(_4063_),
    .A2(\registers[28][0] ),
    .Z(_4111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _8234_ (.A1(_1093_),
    .A2(_1338_),
    .ZN(_4112_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8235_ (.I(_4112_),
    .Z(_4113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8236_ (.I0(_1115_),
    .I1(_4111_),
    .S(_4113_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8237_ (.A1(_4063_),
    .A2(\registers[28][10] ),
    .Z(_4114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8238_ (.I0(_1123_),
    .I1(_4114_),
    .S(_4113_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8239_ (.I(_1639_),
    .Z(_4115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8240_ (.A1(_4115_),
    .A2(\registers[28][11] ),
    .Z(_4116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8241_ (.I0(_1125_),
    .I1(_4116_),
    .S(_4113_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8242_ (.A1(_4115_),
    .A2(\registers[28][12] ),
    .Z(_4117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8243_ (.I0(_1127_),
    .I1(_4117_),
    .S(_4113_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8244_ (.A1(_4115_),
    .A2(\registers[28][13] ),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8245_ (.I0(_1129_),
    .I1(_4118_),
    .S(_4113_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8246_ (.A1(_4115_),
    .A2(\registers[28][14] ),
    .Z(_4119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8247_ (.I0(_1131_),
    .I1(_4119_),
    .S(_4113_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8248_ (.A1(_4115_),
    .A2(\registers[28][15] ),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8249_ (.I0(_1133_),
    .I1(_4120_),
    .S(_4113_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8250_ (.A1(_4115_),
    .A2(\registers[28][16] ),
    .Z(_4121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8251_ (.I0(_1135_),
    .I1(_4121_),
    .S(_4113_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8252_ (.A1(_4115_),
    .A2(\registers[28][17] ),
    .Z(_4122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8253_ (.I0(_1137_),
    .I1(_4122_),
    .S(_4113_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8254_ (.A1(_4115_),
    .A2(\registers[28][18] ),
    .Z(_4123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8255_ (.I0(_1139_),
    .I1(_4123_),
    .S(_4113_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8256_ (.A1(_4115_),
    .A2(\registers[28][19] ),
    .Z(_4124_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8257_ (.I(_4112_),
    .Z(_4125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8258_ (.I0(_1142_),
    .I1(_4124_),
    .S(_4125_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8259_ (.A1(_4115_),
    .A2(\registers[28][1] ),
    .Z(_4126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8260_ (.I0(_1145_),
    .I1(_4126_),
    .S(_4125_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8261_ (.I(_1639_),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8262_ (.A1(_4127_),
    .A2(\registers[28][20] ),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8263_ (.I0(_1147_),
    .I1(_4128_),
    .S(_4125_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8264_ (.A1(_4127_),
    .A2(\registers[28][21] ),
    .Z(_4129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8265_ (.I0(_1149_),
    .I1(_4129_),
    .S(_4125_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8266_ (.A1(_4127_),
    .A2(\registers[28][22] ),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8267_ (.I0(_1151_),
    .I1(_4130_),
    .S(_4125_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8268_ (.A1(_4127_),
    .A2(\registers[28][23] ),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8269_ (.I0(_1153_),
    .I1(_4131_),
    .S(_4125_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8270_ (.A1(_4127_),
    .A2(\registers[28][24] ),
    .Z(_4132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8271_ (.I0(_1155_),
    .I1(_4132_),
    .S(_4125_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8272_ (.A1(_4127_),
    .A2(\registers[28][25] ),
    .Z(_4133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8273_ (.I0(_1157_),
    .I1(_4133_),
    .S(_4125_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8274_ (.A1(_4127_),
    .A2(\registers[28][26] ),
    .Z(_4134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8275_ (.I0(_1159_),
    .I1(_4134_),
    .S(_4125_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8276_ (.A1(_4127_),
    .A2(\registers[28][27] ),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8277_ (.I0(_1161_),
    .I1(_4135_),
    .S(_4125_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8278_ (.A1(_4127_),
    .A2(\registers[28][28] ),
    .Z(_4136_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _8279_ (.I(_4112_),
    .Z(_4137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8280_ (.I0(_1164_),
    .I1(_4136_),
    .S(_4137_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8281_ (.A1(_4127_),
    .A2(\registers[28][29] ),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8282_ (.I0(_1167_),
    .I1(_4138_),
    .S(_4137_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8283_ (.I(_1639_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8284_ (.A1(_4139_),
    .A2(\registers[28][2] ),
    .Z(_4140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8285_ (.I0(_1169_),
    .I1(_4140_),
    .S(_4137_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8286_ (.A1(_4139_),
    .A2(\registers[28][30] ),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8287_ (.I0(_1171_),
    .I1(_4141_),
    .S(_4137_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8288_ (.A1(_4139_),
    .A2(\registers[28][31] ),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8289_ (.I0(_1173_),
    .I1(_4142_),
    .S(_4137_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8290_ (.A1(_4139_),
    .A2(\registers[28][3] ),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8291_ (.I0(_1175_),
    .I1(_4143_),
    .S(_4137_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8292_ (.A1(_4139_),
    .A2(\registers[28][4] ),
    .Z(_4144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8293_ (.I0(_1177_),
    .I1(_4144_),
    .S(_4137_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8294_ (.A1(_4139_),
    .A2(\registers[28][5] ),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8295_ (.I0(_1179_),
    .I1(_4145_),
    .S(_4137_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8296_ (.A1(_4139_),
    .A2(\registers[28][6] ),
    .Z(_4146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8297_ (.I0(_1181_),
    .I1(_4146_),
    .S(_4137_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8298_ (.A1(_4139_),
    .A2(\registers[28][7] ),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8299_ (.I0(_1183_),
    .I1(_4147_),
    .S(_4137_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8300_ (.A1(_4139_),
    .A2(\registers[28][8] ),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8301_ (.I0(_1186_),
    .I1(_4148_),
    .S(_4112_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8302_ (.A1(_4139_),
    .A2(\registers[28][9] ),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8303_ (.I0(_1188_),
    .I1(_4149_),
    .S(_4112_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8304_ (.I(_1639_),
    .Z(_4150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8305_ (.A1(_4150_),
    .A2(\registers[29][0] ),
    .Z(_4151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8306_ (.I0(_1115_),
    .I1(_4151_),
    .S(_1097_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8307_ (.A1(_4150_),
    .A2(\registers[29][10] ),
    .Z(_4152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8308_ (.I0(_1123_),
    .I1(_4152_),
    .S(_1097_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8309_ (.A1(_4150_),
    .A2(\registers[29][11] ),
    .Z(_4153_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8310_ (.I(_1096_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8311_ (.I0(_1125_),
    .I1(_4153_),
    .S(_4154_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8312_ (.A1(_4150_),
    .A2(\registers[29][12] ),
    .Z(_4155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8313_ (.I0(_1127_),
    .I1(_4155_),
    .S(_4154_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8314_ (.A1(_4150_),
    .A2(\registers[29][13] ),
    .Z(_4156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8315_ (.I0(_1129_),
    .I1(_4156_),
    .S(_4154_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8316_ (.A1(_4150_),
    .A2(\registers[29][14] ),
    .Z(_4157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8317_ (.I0(_1131_),
    .I1(_4157_),
    .S(_4154_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8318_ (.A1(_4150_),
    .A2(\registers[29][15] ),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8319_ (.I0(_1133_),
    .I1(_4158_),
    .S(_4154_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8320_ (.A1(_4150_),
    .A2(\registers[29][16] ),
    .Z(_4159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8321_ (.I0(_1135_),
    .I1(_4159_),
    .S(_4154_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8322_ (.A1(_4150_),
    .A2(\registers[29][17] ),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8323_ (.I0(_1137_),
    .I1(_4160_),
    .S(_4154_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8324_ (.A1(_4150_),
    .A2(\registers[29][18] ),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8325_ (.I0(_1139_),
    .I1(_4161_),
    .S(_4154_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _8326_ (.I(_1639_),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8327_ (.A1(_4162_),
    .A2(\registers[29][19] ),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8328_ (.I0(_1142_),
    .I1(_4163_),
    .S(_4154_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8329_ (.A1(_4162_),
    .A2(\registers[29][1] ),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8330_ (.I0(_1145_),
    .I1(_4164_),
    .S(_4154_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8331_ (.A1(_4162_),
    .A2(\registers[29][20] ),
    .Z(_4165_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _8332_ (.I(_1096_),
    .Z(_4166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8333_ (.I0(_1147_),
    .I1(_4165_),
    .S(_4166_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8334_ (.A1(_4162_),
    .A2(\registers[29][21] ),
    .Z(_4167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8335_ (.I0(_1149_),
    .I1(_4167_),
    .S(_4166_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8336_ (.A1(_4162_),
    .A2(\registers[29][22] ),
    .Z(_4168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8337_ (.I0(_1151_),
    .I1(_4168_),
    .S(_4166_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8338_ (.A1(_4162_),
    .A2(\registers[29][23] ),
    .Z(_4169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8339_ (.I0(_1153_),
    .I1(_4169_),
    .S(_4166_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8340_ (.A1(_4162_),
    .A2(\registers[29][24] ),
    .Z(_4170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8341_ (.I0(_1155_),
    .I1(_4170_),
    .S(_4166_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8342_ (.A1(_4162_),
    .A2(\registers[29][25] ),
    .Z(_4171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8343_ (.I0(_1157_),
    .I1(_4171_),
    .S(_4166_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8344_ (.A1(_4162_),
    .A2(\registers[29][26] ),
    .Z(_4172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8345_ (.I0(_1159_),
    .I1(_4172_),
    .S(_4166_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8346_ (.A1(_4162_),
    .A2(\registers[29][27] ),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8347_ (.I0(_1161_),
    .I1(_4173_),
    .S(_4166_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8348_ (.A1(_1112_),
    .A2(\registers[29][28] ),
    .Z(_4174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8349_ (.I0(_1164_),
    .I1(_4174_),
    .S(_4166_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8350_ (.A1(_1112_),
    .A2(\registers[29][29] ),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8351_ (.I0(_1167_),
    .I1(_4175_),
    .S(_4166_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8352_ (.A1(_1112_),
    .A2(\registers[29][2] ),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8353_ (.I0(_1169_),
    .I1(_4176_),
    .S(_1096_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _8354_ (.A1(_1112_),
    .A2(\registers[29][30] ),
    .Z(_4177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _8355_ (.I0(_1171_),
    .I1(_4177_),
    .S(_1096_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[0]$_SDFFCE_PN0P_  (.D(_0329_),
    .CLK(clknet_leaf_28_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[10]$_SDFFCE_PN0P_  (.D(_0330_),
    .CLK(clknet_leaf_28_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[11]$_SDFFCE_PN0P_  (.D(_0331_),
    .CLK(clknet_leaf_24_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[12]$_SDFFCE_PN0P_  (.D(_0332_),
    .CLK(clknet_leaf_24_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[13]$_SDFFCE_PN0P_  (.D(_0333_),
    .CLK(clknet_leaf_24_clk),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[14]$_SDFFCE_PN0P_  (.D(_0334_),
    .CLK(clknet_leaf_25_clk),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[15]$_SDFFCE_PN0P_  (.D(_0335_),
    .CLK(clknet_leaf_20_clk),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[16]$_SDFFCE_PN0P_  (.D(_0336_),
    .CLK(clknet_leaf_19_clk),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[17]$_SDFFCE_PN0P_  (.D(_0337_),
    .CLK(clknet_leaf_19_clk),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[18]$_SDFFCE_PN0P_  (.D(_0338_),
    .CLK(clknet_leaf_20_clk),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[19]$_SDFFCE_PN0P_  (.D(_0339_),
    .CLK(clknet_leaf_18_clk),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[1]$_SDFFCE_PN0P_  (.D(_0340_),
    .CLK(clknet_leaf_18_clk),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[20]$_SDFFCE_PN0P_  (.D(_0341_),
    .CLK(clknet_leaf_12_clk),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[21]$_SDFFCE_PN0P_  (.D(_0342_),
    .CLK(clknet_leaf_12_clk),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[22]$_SDFFCE_PN0P_  (.D(_0343_),
    .CLK(clknet_leaf_10_clk),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[23]$_SDFFCE_PN0P_  (.D(_0344_),
    .CLK(clknet_leaf_10_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[24]$_SDFFCE_PN0P_  (.D(_0345_),
    .CLK(clknet_leaf_8_clk),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[25]$_SDFFCE_PN0P_  (.D(_0346_),
    .CLK(clknet_leaf_8_clk),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[26]$_SDFFCE_PN0P_  (.D(_0347_),
    .CLK(clknet_leaf_7_clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[27]$_SDFFCE_PN0P_  (.D(_0348_),
    .CLK(clknet_leaf_8_clk),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[28]$_SDFFCE_PN0P_  (.D(_0349_),
    .CLK(clknet_leaf_2_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[29]$_SDFFCE_PN0P_  (.D(_0350_),
    .CLK(clknet_leaf_1_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[2]$_SDFFCE_PN0P_  (.D(_0351_),
    .CLK(clknet_leaf_1_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[30]$_SDFFCE_PN0P_  (.D(_0352_),
    .CLK(clknet_leaf_1_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[31]$_SDFFCE_PN0P_  (.D(_0353_),
    .CLK(clknet_leaf_4_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[3]$_SDFFCE_PN0P_  (.D(_0354_),
    .CLK(clknet_leaf_37_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[4]$_SDFFCE_PN0P_  (.D(_0355_),
    .CLK(clknet_leaf_38_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[5]$_SDFFCE_PN0P_  (.D(_0356_),
    .CLK(clknet_leaf_33_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[6]$_SDFFCE_PN0P_  (.D(_0357_),
    .CLK(clknet_leaf_34_clk),
    .Q(net76));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[7]$_SDFFCE_PN0P_  (.D(_0358_),
    .CLK(clknet_leaf_34_clk),
    .Q(net77));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[8]$_SDFFCE_PN0P_  (.D(_0359_),
    .CLK(clknet_leaf_34_clk),
    .Q(net78));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data1[9]$_SDFFCE_PN0P_  (.D(_0360_),
    .CLK(clknet_leaf_34_clk),
    .Q(net79));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[0]$_SDFFCE_PN0P_  (.D(_0361_),
    .CLK(clknet_leaf_28_clk),
    .Q(net80));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[10]$_SDFFCE_PN0P_  (.D(_0362_),
    .CLK(clknet_leaf_28_clk),
    .Q(net81));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[11]$_SDFFCE_PN0P_  (.D(_0363_),
    .CLK(clknet_leaf_24_clk),
    .Q(net82));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[12]$_SDFFCE_PN0P_  (.D(_0364_),
    .CLK(clknet_leaf_28_clk),
    .Q(net83));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[13]$_SDFFCE_PN0P_  (.D(_0365_),
    .CLK(clknet_leaf_24_clk),
    .Q(net84));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[14]$_SDFFCE_PN0P_  (.D(_0366_),
    .CLK(clknet_leaf_25_clk),
    .Q(net85));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[15]$_SDFFCE_PN0P_  (.D(_0367_),
    .CLK(clknet_leaf_17_clk),
    .Q(net86));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[16]$_SDFFCE_PN0P_  (.D(_0368_),
    .CLK(clknet_leaf_20_clk),
    .Q(net87));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[17]$_SDFFCE_PN0P_  (.D(_0369_),
    .CLK(clknet_leaf_20_clk),
    .Q(net88));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[18]$_SDFFCE_PN0P_  (.D(_0370_),
    .CLK(clknet_leaf_20_clk),
    .Q(net89));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[19]$_SDFFCE_PN0P_  (.D(_0371_),
    .CLK(clknet_leaf_18_clk),
    .Q(net90));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[1]$_SDFFCE_PN0P_  (.D(_0372_),
    .CLK(clknet_leaf_17_clk),
    .Q(net91));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[20]$_SDFFCE_PN0P_  (.D(_0373_),
    .CLK(clknet_leaf_13_clk),
    .Q(net92));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[21]$_SDFFCE_PN0P_  (.D(_0374_),
    .CLK(clknet_leaf_14_clk),
    .Q(net93));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[22]$_SDFFCE_PN0P_  (.D(_0375_),
    .CLK(clknet_leaf_9_clk),
    .Q(net94));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[23]$_SDFFCE_PN0P_  (.D(_0376_),
    .CLK(clknet_leaf_11_clk),
    .Q(net95));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[24]$_SDFFCE_PN0P_  (.D(_0377_),
    .CLK(clknet_leaf_9_clk),
    .Q(net96));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[25]$_SDFFCE_PN0P_  (.D(_0378_),
    .CLK(clknet_leaf_9_clk),
    .Q(net97));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[26]$_SDFFCE_PN0P_  (.D(_0379_),
    .CLK(clknet_leaf_8_clk),
    .Q(net98));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[27]$_SDFFCE_PN0P_  (.D(_0380_),
    .CLK(clknet_leaf_8_clk),
    .Q(net99));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[28]$_SDFFCE_PN0P_  (.D(_0381_),
    .CLK(clknet_leaf_1_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[29]$_SDFFCE_PN0P_  (.D(_0382_),
    .CLK(clknet_leaf_1_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[2]$_SDFFCE_PN0P_  (.D(_0383_),
    .CLK(clknet_leaf_3_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[30]$_SDFFCE_PN0P_  (.D(_0384_),
    .CLK(clknet_leaf_1_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[31]$_SDFFCE_PN0P_  (.D(_0385_),
    .CLK(clknet_leaf_4_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[3]$_SDFFCE_PN0P_  (.D(_0386_),
    .CLK(clknet_leaf_37_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[4]$_SDFFCE_PN0P_  (.D(_0387_),
    .CLK(clknet_leaf_36_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[5]$_SDFFCE_PN0P_  (.D(_0388_),
    .CLK(clknet_leaf_38_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[6]$_SDFFCE_PN0P_  (.D(_0389_),
    .CLK(clknet_leaf_36_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[7]$_SDFFCE_PN0P_  (.D(_0390_),
    .CLK(clknet_leaf_33_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[8]$_SDFFCE_PN0P_  (.D(_0391_),
    .CLK(clknet_leaf_34_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \read_data2[9]$_SDFFCE_PN0P_  (.D(_0392_),
    .CLK(clknet_leaf_34_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][0]$_SDFFCE_PN0P_  (.D(_0393_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][10]$_SDFFCE_PN0P_  (.D(_0394_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][11]$_SDFFCE_PN0P_  (.D(_0395_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][12]$_SDFFCE_PN0P_  (.D(_0396_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][13]$_SDFFCE_PN0P_  (.D(_0397_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][14]$_SDFFCE_PN0P_  (.D(_0398_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][15]$_SDFFCE_PN0P_  (.D(_0399_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][16]$_SDFFCE_PN0P_  (.D(_0400_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][17]$_SDFFCE_PN0P_  (.D(_0401_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][18]$_SDFFCE_PN0P_  (.D(_0402_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][19]$_SDFFCE_PN0P_  (.D(_0403_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][1]$_SDFFCE_PN0P_  (.D(_0404_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][20]$_SDFFCE_PN0P_  (.D(_0405_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][21]$_SDFFCE_PN0P_  (.D(_0406_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][22]$_SDFFCE_PN0P_  (.D(_0407_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][23]$_SDFFCE_PN0P_  (.D(_0408_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][24]$_SDFFCE_PN0P_  (.D(_0409_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][25]$_SDFFCE_PN0P_  (.D(_0410_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][26]$_SDFFCE_PN0P_  (.D(_0411_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][27]$_SDFFCE_PN0P_  (.D(_0412_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][28]$_SDFFCE_PN0P_  (.D(_0413_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][29]$_SDFFCE_PN0P_  (.D(_0414_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][2]$_SDFFCE_PN0P_  (.D(_0415_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][30]$_SDFFCE_PN0P_  (.D(_0416_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][31]$_SDFFCE_PN0P_  (.D(_0417_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][3]$_SDFFCE_PN0P_  (.D(_0418_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][4]$_SDFFCE_PN0P_  (.D(_0419_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][5]$_SDFFCE_PN0P_  (.D(_0420_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][6]$_SDFFCE_PN0P_  (.D(_0421_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][7]$_SDFFCE_PN0P_  (.D(_0422_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][8]$_SDFFCE_PN0P_  (.D(_0423_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[0][9]$_SDFFCE_PN0P_  (.D(_0424_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][0]$_SDFFCE_PN0P_  (.D(_0425_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[10][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][10]$_SDFFCE_PN0P_  (.D(_0426_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[10][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][11]$_SDFFCE_PN0P_  (.D(_0427_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[10][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][12]$_SDFFCE_PN0P_  (.D(_0428_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[10][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][13]$_SDFFCE_PN0P_  (.D(_0429_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[10][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][14]$_SDFFCE_PN0P_  (.D(_0430_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[10][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][15]$_SDFFCE_PN0P_  (.D(_0431_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[10][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][16]$_SDFFCE_PN0P_  (.D(_0432_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[10][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][17]$_SDFFCE_PN0P_  (.D(_0433_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[10][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][18]$_SDFFCE_PN0P_  (.D(_0434_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[10][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][19]$_SDFFCE_PN0P_  (.D(_0435_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[10][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][1]$_SDFFCE_PN0P_  (.D(_0436_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[10][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][20]$_SDFFCE_PN0P_  (.D(_0437_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[10][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][21]$_SDFFCE_PN0P_  (.D(_0438_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[10][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][22]$_SDFFCE_PN0P_  (.D(_0439_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[10][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][23]$_SDFFCE_PN0P_  (.D(_0440_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[10][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][24]$_SDFFCE_PN0P_  (.D(_0441_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[10][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][25]$_SDFFCE_PN0P_  (.D(_0442_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[10][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][26]$_SDFFCE_PN0P_  (.D(_0443_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[10][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][27]$_SDFFCE_PN0P_  (.D(_0444_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[10][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][28]$_SDFFCE_PN0P_  (.D(_0445_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[10][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][29]$_SDFFCE_PN0P_  (.D(_0446_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[10][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][2]$_SDFFCE_PN0P_  (.D(_0447_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[10][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][30]$_SDFFCE_PN0P_  (.D(_0448_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[10][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][31]$_SDFFCE_PN0P_  (.D(_0449_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[10][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][3]$_SDFFCE_PN0P_  (.D(_0450_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[10][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][4]$_SDFFCE_PN0P_  (.D(_0451_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[10][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][5]$_SDFFCE_PN0P_  (.D(_0452_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[10][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][6]$_SDFFCE_PN0P_  (.D(_0453_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[10][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][7]$_SDFFCE_PN0P_  (.D(_0454_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[10][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][8]$_SDFFCE_PN0P_  (.D(_0455_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[10][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[10][9]$_SDFFCE_PN0P_  (.D(_0456_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[10][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][0]$_SDFFCE_PN0P_  (.D(_0457_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[11][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][10]$_SDFFCE_PN0P_  (.D(_0458_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[11][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][11]$_SDFFCE_PN0P_  (.D(_0459_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[11][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][12]$_SDFFCE_PN0P_  (.D(_0460_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[11][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][13]$_SDFFCE_PN0P_  (.D(_0461_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[11][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][14]$_SDFFCE_PN0P_  (.D(_0462_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[11][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][15]$_SDFFCE_PN0P_  (.D(_0463_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[11][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][16]$_SDFFCE_PN0P_  (.D(_0464_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[11][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][17]$_SDFFCE_PN0P_  (.D(_0465_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[11][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][18]$_SDFFCE_PN0P_  (.D(_0466_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[11][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][19]$_SDFFCE_PN0P_  (.D(_0467_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[11][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][1]$_SDFFCE_PN0P_  (.D(_0468_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[11][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][20]$_SDFFCE_PN0P_  (.D(_0469_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[11][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][21]$_SDFFCE_PN0P_  (.D(_0470_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[11][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][22]$_SDFFCE_PN0P_  (.D(_0471_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[11][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][23]$_SDFFCE_PN0P_  (.D(_0472_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[11][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][24]$_SDFFCE_PN0P_  (.D(_0473_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[11][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][25]$_SDFFCE_PN0P_  (.D(_0474_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[11][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][26]$_SDFFCE_PN0P_  (.D(_0475_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[11][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][27]$_SDFFCE_PN0P_  (.D(_0476_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[11][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][28]$_SDFFCE_PN0P_  (.D(_0477_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[11][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][29]$_SDFFCE_PN0P_  (.D(_0478_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[11][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][2]$_SDFFCE_PN0P_  (.D(_0479_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[11][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][30]$_SDFFCE_PN0P_  (.D(_0480_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[11][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][31]$_SDFFCE_PN0P_  (.D(_0481_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[11][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][3]$_SDFFCE_PN0P_  (.D(_0482_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[11][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][4]$_SDFFCE_PN0P_  (.D(_0483_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[11][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][5]$_SDFFCE_PN0P_  (.D(_0484_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[11][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][6]$_SDFFCE_PN0P_  (.D(_0485_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[11][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][7]$_SDFFCE_PN0P_  (.D(_0486_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[11][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][8]$_SDFFCE_PN0P_  (.D(_0487_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[11][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[11][9]$_SDFFCE_PN0P_  (.D(_0488_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[11][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][0]$_SDFFCE_PN0P_  (.D(_0489_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[12][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][10]$_SDFFCE_PN0P_  (.D(_0490_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[12][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][11]$_SDFFCE_PN0P_  (.D(_0491_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[12][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][12]$_SDFFCE_PN0P_  (.D(_0492_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[12][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][13]$_SDFFCE_PN0P_  (.D(_0493_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[12][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][14]$_SDFFCE_PN0P_  (.D(_0494_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[12][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][15]$_SDFFCE_PN0P_  (.D(_0495_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[12][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][16]$_SDFFCE_PN0P_  (.D(_0496_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[12][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][17]$_SDFFCE_PN0P_  (.D(_0497_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[12][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][18]$_SDFFCE_PN0P_  (.D(_0498_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[12][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][19]$_SDFFCE_PN0P_  (.D(_0499_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[12][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][1]$_SDFFCE_PN0P_  (.D(_0500_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[12][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][20]$_SDFFCE_PN0P_  (.D(_0501_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[12][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][21]$_SDFFCE_PN0P_  (.D(_0502_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[12][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][22]$_SDFFCE_PN0P_  (.D(_0503_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[12][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][23]$_SDFFCE_PN0P_  (.D(_0504_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[12][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][24]$_SDFFCE_PN0P_  (.D(_0505_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[12][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][25]$_SDFFCE_PN0P_  (.D(_0506_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[12][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][26]$_SDFFCE_PN0P_  (.D(_0507_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[12][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][27]$_SDFFCE_PN0P_  (.D(_0508_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[12][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][28]$_SDFFCE_PN0P_  (.D(_0509_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[12][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][29]$_SDFFCE_PN0P_  (.D(_0510_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[12][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][2]$_SDFFCE_PN0P_  (.D(_0511_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[12][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][30]$_SDFFCE_PN0P_  (.D(_0512_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[12][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][31]$_SDFFCE_PN0P_  (.D(_0513_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[12][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][3]$_SDFFCE_PN0P_  (.D(_0514_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[12][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][4]$_SDFFCE_PN0P_  (.D(_0515_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[12][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][5]$_SDFFCE_PN0P_  (.D(_0516_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[12][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][6]$_SDFFCE_PN0P_  (.D(_0517_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[12][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][7]$_SDFFCE_PN0P_  (.D(_0518_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[12][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][8]$_SDFFCE_PN0P_  (.D(_0519_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[12][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[12][9]$_SDFFCE_PN0P_  (.D(_0520_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[12][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][0]$_SDFFCE_PN0P_  (.D(_0521_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[13][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][10]$_SDFFCE_PN0P_  (.D(_0522_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[13][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][11]$_SDFFCE_PN0P_  (.D(_0523_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[13][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][12]$_SDFFCE_PN0P_  (.D(_0524_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[13][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][13]$_SDFFCE_PN0P_  (.D(_0525_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[13][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][14]$_SDFFCE_PN0P_  (.D(_0526_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[13][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][15]$_SDFFCE_PN0P_  (.D(_0527_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[13][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][16]$_SDFFCE_PN0P_  (.D(_0528_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[13][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][17]$_SDFFCE_PN0P_  (.D(_0529_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[13][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][18]$_SDFFCE_PN0P_  (.D(_0530_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[13][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][19]$_SDFFCE_PN0P_  (.D(_0531_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[13][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][1]$_SDFFCE_PN0P_  (.D(_0532_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[13][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][20]$_SDFFCE_PN0P_  (.D(_0533_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[13][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][21]$_SDFFCE_PN0P_  (.D(_0534_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[13][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][22]$_SDFFCE_PN0P_  (.D(_0535_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[13][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][23]$_SDFFCE_PN0P_  (.D(_0536_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[13][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][24]$_SDFFCE_PN0P_  (.D(_0537_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[13][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][25]$_SDFFCE_PN0P_  (.D(_0538_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[13][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][26]$_SDFFCE_PN0P_  (.D(_0539_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[13][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][27]$_SDFFCE_PN0P_  (.D(_0540_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[13][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][28]$_SDFFCE_PN0P_  (.D(_0541_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[13][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][29]$_SDFFCE_PN0P_  (.D(_0542_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[13][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][2]$_SDFFCE_PN0P_  (.D(_0543_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[13][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][30]$_SDFFCE_PN0P_  (.D(_0544_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[13][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][31]$_SDFFCE_PN0P_  (.D(_0545_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[13][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][3]$_SDFFCE_PN0P_  (.D(_0546_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[13][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][4]$_SDFFCE_PN0P_  (.D(_0547_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[13][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][5]$_SDFFCE_PN0P_  (.D(_0548_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[13][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][6]$_SDFFCE_PN0P_  (.D(_0549_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[13][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][7]$_SDFFCE_PN0P_  (.D(_0550_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[13][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][8]$_SDFFCE_PN0P_  (.D(_0551_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[13][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[13][9]$_SDFFCE_PN0P_  (.D(_0552_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[13][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][0]$_SDFFCE_PN0P_  (.D(_0553_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[14][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][10]$_SDFFCE_PN0P_  (.D(_0554_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[14][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][11]$_SDFFCE_PN0P_  (.D(_0555_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[14][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][12]$_SDFFCE_PN0P_  (.D(_0556_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[14][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][13]$_SDFFCE_PN0P_  (.D(_0557_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[14][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][14]$_SDFFCE_PN0P_  (.D(_0558_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[14][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][15]$_SDFFCE_PN0P_  (.D(_0559_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[14][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][16]$_SDFFCE_PN0P_  (.D(_0560_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[14][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][17]$_SDFFCE_PN0P_  (.D(_0561_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[14][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][18]$_SDFFCE_PN0P_  (.D(_0562_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[14][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][19]$_SDFFCE_PN0P_  (.D(_0563_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[14][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][1]$_SDFFCE_PN0P_  (.D(_0564_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[14][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][20]$_SDFFCE_PN0P_  (.D(_0565_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[14][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][21]$_SDFFCE_PN0P_  (.D(_0566_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[14][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][22]$_SDFFCE_PN0P_  (.D(_0567_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[14][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][23]$_SDFFCE_PN0P_  (.D(_0568_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[14][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][24]$_SDFFCE_PN0P_  (.D(_0569_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[14][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][25]$_SDFFCE_PN0P_  (.D(_0570_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[14][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][26]$_SDFFCE_PN0P_  (.D(_0571_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[14][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][27]$_SDFFCE_PN0P_  (.D(_0572_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[14][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][28]$_SDFFCE_PN0P_  (.D(_0573_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[14][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][29]$_SDFFCE_PN0P_  (.D(_0574_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[14][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][2]$_SDFFCE_PN0P_  (.D(_0575_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[14][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][30]$_SDFFCE_PN0P_  (.D(_0576_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[14][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][31]$_SDFFCE_PN0P_  (.D(_0577_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[14][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][3]$_SDFFCE_PN0P_  (.D(_0578_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[14][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][4]$_SDFFCE_PN0P_  (.D(_0579_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[14][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][5]$_SDFFCE_PN0P_  (.D(_0580_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[14][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][6]$_SDFFCE_PN0P_  (.D(_0581_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[14][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][7]$_SDFFCE_PN0P_  (.D(_0582_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[14][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][8]$_SDFFCE_PN0P_  (.D(_0583_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[14][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[14][9]$_SDFFCE_PN0P_  (.D(_0584_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[14][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][0]$_SDFFCE_PN0P_  (.D(_0585_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[15][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][10]$_SDFFCE_PN0P_  (.D(_0586_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[15][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][11]$_SDFFCE_PN0P_  (.D(_0587_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[15][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][12]$_SDFFCE_PN0P_  (.D(_0588_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[15][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][13]$_SDFFCE_PN0P_  (.D(_0589_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[15][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][14]$_SDFFCE_PN0P_  (.D(_0590_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[15][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][15]$_SDFFCE_PN0P_  (.D(_0591_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[15][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][16]$_SDFFCE_PN0P_  (.D(_0592_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[15][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][17]$_SDFFCE_PN0P_  (.D(_0593_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[15][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][18]$_SDFFCE_PN0P_  (.D(_0594_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[15][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][19]$_SDFFCE_PN0P_  (.D(_0595_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[15][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][1]$_SDFFCE_PN0P_  (.D(_0596_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[15][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][20]$_SDFFCE_PN0P_  (.D(_0597_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[15][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][21]$_SDFFCE_PN0P_  (.D(_0598_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[15][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][22]$_SDFFCE_PN0P_  (.D(_0599_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[15][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][23]$_SDFFCE_PN0P_  (.D(_0600_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[15][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][24]$_SDFFCE_PN0P_  (.D(_0601_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[15][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][25]$_SDFFCE_PN0P_  (.D(_0602_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[15][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][26]$_SDFFCE_PN0P_  (.D(_0603_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[15][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][27]$_SDFFCE_PN0P_  (.D(_0604_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[15][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][28]$_SDFFCE_PN0P_  (.D(_0605_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[15][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][29]$_SDFFCE_PN0P_  (.D(_0606_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[15][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][2]$_SDFFCE_PN0P_  (.D(_0607_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[15][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][30]$_SDFFCE_PN0P_  (.D(_0608_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[15][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][31]$_SDFFCE_PN0P_  (.D(_0609_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[15][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][3]$_SDFFCE_PN0P_  (.D(_0610_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[15][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][4]$_SDFFCE_PN0P_  (.D(_0611_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[15][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][5]$_SDFFCE_PN0P_  (.D(_0612_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[15][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][6]$_SDFFCE_PN0P_  (.D(_0613_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[15][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][7]$_SDFFCE_PN0P_  (.D(_0614_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[15][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][8]$_SDFFCE_PN0P_  (.D(_0615_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[15][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[15][9]$_SDFFCE_PN0P_  (.D(_0616_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[15][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][0]$_SDFFCE_PN0P_  (.D(_0617_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[16][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][10]$_SDFFCE_PN0P_  (.D(_0618_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[16][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][11]$_SDFFCE_PN0P_  (.D(_0619_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[16][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][12]$_SDFFCE_PN0P_  (.D(_0620_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[16][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][13]$_SDFFCE_PN0P_  (.D(_0621_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[16][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][14]$_SDFFCE_PN0P_  (.D(_0622_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[16][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][15]$_SDFFCE_PN0P_  (.D(_0623_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[16][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][16]$_SDFFCE_PN0P_  (.D(_0624_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[16][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][17]$_SDFFCE_PN0P_  (.D(_0625_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[16][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][18]$_SDFFCE_PN0P_  (.D(_0626_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[16][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][19]$_SDFFCE_PN0P_  (.D(_0627_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[16][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][1]$_SDFFCE_PN0P_  (.D(_0628_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[16][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][20]$_SDFFCE_PN0P_  (.D(_0629_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[16][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][21]$_SDFFCE_PN0P_  (.D(_0630_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[16][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][22]$_SDFFCE_PN0P_  (.D(_0631_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[16][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][23]$_SDFFCE_PN0P_  (.D(_0632_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[16][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][24]$_SDFFCE_PN0P_  (.D(_0633_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[16][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][25]$_SDFFCE_PN0P_  (.D(_0634_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[16][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][26]$_SDFFCE_PN0P_  (.D(_0635_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[16][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][27]$_SDFFCE_PN0P_  (.D(_0636_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[16][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][28]$_SDFFCE_PN0P_  (.D(_0637_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[16][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][29]$_SDFFCE_PN0P_  (.D(_0638_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[16][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][2]$_SDFFCE_PN0P_  (.D(_0639_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[16][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][30]$_SDFFCE_PN0P_  (.D(_0640_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[16][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][31]$_SDFFCE_PN0P_  (.D(_0641_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[16][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][3]$_SDFFCE_PN0P_  (.D(_0642_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[16][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][4]$_SDFFCE_PN0P_  (.D(_0643_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[16][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][5]$_SDFFCE_PN0P_  (.D(_0644_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[16][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][6]$_SDFFCE_PN0P_  (.D(_0645_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[16][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][7]$_SDFFCE_PN0P_  (.D(_0646_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[16][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][8]$_SDFFCE_PN0P_  (.D(_0647_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[16][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[16][9]$_SDFFCE_PN0P_  (.D(_0648_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[16][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][0]$_SDFFCE_PN0P_  (.D(_0649_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[17][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][10]$_SDFFCE_PN0P_  (.D(_0650_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[17][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][11]$_SDFFCE_PN0P_  (.D(_0651_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[17][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][12]$_SDFFCE_PN0P_  (.D(_0652_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[17][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][13]$_SDFFCE_PN0P_  (.D(_0653_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[17][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][14]$_SDFFCE_PN0P_  (.D(_0654_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[17][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][15]$_SDFFCE_PN0P_  (.D(_0655_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[17][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][16]$_SDFFCE_PN0P_  (.D(_0656_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[17][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][17]$_SDFFCE_PN0P_  (.D(_0657_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[17][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][18]$_SDFFCE_PN0P_  (.D(_0658_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[17][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][19]$_SDFFCE_PN0P_  (.D(_0659_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[17][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][1]$_SDFFCE_PN0P_  (.D(_0660_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[17][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][20]$_SDFFCE_PN0P_  (.D(_0661_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[17][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][21]$_SDFFCE_PN0P_  (.D(_0662_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[17][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][22]$_SDFFCE_PN0P_  (.D(_0663_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[17][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][23]$_SDFFCE_PN0P_  (.D(_0664_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[17][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][24]$_SDFFCE_PN0P_  (.D(_0665_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[17][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][25]$_SDFFCE_PN0P_  (.D(_0666_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[17][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][26]$_SDFFCE_PN0P_  (.D(_0667_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[17][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][27]$_SDFFCE_PN0P_  (.D(_0668_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[17][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][28]$_SDFFCE_PN0P_  (.D(_0669_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[17][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][29]$_SDFFCE_PN0P_  (.D(_0670_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[17][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][2]$_SDFFCE_PN0P_  (.D(_0671_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[17][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][30]$_SDFFCE_PN0P_  (.D(_0672_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[17][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][31]$_SDFFCE_PN0P_  (.D(_0673_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[17][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][3]$_SDFFCE_PN0P_  (.D(_0674_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[17][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][4]$_SDFFCE_PN0P_  (.D(_0675_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[17][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][5]$_SDFFCE_PN0P_  (.D(_0676_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[17][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][6]$_SDFFCE_PN0P_  (.D(_0677_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[17][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][7]$_SDFFCE_PN0P_  (.D(_0678_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[17][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][8]$_SDFFCE_PN0P_  (.D(_0679_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[17][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[17][9]$_SDFFCE_PN0P_  (.D(_0680_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[17][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][0]$_SDFFCE_PN0P_  (.D(_0681_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[18][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][10]$_SDFFCE_PN0P_  (.D(_0682_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[18][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][11]$_SDFFCE_PN0P_  (.D(_0683_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[18][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][12]$_SDFFCE_PN0P_  (.D(_0684_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[18][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][13]$_SDFFCE_PN0P_  (.D(_0685_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[18][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][14]$_SDFFCE_PN0P_  (.D(_0686_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[18][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][15]$_SDFFCE_PN0P_  (.D(_0687_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[18][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][16]$_SDFFCE_PN0P_  (.D(_0688_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[18][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][17]$_SDFFCE_PN0P_  (.D(_0689_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[18][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][18]$_SDFFCE_PN0P_  (.D(_0690_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[18][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][19]$_SDFFCE_PN0P_  (.D(_0691_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[18][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][1]$_SDFFCE_PN0P_  (.D(_0692_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[18][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][20]$_SDFFCE_PN0P_  (.D(_0693_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[18][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][21]$_SDFFCE_PN0P_  (.D(_0694_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[18][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][22]$_SDFFCE_PN0P_  (.D(_0695_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[18][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][23]$_SDFFCE_PN0P_  (.D(_0696_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[18][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][24]$_SDFFCE_PN0P_  (.D(_0697_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[18][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][25]$_SDFFCE_PN0P_  (.D(_0698_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[18][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][26]$_SDFFCE_PN0P_  (.D(_0699_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[18][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][27]$_SDFFCE_PN0P_  (.D(_0700_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[18][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][28]$_SDFFCE_PN0P_  (.D(_0701_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[18][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][29]$_SDFFCE_PN0P_  (.D(_0702_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[18][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][2]$_SDFFCE_PN0P_  (.D(_0703_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[18][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][30]$_SDFFCE_PN0P_  (.D(_0704_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[18][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][31]$_SDFFCE_PN0P_  (.D(_0705_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[18][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][3]$_SDFFCE_PN0P_  (.D(_0706_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[18][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][4]$_SDFFCE_PN0P_  (.D(_0707_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[18][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][5]$_SDFFCE_PN0P_  (.D(_0708_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[18][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][6]$_SDFFCE_PN0P_  (.D(_0709_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[18][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][7]$_SDFFCE_PN0P_  (.D(_0710_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[18][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][8]$_SDFFCE_PN0P_  (.D(_0711_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[18][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[18][9]$_SDFFCE_PN0P_  (.D(_0712_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[18][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][0]$_SDFFCE_PN0P_  (.D(_0713_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[19][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][10]$_SDFFCE_PN0P_  (.D(_0714_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[19][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][11]$_SDFFCE_PN0P_  (.D(_0715_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[19][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][12]$_SDFFCE_PN0P_  (.D(_0716_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[19][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][13]$_SDFFCE_PN0P_  (.D(_0717_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[19][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][14]$_SDFFCE_PN0P_  (.D(_0718_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[19][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][15]$_SDFFCE_PN0P_  (.D(_0719_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[19][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][16]$_SDFFCE_PN0P_  (.D(_0720_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[19][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][17]$_SDFFCE_PN0P_  (.D(_0721_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[19][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][18]$_SDFFCE_PN0P_  (.D(_0722_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[19][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][19]$_SDFFCE_PN0P_  (.D(_0723_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[19][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][1]$_SDFFCE_PN0P_  (.D(_0724_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[19][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][20]$_SDFFCE_PN0P_  (.D(_0725_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[19][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][21]$_SDFFCE_PN0P_  (.D(_0726_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[19][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][22]$_SDFFCE_PN0P_  (.D(_0727_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[19][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][23]$_SDFFCE_PN0P_  (.D(_0728_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[19][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][24]$_SDFFCE_PN0P_  (.D(_0729_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[19][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][25]$_SDFFCE_PN0P_  (.D(_0730_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[19][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][26]$_SDFFCE_PN0P_  (.D(_0731_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[19][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][27]$_SDFFCE_PN0P_  (.D(_0732_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[19][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][28]$_SDFFCE_PN0P_  (.D(_0733_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[19][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][29]$_SDFFCE_PN0P_  (.D(_0734_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[19][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][2]$_SDFFCE_PN0P_  (.D(_0735_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[19][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][30]$_SDFFCE_PN0P_  (.D(_0736_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[19][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][31]$_SDFFCE_PN0P_  (.D(_0737_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[19][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][3]$_SDFFCE_PN0P_  (.D(_0738_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[19][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][4]$_SDFFCE_PN0P_  (.D(_0739_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[19][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][5]$_SDFFCE_PN0P_  (.D(_0740_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[19][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][6]$_SDFFCE_PN0P_  (.D(_0741_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[19][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][7]$_SDFFCE_PN0P_  (.D(_0742_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[19][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][8]$_SDFFCE_PN0P_  (.D(_0743_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[19][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[19][9]$_SDFFCE_PN0P_  (.D(_0744_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[19][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][0]$_SDFFCE_PN0P_  (.D(_0745_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][10]$_SDFFCE_PN0P_  (.D(_0746_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][11]$_SDFFCE_PN0P_  (.D(_0747_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][12]$_SDFFCE_PN0P_  (.D(_0748_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][13]$_SDFFCE_PN0P_  (.D(_0749_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][14]$_SDFFCE_PN0P_  (.D(_0750_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][15]$_SDFFCE_PN0P_  (.D(_0751_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][16]$_SDFFCE_PN0P_  (.D(_0752_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][17]$_SDFFCE_PN0P_  (.D(_0753_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][18]$_SDFFCE_PN0P_  (.D(_0754_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][19]$_SDFFCE_PN0P_  (.D(_0755_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][1]$_SDFFCE_PN0P_  (.D(_0756_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][20]$_SDFFCE_PN0P_  (.D(_0757_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][21]$_SDFFCE_PN0P_  (.D(_0758_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][22]$_SDFFCE_PN0P_  (.D(_0759_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][23]$_SDFFCE_PN0P_  (.D(_0760_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][24]$_SDFFCE_PN0P_  (.D(_0761_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][25]$_SDFFCE_PN0P_  (.D(_0762_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][26]$_SDFFCE_PN0P_  (.D(_0763_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][27]$_SDFFCE_PN0P_  (.D(_0764_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][28]$_SDFFCE_PN0P_  (.D(_0765_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][29]$_SDFFCE_PN0P_  (.D(_0766_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][2]$_SDFFCE_PN0P_  (.D(_0767_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][30]$_SDFFCE_PN0P_  (.D(_0768_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][31]$_SDFFCE_PN0P_  (.D(_0769_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][3]$_SDFFCE_PN0P_  (.D(_0770_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][4]$_SDFFCE_PN0P_  (.D(_0771_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][5]$_SDFFCE_PN0P_  (.D(_0772_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][6]$_SDFFCE_PN0P_  (.D(_0773_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][7]$_SDFFCE_PN0P_  (.D(_0774_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][8]$_SDFFCE_PN0P_  (.D(_0775_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[1][9]$_SDFFCE_PN0P_  (.D(_0776_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][0]$_SDFFCE_PN0P_  (.D(_0777_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[20][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][10]$_SDFFCE_PN0P_  (.D(_0778_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[20][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][11]$_SDFFCE_PN0P_  (.D(_0779_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[20][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][12]$_SDFFCE_PN0P_  (.D(_0780_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[20][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][13]$_SDFFCE_PN0P_  (.D(_0781_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[20][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][14]$_SDFFCE_PN0P_  (.D(_0782_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[20][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][15]$_SDFFCE_PN0P_  (.D(_0783_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[20][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][16]$_SDFFCE_PN0P_  (.D(_0784_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[20][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][17]$_SDFFCE_PN0P_  (.D(_0785_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[20][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][18]$_SDFFCE_PN0P_  (.D(_0786_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[20][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][19]$_SDFFCE_PN0P_  (.D(_0787_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[20][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][1]$_SDFFCE_PN0P_  (.D(_0788_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[20][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][20]$_SDFFCE_PN0P_  (.D(_0789_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[20][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][21]$_SDFFCE_PN0P_  (.D(_0790_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[20][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][22]$_SDFFCE_PN0P_  (.D(_0791_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[20][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][23]$_SDFFCE_PN0P_  (.D(_0792_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[20][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][24]$_SDFFCE_PN0P_  (.D(_0793_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[20][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][25]$_SDFFCE_PN0P_  (.D(_0794_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[20][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][26]$_SDFFCE_PN0P_  (.D(_0795_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[20][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][27]$_SDFFCE_PN0P_  (.D(_0796_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[20][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][28]$_SDFFCE_PN0P_  (.D(_0797_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[20][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][29]$_SDFFCE_PN0P_  (.D(_0798_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[20][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][2]$_SDFFCE_PN0P_  (.D(_0799_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[20][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][30]$_SDFFCE_PN0P_  (.D(_0800_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[20][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][31]$_SDFFCE_PN0P_  (.D(_0801_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[20][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][3]$_SDFFCE_PN0P_  (.D(_0802_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[20][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][4]$_SDFFCE_PN0P_  (.D(_0803_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[20][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][5]$_SDFFCE_PN0P_  (.D(_0804_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[20][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][6]$_SDFFCE_PN0P_  (.D(_0805_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[20][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][7]$_SDFFCE_PN0P_  (.D(_0806_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[20][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][8]$_SDFFCE_PN0P_  (.D(_0807_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[20][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[20][9]$_SDFFCE_PN0P_  (.D(_0808_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[20][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][0]$_SDFFCE_PN0P_  (.D(_0809_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[21][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][10]$_SDFFCE_PN0P_  (.D(_0810_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[21][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][11]$_SDFFCE_PN0P_  (.D(_0811_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[21][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][12]$_SDFFCE_PN0P_  (.D(_0812_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[21][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][13]$_SDFFCE_PN0P_  (.D(_0813_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[21][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][14]$_SDFFCE_PN0P_  (.D(_0814_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[21][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][15]$_SDFFCE_PN0P_  (.D(_0815_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[21][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][16]$_SDFFCE_PN0P_  (.D(_0816_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[21][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][17]$_SDFFCE_PN0P_  (.D(_0817_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[21][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][18]$_SDFFCE_PN0P_  (.D(_0818_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[21][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][19]$_SDFFCE_PN0P_  (.D(_0819_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[21][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][1]$_SDFFCE_PN0P_  (.D(_0820_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[21][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][20]$_SDFFCE_PN0P_  (.D(_0821_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[21][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][21]$_SDFFCE_PN0P_  (.D(_0822_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[21][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][22]$_SDFFCE_PN0P_  (.D(_0823_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[21][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][23]$_SDFFCE_PN0P_  (.D(_0824_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[21][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][24]$_SDFFCE_PN0P_  (.D(_0825_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[21][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][25]$_SDFFCE_PN0P_  (.D(_0826_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[21][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][26]$_SDFFCE_PN0P_  (.D(_0827_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[21][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][27]$_SDFFCE_PN0P_  (.D(_0828_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[21][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][28]$_SDFFCE_PN0P_  (.D(_0829_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[21][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][29]$_SDFFCE_PN0P_  (.D(_0830_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[21][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][2]$_SDFFCE_PN0P_  (.D(_0831_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[21][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][30]$_SDFFCE_PN0P_  (.D(_0832_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[21][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][31]$_SDFFCE_PN0P_  (.D(_0833_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[21][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][3]$_SDFFCE_PN0P_  (.D(_0834_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[21][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][4]$_SDFFCE_PN0P_  (.D(_0835_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[21][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][5]$_SDFFCE_PN0P_  (.D(_0836_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[21][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][6]$_SDFFCE_PN0P_  (.D(_0837_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[21][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][7]$_SDFFCE_PN0P_  (.D(_0838_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[21][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][8]$_SDFFCE_PN0P_  (.D(_0839_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[21][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[21][9]$_SDFFCE_PN0P_  (.D(_0840_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[21][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][0]$_SDFFCE_PN0P_  (.D(_0841_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[22][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][10]$_SDFFCE_PN0P_  (.D(_0842_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[22][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][11]$_SDFFCE_PN0P_  (.D(_0843_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[22][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][12]$_SDFFCE_PN0P_  (.D(_0844_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[22][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][13]$_SDFFCE_PN0P_  (.D(_0845_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[22][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][14]$_SDFFCE_PN0P_  (.D(_0846_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[22][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][15]$_SDFFCE_PN0P_  (.D(_0847_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[22][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][16]$_SDFFCE_PN0P_  (.D(_0848_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[22][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][17]$_SDFFCE_PN0P_  (.D(_0849_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[22][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][18]$_SDFFCE_PN0P_  (.D(_0850_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[22][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][19]$_SDFFCE_PN0P_  (.D(_0851_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[22][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][1]$_SDFFCE_PN0P_  (.D(_0852_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[22][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][20]$_SDFFCE_PN0P_  (.D(_0853_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[22][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][21]$_SDFFCE_PN0P_  (.D(_0854_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[22][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][22]$_SDFFCE_PN0P_  (.D(_0855_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[22][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][23]$_SDFFCE_PN0P_  (.D(_0856_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[22][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][24]$_SDFFCE_PN0P_  (.D(_0857_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[22][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][25]$_SDFFCE_PN0P_  (.D(_0858_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[22][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][26]$_SDFFCE_PN0P_  (.D(_0859_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[22][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][27]$_SDFFCE_PN0P_  (.D(_0860_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[22][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][28]$_SDFFCE_PN0P_  (.D(_0861_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[22][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][29]$_SDFFCE_PN0P_  (.D(_0862_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[22][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][2]$_SDFFCE_PN0P_  (.D(_0863_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[22][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][30]$_SDFFCE_PN0P_  (.D(_0864_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[22][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][31]$_SDFFCE_PN0P_  (.D(_0865_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[22][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][3]$_SDFFCE_PN0P_  (.D(_0866_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[22][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][4]$_SDFFCE_PN0P_  (.D(_0867_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[22][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][5]$_SDFFCE_PN0P_  (.D(_0868_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[22][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][6]$_SDFFCE_PN0P_  (.D(_0869_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[22][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][7]$_SDFFCE_PN0P_  (.D(_0870_),
    .CLK(clknet_leaf_34_clk),
    .Q(\registers[22][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][8]$_SDFFCE_PN0P_  (.D(_0871_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[22][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[22][9]$_SDFFCE_PN0P_  (.D(_0872_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[22][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][0]$_SDFFCE_PN0P_  (.D(_0873_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[23][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][10]$_SDFFCE_PN0P_  (.D(_0874_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[23][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][11]$_SDFFCE_PN0P_  (.D(_0875_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[23][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][12]$_SDFFCE_PN0P_  (.D(_0876_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[23][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][13]$_SDFFCE_PN0P_  (.D(_0877_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[23][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][14]$_SDFFCE_PN0P_  (.D(_0878_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[23][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][15]$_SDFFCE_PN0P_  (.D(_0879_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[23][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][16]$_SDFFCE_PN0P_  (.D(_0880_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[23][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][17]$_SDFFCE_PN0P_  (.D(_0881_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[23][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][18]$_SDFFCE_PN0P_  (.D(_0882_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[23][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][19]$_SDFFCE_PN0P_  (.D(_0883_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[23][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][1]$_SDFFCE_PN0P_  (.D(_0884_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[23][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][20]$_SDFFCE_PN0P_  (.D(_0885_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[23][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][21]$_SDFFCE_PN0P_  (.D(_0886_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[23][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][22]$_SDFFCE_PN0P_  (.D(_0887_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[23][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][23]$_SDFFCE_PN0P_  (.D(_0888_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[23][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][24]$_SDFFCE_PN0P_  (.D(_0889_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[23][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][25]$_SDFFCE_PN0P_  (.D(_0890_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[23][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][26]$_SDFFCE_PN0P_  (.D(_0891_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[23][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][27]$_SDFFCE_PN0P_  (.D(_0892_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[23][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][28]$_SDFFCE_PN0P_  (.D(_0893_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[23][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][29]$_SDFFCE_PN0P_  (.D(_0894_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[23][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][2]$_SDFFCE_PN0P_  (.D(_0895_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[23][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][30]$_SDFFCE_PN0P_  (.D(_0896_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[23][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][31]$_SDFFCE_PN0P_  (.D(_0897_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[23][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][3]$_SDFFCE_PN0P_  (.D(_0898_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[23][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][4]$_SDFFCE_PN0P_  (.D(_0899_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[23][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][5]$_SDFFCE_PN0P_  (.D(_0900_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[23][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][6]$_SDFFCE_PN0P_  (.D(_0901_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[23][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][7]$_SDFFCE_PN0P_  (.D(_0902_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[23][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][8]$_SDFFCE_PN0P_  (.D(_0903_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[23][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[23][9]$_SDFFCE_PN0P_  (.D(_0904_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[23][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][0]$_SDFFCE_PN0P_  (.D(_0905_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[24][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][10]$_SDFFCE_PN0P_  (.D(_0906_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[24][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][11]$_SDFFCE_PN0P_  (.D(_0907_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[24][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][12]$_SDFFCE_PN0P_  (.D(_0908_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[24][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][13]$_SDFFCE_PN0P_  (.D(_0909_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[24][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][14]$_SDFFCE_PN0P_  (.D(_0910_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[24][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][15]$_SDFFCE_PN0P_  (.D(_0911_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[24][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][16]$_SDFFCE_PN0P_  (.D(_0912_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[24][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][17]$_SDFFCE_PN0P_  (.D(_0913_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[24][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][18]$_SDFFCE_PN0P_  (.D(_0914_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[24][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][19]$_SDFFCE_PN0P_  (.D(_0915_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[24][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][1]$_SDFFCE_PN0P_  (.D(_0916_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[24][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][20]$_SDFFCE_PN0P_  (.D(_0917_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[24][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][21]$_SDFFCE_PN0P_  (.D(_0918_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[24][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][22]$_SDFFCE_PN0P_  (.D(_0919_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[24][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][23]$_SDFFCE_PN0P_  (.D(_0920_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[24][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][24]$_SDFFCE_PN0P_  (.D(_0921_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[24][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][25]$_SDFFCE_PN0P_  (.D(_0922_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[24][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][26]$_SDFFCE_PN0P_  (.D(_0923_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[24][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][27]$_SDFFCE_PN0P_  (.D(_0924_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[24][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][28]$_SDFFCE_PN0P_  (.D(_0925_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[24][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][29]$_SDFFCE_PN0P_  (.D(_0926_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[24][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][2]$_SDFFCE_PN0P_  (.D(_0927_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[24][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][30]$_SDFFCE_PN0P_  (.D(_0928_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[24][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][31]$_SDFFCE_PN0P_  (.D(_0929_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[24][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][3]$_SDFFCE_PN0P_  (.D(_0930_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[24][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][4]$_SDFFCE_PN0P_  (.D(_0931_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[24][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][5]$_SDFFCE_PN0P_  (.D(_0932_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[24][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][6]$_SDFFCE_PN0P_  (.D(_0933_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[24][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][7]$_SDFFCE_PN0P_  (.D(_0934_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[24][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][8]$_SDFFCE_PN0P_  (.D(_0935_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[24][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[24][9]$_SDFFCE_PN0P_  (.D(_0936_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[24][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][0]$_SDFFCE_PN0P_  (.D(_0937_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[25][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][10]$_SDFFCE_PN0P_  (.D(_0938_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[25][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][11]$_SDFFCE_PN0P_  (.D(_0939_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[25][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][12]$_SDFFCE_PN0P_  (.D(_0940_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[25][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][13]$_SDFFCE_PN0P_  (.D(_0941_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[25][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][14]$_SDFFCE_PN0P_  (.D(_0942_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[25][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][15]$_SDFFCE_PN0P_  (.D(_0943_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[25][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][16]$_SDFFCE_PN0P_  (.D(_0944_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[25][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][17]$_SDFFCE_PN0P_  (.D(_0945_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[25][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][18]$_SDFFCE_PN0P_  (.D(_0946_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[25][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][19]$_SDFFCE_PN0P_  (.D(_0947_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[25][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][1]$_SDFFCE_PN0P_  (.D(_0948_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[25][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][20]$_SDFFCE_PN0P_  (.D(_0949_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[25][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][21]$_SDFFCE_PN0P_  (.D(_0950_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[25][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][22]$_SDFFCE_PN0P_  (.D(_0951_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[25][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][23]$_SDFFCE_PN0P_  (.D(_0952_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[25][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][24]$_SDFFCE_PN0P_  (.D(_0953_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[25][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][25]$_SDFFCE_PN0P_  (.D(_0954_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[25][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][26]$_SDFFCE_PN0P_  (.D(_0955_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[25][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][27]$_SDFFCE_PN0P_  (.D(_0956_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[25][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][28]$_SDFFCE_PN0P_  (.D(_0957_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[25][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][29]$_SDFFCE_PN0P_  (.D(_0958_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[25][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][2]$_SDFFCE_PN0P_  (.D(_0959_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[25][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][30]$_SDFFCE_PN0P_  (.D(_0960_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[25][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][31]$_SDFFCE_PN0P_  (.D(_0961_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[25][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][3]$_SDFFCE_PN0P_  (.D(_0962_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[25][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][4]$_SDFFCE_PN0P_  (.D(_0963_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[25][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][5]$_SDFFCE_PN0P_  (.D(_0964_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[25][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][6]$_SDFFCE_PN0P_  (.D(_0965_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[25][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][7]$_SDFFCE_PN0P_  (.D(_0966_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[25][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][8]$_SDFFCE_PN0P_  (.D(_0967_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[25][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[25][9]$_SDFFCE_PN0P_  (.D(_0968_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[25][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][0]$_SDFFCE_PN0P_  (.D(_0969_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[26][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][10]$_SDFFCE_PN0P_  (.D(_0970_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[26][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][11]$_SDFFCE_PN0P_  (.D(_0971_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[26][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][12]$_SDFFCE_PN0P_  (.D(_0972_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[26][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][13]$_SDFFCE_PN0P_  (.D(_0973_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[26][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][14]$_SDFFCE_PN0P_  (.D(_0974_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[26][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][15]$_SDFFCE_PN0P_  (.D(_0975_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[26][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][16]$_SDFFCE_PN0P_  (.D(_0976_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[26][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][17]$_SDFFCE_PN0P_  (.D(_0977_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[26][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][18]$_SDFFCE_PN0P_  (.D(_0978_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[26][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][19]$_SDFFCE_PN0P_  (.D(_0979_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[26][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][1]$_SDFFCE_PN0P_  (.D(_0980_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[26][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][20]$_SDFFCE_PN0P_  (.D(_0981_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[26][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][21]$_SDFFCE_PN0P_  (.D(_0982_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[26][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][22]$_SDFFCE_PN0P_  (.D(_0983_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[26][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][23]$_SDFFCE_PN0P_  (.D(_0984_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[26][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][24]$_SDFFCE_PN0P_  (.D(_0985_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[26][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][25]$_SDFFCE_PN0P_  (.D(_0986_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[26][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][26]$_SDFFCE_PN0P_  (.D(_0987_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[26][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][27]$_SDFFCE_PN0P_  (.D(_0988_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[26][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][28]$_SDFFCE_PN0P_  (.D(_0989_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[26][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][29]$_SDFFCE_PN0P_  (.D(_0990_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[26][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][2]$_SDFFCE_PN0P_  (.D(_0991_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[26][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][30]$_SDFFCE_PN0P_  (.D(_0992_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[26][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][31]$_SDFFCE_PN0P_  (.D(_0993_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[26][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][3]$_SDFFCE_PN0P_  (.D(_0994_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[26][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][4]$_SDFFCE_PN0P_  (.D(_0995_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[26][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][5]$_SDFFCE_PN0P_  (.D(_0996_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[26][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][6]$_SDFFCE_PN0P_  (.D(_0997_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[26][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][7]$_SDFFCE_PN0P_  (.D(_0998_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[26][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][8]$_SDFFCE_PN0P_  (.D(_0999_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[26][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[26][9]$_SDFFCE_PN0P_  (.D(_1000_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[26][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][0]$_SDFFCE_PN0P_  (.D(_1001_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[27][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][10]$_SDFFCE_PN0P_  (.D(_1002_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[27][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][11]$_SDFFCE_PN0P_  (.D(_1003_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[27][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][12]$_SDFFCE_PN0P_  (.D(_1004_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[27][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][13]$_SDFFCE_PN0P_  (.D(_1005_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[27][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][14]$_SDFFCE_PN0P_  (.D(_1006_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[27][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][15]$_SDFFCE_PN0P_  (.D(_1007_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[27][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][16]$_SDFFCE_PN0P_  (.D(_1008_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[27][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][17]$_SDFFCE_PN0P_  (.D(_1009_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[27][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][18]$_SDFFCE_PN0P_  (.D(_1010_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[27][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][19]$_SDFFCE_PN0P_  (.D(_1011_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[27][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][1]$_SDFFCE_PN0P_  (.D(_1012_),
    .CLK(clknet_leaf_18_clk),
    .Q(\registers[27][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][20]$_SDFFCE_PN0P_  (.D(_1013_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[27][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][21]$_SDFFCE_PN0P_  (.D(_1014_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[27][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][22]$_SDFFCE_PN0P_  (.D(_1015_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[27][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][23]$_SDFFCE_PN0P_  (.D(_1016_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[27][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][24]$_SDFFCE_PN0P_  (.D(_1017_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[27][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][25]$_SDFFCE_PN0P_  (.D(_1018_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[27][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][26]$_SDFFCE_PN0P_  (.D(_1019_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[27][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][27]$_SDFFCE_PN0P_  (.D(_1020_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[27][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][28]$_SDFFCE_PN0P_  (.D(_1021_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[27][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][29]$_SDFFCE_PN0P_  (.D(_1022_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[27][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][2]$_SDFFCE_PN0P_  (.D(_1023_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[27][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][30]$_SDFFCE_PN0P_  (.D(_1024_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[27][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][31]$_SDFFCE_PN0P_  (.D(_1025_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[27][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][3]$_SDFFCE_PN0P_  (.D(_1026_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[27][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][4]$_SDFFCE_PN0P_  (.D(_1027_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[27][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][5]$_SDFFCE_PN0P_  (.D(_1028_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[27][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][6]$_SDFFCE_PN0P_  (.D(_1029_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[27][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][7]$_SDFFCE_PN0P_  (.D(_1030_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[27][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][8]$_SDFFCE_PN0P_  (.D(_1031_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[27][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[27][9]$_SDFFCE_PN0P_  (.D(_1032_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[27][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][0]$_SDFFCE_PN0P_  (.D(_1033_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[28][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][10]$_SDFFCE_PN0P_  (.D(_1034_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[28][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][11]$_SDFFCE_PN0P_  (.D(_1035_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[28][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][12]$_SDFFCE_PN0P_  (.D(_1036_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[28][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][13]$_SDFFCE_PN0P_  (.D(_1037_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[28][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][14]$_SDFFCE_PN0P_  (.D(_1038_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[28][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][15]$_SDFFCE_PN0P_  (.D(_1039_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[28][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][16]$_SDFFCE_PN0P_  (.D(_1040_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[28][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][17]$_SDFFCE_PN0P_  (.D(_1041_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[28][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][18]$_SDFFCE_PN0P_  (.D(_1042_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[28][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][19]$_SDFFCE_PN0P_  (.D(_1043_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[28][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][1]$_SDFFCE_PN0P_  (.D(_1044_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[28][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][20]$_SDFFCE_PN0P_  (.D(_1045_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[28][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][21]$_SDFFCE_PN0P_  (.D(_1046_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[28][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][22]$_SDFFCE_PN0P_  (.D(_1047_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[28][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][23]$_SDFFCE_PN0P_  (.D(_1048_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[28][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][24]$_SDFFCE_PN0P_  (.D(_1049_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[28][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][25]$_SDFFCE_PN0P_  (.D(_1050_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[28][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][26]$_SDFFCE_PN0P_  (.D(_1051_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[28][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][27]$_SDFFCE_PN0P_  (.D(_1052_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[28][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][28]$_SDFFCE_PN0P_  (.D(_1053_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[28][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][29]$_SDFFCE_PN0P_  (.D(_1054_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[28][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][2]$_SDFFCE_PN0P_  (.D(_1055_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[28][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][30]$_SDFFCE_PN0P_  (.D(_1056_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[28][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][31]$_SDFFCE_PN0P_  (.D(_1057_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[28][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][3]$_SDFFCE_PN0P_  (.D(_1058_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[28][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][4]$_SDFFCE_PN0P_  (.D(_1059_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[28][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][5]$_SDFFCE_PN0P_  (.D(_1060_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[28][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][6]$_SDFFCE_PN0P_  (.D(_1061_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[28][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][7]$_SDFFCE_PN0P_  (.D(_1062_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[28][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][8]$_SDFFCE_PN0P_  (.D(_1063_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[28][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[28][9]$_SDFFCE_PN0P_  (.D(_1064_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[28][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][0]$_SDFFCE_PN0P_  (.D(_1065_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[29][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][10]$_SDFFCE_PN0P_  (.D(_1066_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[29][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][11]$_SDFFCE_PN0P_  (.D(_1067_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[29][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][12]$_SDFFCE_PN0P_  (.D(_1068_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[29][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][13]$_SDFFCE_PN0P_  (.D(_1069_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[29][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][14]$_SDFFCE_PN0P_  (.D(_1070_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[29][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][15]$_SDFFCE_PN0P_  (.D(_1071_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[29][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][16]$_SDFFCE_PN0P_  (.D(_1072_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[29][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][17]$_SDFFCE_PN0P_  (.D(_1073_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[29][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][18]$_SDFFCE_PN0P_  (.D(_1074_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[29][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][19]$_SDFFCE_PN0P_  (.D(_1075_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[29][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][1]$_SDFFCE_PN0P_  (.D(_1076_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[29][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][20]$_SDFFCE_PN0P_  (.D(_1077_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[29][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][21]$_SDFFCE_PN0P_  (.D(_1078_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[29][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][22]$_SDFFCE_PN0P_  (.D(_1079_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[29][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][23]$_SDFFCE_PN0P_  (.D(_1080_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[29][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][24]$_SDFFCE_PN0P_  (.D(_1081_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[29][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][25]$_SDFFCE_PN0P_  (.D(_1082_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[29][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][26]$_SDFFCE_PN0P_  (.D(_1083_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[29][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][27]$_SDFFCE_PN0P_  (.D(_1084_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[29][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][28]$_SDFFCE_PN0P_  (.D(_1085_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[29][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][29]$_SDFFCE_PN0P_  (.D(_1086_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[29][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][2]$_SDFFCE_PN0P_  (.D(_1087_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[29][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][30]$_SDFFCE_PN0P_  (.D(_0000_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[29][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][31]$_SDFFCE_PN0P_  (.D(_0001_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[29][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][3]$_SDFFCE_PN0P_  (.D(_0002_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[29][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][4]$_SDFFCE_PN0P_  (.D(_0003_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[29][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][5]$_SDFFCE_PN0P_  (.D(_0004_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[29][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][6]$_SDFFCE_PN0P_  (.D(_0005_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[29][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][7]$_SDFFCE_PN0P_  (.D(_0006_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[29][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][8]$_SDFFCE_PN0P_  (.D(_0007_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[29][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[29][9]$_SDFFCE_PN0P_  (.D(_0008_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[29][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][0]$_SDFFCE_PN0P_  (.D(_0009_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][10]$_SDFFCE_PN0P_  (.D(_0010_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][11]$_SDFFCE_PN0P_  (.D(_0011_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][12]$_SDFFCE_PN0P_  (.D(_0012_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][13]$_SDFFCE_PN0P_  (.D(_0013_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][14]$_SDFFCE_PN0P_  (.D(_0014_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][15]$_SDFFCE_PN0P_  (.D(_0015_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][16]$_SDFFCE_PN0P_  (.D(_0016_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][17]$_SDFFCE_PN0P_  (.D(_0017_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][18]$_SDFFCE_PN0P_  (.D(_0018_),
    .CLK(clknet_leaf_20_clk),
    .Q(\registers[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][19]$_SDFFCE_PN0P_  (.D(_0019_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][1]$_SDFFCE_PN0P_  (.D(_0020_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][20]$_SDFFCE_PN0P_  (.D(_0021_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][21]$_SDFFCE_PN0P_  (.D(_0022_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][22]$_SDFFCE_PN0P_  (.D(_0023_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][23]$_SDFFCE_PN0P_  (.D(_0024_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][24]$_SDFFCE_PN0P_  (.D(_0025_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][25]$_SDFFCE_PN0P_  (.D(_0026_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][26]$_SDFFCE_PN0P_  (.D(_0027_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][27]$_SDFFCE_PN0P_  (.D(_0028_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][28]$_SDFFCE_PN0P_  (.D(_0029_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][29]$_SDFFCE_PN0P_  (.D(_0030_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][2]$_SDFFCE_PN0P_  (.D(_0031_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][30]$_SDFFCE_PN0P_  (.D(_0032_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][31]$_SDFFCE_PN0P_  (.D(_0033_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][3]$_SDFFCE_PN0P_  (.D(_0034_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][4]$_SDFFCE_PN0P_  (.D(_0035_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][5]$_SDFFCE_PN0P_  (.D(_0036_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][6]$_SDFFCE_PN0P_  (.D(_0037_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][7]$_SDFFCE_PN0P_  (.D(_0038_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][8]$_SDFFCE_PN0P_  (.D(_0039_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[2][9]$_SDFFCE_PN0P_  (.D(_0040_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][0]$_SDFFCE_PN0P_  (.D(_0041_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[30][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][10]$_SDFFCE_PN0P_  (.D(_0042_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[30][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][11]$_SDFFCE_PN0P_  (.D(_0043_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[30][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][12]$_SDFFCE_PN0P_  (.D(_0044_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[30][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][13]$_SDFFCE_PN0P_  (.D(_0045_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[30][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][14]$_SDFFCE_PN0P_  (.D(_0046_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[30][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][15]$_SDFFCE_PN0P_  (.D(_0047_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[30][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][16]$_SDFFCE_PN0P_  (.D(_0048_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[30][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][17]$_SDFFCE_PN0P_  (.D(_0049_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[30][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][18]$_SDFFCE_PN0P_  (.D(_0050_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[30][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][19]$_SDFFCE_PN0P_  (.D(_0051_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[30][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][1]$_SDFFCE_PN0P_  (.D(_0052_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[30][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][20]$_SDFFCE_PN0P_  (.D(_0053_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[30][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][21]$_SDFFCE_PN0P_  (.D(_0054_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[30][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][22]$_SDFFCE_PN0P_  (.D(_0055_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[30][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][23]$_SDFFCE_PN0P_  (.D(_0056_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[30][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][24]$_SDFFCE_PN0P_  (.D(_0057_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[30][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][25]$_SDFFCE_PN0P_  (.D(_0058_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[30][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][26]$_SDFFCE_PN0P_  (.D(_0059_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[30][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][27]$_SDFFCE_PN0P_  (.D(_0060_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[30][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][28]$_SDFFCE_PN0P_  (.D(_0061_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[30][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][29]$_SDFFCE_PN0P_  (.D(_0062_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[30][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][2]$_SDFFCE_PN0P_  (.D(_0063_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[30][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][30]$_SDFFCE_PN0P_  (.D(_0064_),
    .CLK(clknet_leaf_41_clk),
    .Q(\registers[30][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][31]$_SDFFCE_PN0P_  (.D(_0065_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[30][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][3]$_SDFFCE_PN0P_  (.D(_0066_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[30][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][4]$_SDFFCE_PN0P_  (.D(_0067_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[30][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][5]$_SDFFCE_PN0P_  (.D(_0068_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[30][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][6]$_SDFFCE_PN0P_  (.D(_0069_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[30][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][7]$_SDFFCE_PN0P_  (.D(_0070_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[30][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][8]$_SDFFCE_PN0P_  (.D(_0071_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[30][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[30][9]$_SDFFCE_PN0P_  (.D(_0072_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[30][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][0]$_SDFFCE_PN0P_  (.D(_0073_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[31][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][10]$_SDFFCE_PN0P_  (.D(_0074_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[31][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][11]$_SDFFCE_PN0P_  (.D(_0075_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[31][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][12]$_SDFFCE_PN0P_  (.D(_0076_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[31][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][13]$_SDFFCE_PN0P_  (.D(_0077_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[31][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][14]$_SDFFCE_PN0P_  (.D(_0078_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[31][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][15]$_SDFFCE_PN0P_  (.D(_0079_),
    .CLK(clknet_leaf_21_clk),
    .Q(\registers[31][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][16]$_SDFFCE_PN0P_  (.D(_0080_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[31][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][17]$_SDFFCE_PN0P_  (.D(_0081_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[31][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][18]$_SDFFCE_PN0P_  (.D(_0082_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[31][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][19]$_SDFFCE_PN0P_  (.D(_0083_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[31][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][1]$_SDFFCE_PN0P_  (.D(_0084_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[31][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][20]$_SDFFCE_PN0P_  (.D(_0085_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[31][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][21]$_SDFFCE_PN0P_  (.D(_0086_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[31][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][22]$_SDFFCE_PN0P_  (.D(_0087_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[31][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][23]$_SDFFCE_PN0P_  (.D(_0088_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[31][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][24]$_SDFFCE_PN0P_  (.D(_0089_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[31][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][25]$_SDFFCE_PN0P_  (.D(_0090_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[31][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][26]$_SDFFCE_PN0P_  (.D(_0091_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[31][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][27]$_SDFFCE_PN0P_  (.D(_0092_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[31][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][28]$_SDFFCE_PN0P_  (.D(_0093_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[31][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][29]$_SDFFCE_PN0P_  (.D(_0094_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[31][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][2]$_SDFFCE_PN0P_  (.D(_0095_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[31][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][30]$_SDFFCE_PN0P_  (.D(_0096_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[31][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][31]$_SDFFCE_PN0P_  (.D(_0097_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[31][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][3]$_SDFFCE_PN0P_  (.D(_0098_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[31][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][4]$_SDFFCE_PN0P_  (.D(_0099_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[31][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][5]$_SDFFCE_PN0P_  (.D(_0100_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[31][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][6]$_SDFFCE_PN0P_  (.D(_0101_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[31][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][7]$_SDFFCE_PN0P_  (.D(_0102_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[31][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][8]$_SDFFCE_PN0P_  (.D(_0103_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[31][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[31][9]$_SDFFCE_PN0P_  (.D(_0104_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[31][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][0]$_SDFFCE_PN0P_  (.D(_0105_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][10]$_SDFFCE_PN0P_  (.D(_0106_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][11]$_SDFFCE_PN0P_  (.D(_0107_),
    .CLK(clknet_leaf_24_clk),
    .Q(\registers[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][12]$_SDFFCE_PN0P_  (.D(_0108_),
    .CLK(clknet_leaf_28_clk),
    .Q(\registers[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][13]$_SDFFCE_PN0P_  (.D(_0109_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][14]$_SDFFCE_PN0P_  (.D(_0110_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][15]$_SDFFCE_PN0P_  (.D(_0111_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][16]$_SDFFCE_PN0P_  (.D(_0112_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[3][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][17]$_SDFFCE_PN0P_  (.D(_0113_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[3][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][18]$_SDFFCE_PN0P_  (.D(_0114_),
    .CLK(clknet_leaf_19_clk),
    .Q(\registers[3][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][19]$_SDFFCE_PN0P_  (.D(_0115_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[3][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][1]$_SDFFCE_PN0P_  (.D(_0116_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][20]$_SDFFCE_PN0P_  (.D(_0117_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[3][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][21]$_SDFFCE_PN0P_  (.D(_0118_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[3][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][22]$_SDFFCE_PN0P_  (.D(_0119_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[3][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][23]$_SDFFCE_PN0P_  (.D(_0120_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[3][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][24]$_SDFFCE_PN0P_  (.D(_0121_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[3][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][25]$_SDFFCE_PN0P_  (.D(_0122_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[3][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][26]$_SDFFCE_PN0P_  (.D(_0123_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[3][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][27]$_SDFFCE_PN0P_  (.D(_0124_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[3][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][28]$_SDFFCE_PN0P_  (.D(_0125_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[3][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][29]$_SDFFCE_PN0P_  (.D(_0126_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[3][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][2]$_SDFFCE_PN0P_  (.D(_0127_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][30]$_SDFFCE_PN0P_  (.D(_0128_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[3][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][31]$_SDFFCE_PN0P_  (.D(_0129_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[3][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][3]$_SDFFCE_PN0P_  (.D(_0130_),
    .CLK(clknet_leaf_37_clk),
    .Q(\registers[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][4]$_SDFFCE_PN0P_  (.D(_0131_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][5]$_SDFFCE_PN0P_  (.D(_0132_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][6]$_SDFFCE_PN0P_  (.D(_0133_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][7]$_SDFFCE_PN0P_  (.D(_0134_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][8]$_SDFFCE_PN0P_  (.D(_0135_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[3][9]$_SDFFCE_PN0P_  (.D(_0136_),
    .CLK(clknet_leaf_27_clk),
    .Q(\registers[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][0]$_SDFFCE_PN0P_  (.D(_0137_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][10]$_SDFFCE_PN0P_  (.D(_0138_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][11]$_SDFFCE_PN0P_  (.D(_0139_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][12]$_SDFFCE_PN0P_  (.D(_0140_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][13]$_SDFFCE_PN0P_  (.D(_0141_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][14]$_SDFFCE_PN0P_  (.D(_0142_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][15]$_SDFFCE_PN0P_  (.D(_0143_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][16]$_SDFFCE_PN0P_  (.D(_0144_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[4][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][17]$_SDFFCE_PN0P_  (.D(_0145_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[4][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][18]$_SDFFCE_PN0P_  (.D(_0146_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[4][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][19]$_SDFFCE_PN0P_  (.D(_0147_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[4][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][1]$_SDFFCE_PN0P_  (.D(_0148_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][20]$_SDFFCE_PN0P_  (.D(_0149_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[4][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][21]$_SDFFCE_PN0P_  (.D(_0150_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[4][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][22]$_SDFFCE_PN0P_  (.D(_0151_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[4][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][23]$_SDFFCE_PN0P_  (.D(_0152_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[4][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][24]$_SDFFCE_PN0P_  (.D(_0153_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[4][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][25]$_SDFFCE_PN0P_  (.D(_0154_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[4][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][26]$_SDFFCE_PN0P_  (.D(_0155_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[4][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][27]$_SDFFCE_PN0P_  (.D(_0156_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[4][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][28]$_SDFFCE_PN0P_  (.D(_0157_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[4][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][29]$_SDFFCE_PN0P_  (.D(_0158_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[4][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][2]$_SDFFCE_PN0P_  (.D(_0159_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][30]$_SDFFCE_PN0P_  (.D(_0160_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[4][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][31]$_SDFFCE_PN0P_  (.D(_0161_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[4][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][3]$_SDFFCE_PN0P_  (.D(_0162_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][4]$_SDFFCE_PN0P_  (.D(_0163_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][5]$_SDFFCE_PN0P_  (.D(_0164_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][6]$_SDFFCE_PN0P_  (.D(_0165_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][7]$_SDFFCE_PN0P_  (.D(_0166_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][8]$_SDFFCE_PN0P_  (.D(_0167_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[4][9]$_SDFFCE_PN0P_  (.D(_0168_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][0]$_SDFFCE_PN0P_  (.D(_0169_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][10]$_SDFFCE_PN0P_  (.D(_0170_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][11]$_SDFFCE_PN0P_  (.D(_0171_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][12]$_SDFFCE_PN0P_  (.D(_0172_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][13]$_SDFFCE_PN0P_  (.D(_0173_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][14]$_SDFFCE_PN0P_  (.D(_0174_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][15]$_SDFFCE_PN0P_  (.D(_0175_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][16]$_SDFFCE_PN0P_  (.D(_0176_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[5][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][17]$_SDFFCE_PN0P_  (.D(_0177_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[5][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][18]$_SDFFCE_PN0P_  (.D(_0178_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[5][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][19]$_SDFFCE_PN0P_  (.D(_0179_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[5][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][1]$_SDFFCE_PN0P_  (.D(_0180_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][20]$_SDFFCE_PN0P_  (.D(_0181_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[5][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][21]$_SDFFCE_PN0P_  (.D(_0182_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[5][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][22]$_SDFFCE_PN0P_  (.D(_0183_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[5][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][23]$_SDFFCE_PN0P_  (.D(_0184_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[5][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][24]$_SDFFCE_PN0P_  (.D(_0185_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[5][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][25]$_SDFFCE_PN0P_  (.D(_0186_),
    .CLK(clknet_leaf_8_clk),
    .Q(\registers[5][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][26]$_SDFFCE_PN0P_  (.D(_0187_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[5][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][27]$_SDFFCE_PN0P_  (.D(_0188_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[5][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][28]$_SDFFCE_PN0P_  (.D(_0189_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[5][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][29]$_SDFFCE_PN0P_  (.D(_0190_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[5][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][2]$_SDFFCE_PN0P_  (.D(_0191_),
    .CLK(clknet_leaf_2_clk),
    .Q(\registers[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][30]$_SDFFCE_PN0P_  (.D(_0192_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[5][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][31]$_SDFFCE_PN0P_  (.D(_0193_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[5][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][3]$_SDFFCE_PN0P_  (.D(_0194_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][4]$_SDFFCE_PN0P_  (.D(_0195_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][5]$_SDFFCE_PN0P_  (.D(_0196_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][6]$_SDFFCE_PN0P_  (.D(_0197_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][7]$_SDFFCE_PN0P_  (.D(_0198_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][8]$_SDFFCE_PN0P_  (.D(_0199_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[5][9]$_SDFFCE_PN0P_  (.D(_0200_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][0]$_SDFFCE_PN0P_  (.D(_0201_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][10]$_SDFFCE_PN0P_  (.D(_0202_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][11]$_SDFFCE_PN0P_  (.D(_0203_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][12]$_SDFFCE_PN0P_  (.D(_0204_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][13]$_SDFFCE_PN0P_  (.D(_0205_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][14]$_SDFFCE_PN0P_  (.D(_0206_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][15]$_SDFFCE_PN0P_  (.D(_0207_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][16]$_SDFFCE_PN0P_  (.D(_0208_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[6][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][17]$_SDFFCE_PN0P_  (.D(_0209_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[6][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][18]$_SDFFCE_PN0P_  (.D(_0210_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[6][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][19]$_SDFFCE_PN0P_  (.D(_0211_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[6][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][1]$_SDFFCE_PN0P_  (.D(_0212_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][20]$_SDFFCE_PN0P_  (.D(_0213_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[6][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][21]$_SDFFCE_PN0P_  (.D(_0214_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[6][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][22]$_SDFFCE_PN0P_  (.D(_0215_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[6][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][23]$_SDFFCE_PN0P_  (.D(_0216_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[6][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][24]$_SDFFCE_PN0P_  (.D(_0217_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[6][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][25]$_SDFFCE_PN0P_  (.D(_0218_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[6][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][26]$_SDFFCE_PN0P_  (.D(_0219_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[6][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][27]$_SDFFCE_PN0P_  (.D(_0220_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[6][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][28]$_SDFFCE_PN0P_  (.D(_0221_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[6][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][29]$_SDFFCE_PN0P_  (.D(_0222_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[6][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][2]$_SDFFCE_PN0P_  (.D(_0223_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][30]$_SDFFCE_PN0P_  (.D(_0224_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[6][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][31]$_SDFFCE_PN0P_  (.D(_0225_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[6][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][3]$_SDFFCE_PN0P_  (.D(_0226_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][4]$_SDFFCE_PN0P_  (.D(_0227_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][5]$_SDFFCE_PN0P_  (.D(_0228_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][6]$_SDFFCE_PN0P_  (.D(_0229_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][7]$_SDFFCE_PN0P_  (.D(_0230_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][8]$_SDFFCE_PN0P_  (.D(_0231_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[6][9]$_SDFFCE_PN0P_  (.D(_0232_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][0]$_SDFFCE_PN0P_  (.D(_0233_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][10]$_SDFFCE_PN0P_  (.D(_0234_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][11]$_SDFFCE_PN0P_  (.D(_0235_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][12]$_SDFFCE_PN0P_  (.D(_0236_),
    .CLK(clknet_leaf_26_clk),
    .Q(\registers[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][13]$_SDFFCE_PN0P_  (.D(_0237_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][14]$_SDFFCE_PN0P_  (.D(_0238_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][15]$_SDFFCE_PN0P_  (.D(_0239_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][16]$_SDFFCE_PN0P_  (.D(_0240_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[7][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][17]$_SDFFCE_PN0P_  (.D(_0241_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[7][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][18]$_SDFFCE_PN0P_  (.D(_0242_),
    .CLK(clknet_leaf_17_clk),
    .Q(\registers[7][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][19]$_SDFFCE_PN0P_  (.D(_0243_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[7][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][1]$_SDFFCE_PN0P_  (.D(_0244_),
    .CLK(clknet_leaf_13_clk),
    .Q(\registers[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][20]$_SDFFCE_PN0P_  (.D(_0245_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[7][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][21]$_SDFFCE_PN0P_  (.D(_0246_),
    .CLK(clknet_leaf_12_clk),
    .Q(\registers[7][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][22]$_SDFFCE_PN0P_  (.D(_0247_),
    .CLK(clknet_leaf_11_clk),
    .Q(\registers[7][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][23]$_SDFFCE_PN0P_  (.D(_0248_),
    .CLK(clknet_leaf_10_clk),
    .Q(\registers[7][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][24]$_SDFFCE_PN0P_  (.D(_0249_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[7][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][25]$_SDFFCE_PN0P_  (.D(_0250_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[7][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][26]$_SDFFCE_PN0P_  (.D(_0251_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[7][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][27]$_SDFFCE_PN0P_  (.D(_0252_),
    .CLK(clknet_leaf_7_clk),
    .Q(\registers[7][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][28]$_SDFFCE_PN0P_  (.D(_0253_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[7][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][29]$_SDFFCE_PN0P_  (.D(_0254_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[7][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][2]$_SDFFCE_PN0P_  (.D(_0255_),
    .CLK(clknet_leaf_3_clk),
    .Q(\registers[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][30]$_SDFFCE_PN0P_  (.D(_0256_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[7][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][31]$_SDFFCE_PN0P_  (.D(_0257_),
    .CLK(clknet_leaf_4_clk),
    .Q(\registers[7][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][3]$_SDFFCE_PN0P_  (.D(_0258_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][4]$_SDFFCE_PN0P_  (.D(_0259_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][5]$_SDFFCE_PN0P_  (.D(_0260_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][6]$_SDFFCE_PN0P_  (.D(_0261_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][7]$_SDFFCE_PN0P_  (.D(_0262_),
    .CLK(clknet_leaf_36_clk),
    .Q(\registers[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][8]$_SDFFCE_PN0P_  (.D(_0263_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[7][9]$_SDFFCE_PN0P_  (.D(_0264_),
    .CLK(clknet_leaf_35_clk),
    .Q(\registers[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][0]$_SDFFCE_PN0P_  (.D(_0265_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[8][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][10]$_SDFFCE_PN0P_  (.D(_0266_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[8][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][11]$_SDFFCE_PN0P_  (.D(_0267_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[8][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][12]$_SDFFCE_PN0P_  (.D(_0268_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[8][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][13]$_SDFFCE_PN0P_  (.D(_0269_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[8][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][14]$_SDFFCE_PN0P_  (.D(_0270_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[8][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][15]$_SDFFCE_PN0P_  (.D(_0271_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[8][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][16]$_SDFFCE_PN0P_  (.D(_0272_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[8][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][17]$_SDFFCE_PN0P_  (.D(_0273_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[8][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][18]$_SDFFCE_PN0P_  (.D(_0274_),
    .CLK(clknet_leaf_25_clk),
    .Q(\registers[8][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][19]$_SDFFCE_PN0P_  (.D(_0275_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[8][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][1]$_SDFFCE_PN0P_  (.D(_0276_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[8][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][20]$_SDFFCE_PN0P_  (.D(_0277_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[8][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][21]$_SDFFCE_PN0P_  (.D(_0278_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[8][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][22]$_SDFFCE_PN0P_  (.D(_0279_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[8][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][23]$_SDFFCE_PN0P_  (.D(_0280_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[8][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][24]$_SDFFCE_PN0P_  (.D(_0281_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[8][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][25]$_SDFFCE_PN0P_  (.D(_0282_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[8][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][26]$_SDFFCE_PN0P_  (.D(_0283_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[8][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][27]$_SDFFCE_PN0P_  (.D(_0284_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[8][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][28]$_SDFFCE_PN0P_  (.D(_0285_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[8][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][29]$_SDFFCE_PN0P_  (.D(_0286_),
    .CLK(clknet_leaf_1_clk),
    .Q(\registers[8][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][2]$_SDFFCE_PN0P_  (.D(_0287_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[8][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][30]$_SDFFCE_PN0P_  (.D(_0288_),
    .CLK(clknet_leaf_40_clk),
    .Q(\registers[8][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][31]$_SDFFCE_PN0P_  (.D(_0289_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[8][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][3]$_SDFFCE_PN0P_  (.D(_0290_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[8][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][4]$_SDFFCE_PN0P_  (.D(_0291_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[8][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][5]$_SDFFCE_PN0P_  (.D(_0292_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[8][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][6]$_SDFFCE_PN0P_  (.D(_0293_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[8][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][7]$_SDFFCE_PN0P_  (.D(_0294_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[8][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][8]$_SDFFCE_PN0P_  (.D(_0295_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[8][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[8][9]$_SDFFCE_PN0P_  (.D(_0296_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[8][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][0]$_SDFFCE_PN0P_  (.D(_0297_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[9][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][10]$_SDFFCE_PN0P_  (.D(_0298_),
    .CLK(clknet_leaf_30_clk),
    .Q(\registers[9][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][11]$_SDFFCE_PN0P_  (.D(_0299_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[9][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][12]$_SDFFCE_PN0P_  (.D(_0300_),
    .CLK(clknet_leaf_29_clk),
    .Q(\registers[9][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][13]$_SDFFCE_PN0P_  (.D(_0301_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[9][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][14]$_SDFFCE_PN0P_  (.D(_0302_),
    .CLK(clknet_leaf_23_clk),
    .Q(\registers[9][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][15]$_SDFFCE_PN0P_  (.D(_0303_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[9][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][16]$_SDFFCE_PN0P_  (.D(_0304_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[9][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][17]$_SDFFCE_PN0P_  (.D(_0305_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[9][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][18]$_SDFFCE_PN0P_  (.D(_0306_),
    .CLK(clknet_leaf_22_clk),
    .Q(\registers[9][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][19]$_SDFFCE_PN0P_  (.D(_0307_),
    .CLK(clknet_leaf_16_clk),
    .Q(\registers[9][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][1]$_SDFFCE_PN0P_  (.D(_0308_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[9][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][20]$_SDFFCE_PN0P_  (.D(_0309_),
    .CLK(clknet_leaf_15_clk),
    .Q(\registers[9][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][21]$_SDFFCE_PN0P_  (.D(_0310_),
    .CLK(clknet_leaf_14_clk),
    .Q(\registers[9][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][22]$_SDFFCE_PN0P_  (.D(_0311_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[9][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][23]$_SDFFCE_PN0P_  (.D(_0312_),
    .CLK(clknet_leaf_9_clk),
    .Q(\registers[9][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][24]$_SDFFCE_PN0P_  (.D(_0313_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[9][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][25]$_SDFFCE_PN0P_  (.D(_0314_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[9][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][26]$_SDFFCE_PN0P_  (.D(_0315_),
    .CLK(clknet_leaf_5_clk),
    .Q(\registers[9][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][27]$_SDFFCE_PN0P_  (.D(_0316_),
    .CLK(clknet_leaf_6_clk),
    .Q(\registers[9][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][28]$_SDFFCE_PN0P_  (.D(_0317_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[9][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][29]$_SDFFCE_PN0P_  (.D(_0318_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[9][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][2]$_SDFFCE_PN0P_  (.D(_0319_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[9][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][30]$_SDFFCE_PN0P_  (.D(_0320_),
    .CLK(clknet_leaf_0_clk),
    .Q(\registers[9][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][31]$_SDFFCE_PN0P_  (.D(_0321_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[9][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][3]$_SDFFCE_PN0P_  (.D(_0322_),
    .CLK(clknet_leaf_39_clk),
    .Q(\registers[9][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][4]$_SDFFCE_PN0P_  (.D(_0323_),
    .CLK(clknet_leaf_38_clk),
    .Q(\registers[9][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][5]$_SDFFCE_PN0P_  (.D(_0324_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[9][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][6]$_SDFFCE_PN0P_  (.D(_0325_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[9][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][7]$_SDFFCE_PN0P_  (.D(_0326_),
    .CLK(clknet_leaf_33_clk),
    .Q(\registers[9][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][8]$_SDFFCE_PN0P_  (.D(_0327_),
    .CLK(clknet_leaf_32_clk),
    .Q(\registers[9][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \registers[9][9]$_SDFFCE_PN0P_  (.D(_0328_),
    .CLK(clknet_leaf_31_clk),
    .Q(\registers[9][9] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_961 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input1 (.I(read_addr1[2]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input2 (.I(read_addr1[3]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 input3 (.I(net114),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input4 (.I(read_addr2[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input5 (.I(read_addr2[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input6 (.I(read_addr2[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(read_en1),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input8 (.I(read_en2),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input9 (.I(rst_n),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input10 (.I(write_addr[0]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input11 (.I(write_addr[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input12 (.I(write_addr[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input13 (.I(write_addr[3]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input14 (.I(write_addr[4]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input15 (.I(net115),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input16 (.I(net126),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input17 (.I(net116),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input18 (.I(net129),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input19 (.I(net117),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(net124),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input21 (.I(net125),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(net122),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input23 (.I(net137),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input24 (.I(net119),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input25 (.I(net121),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input26 (.I(net131),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input27 (.I(net120),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input28 (.I(net144),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input29 (.I(net140),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input30 (.I(net142),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input31 (.I(net136),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input32 (.I(net141),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input33 (.I(net143),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input34 (.I(net134),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input35 (.I(net123),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input36 (.I(net132),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input37 (.I(net128),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input38 (.I(net118),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input39 (.I(net133),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input40 (.I(net138),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input41 (.I(net113),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input42 (.I(net112),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input43 (.I(net135),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(net127),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input45 (.I(net139),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input46 (.I(net130),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input47 (.I(write_en),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net48),
    .Z(read_data1[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net49),
    .Z(read_data1[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net50),
    .Z(read_data1[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net51),
    .Z(read_data1[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net52),
    .Z(read_data1[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net53),
    .Z(read_data1[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net54),
    .Z(read_data1[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net55),
    .Z(read_data1[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net56),
    .Z(read_data1[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net57),
    .Z(read_data1[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net58),
    .Z(read_data1[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net59),
    .Z(read_data1[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net60),
    .Z(read_data1[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net61),
    .Z(read_data1[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net62),
    .Z(read_data1[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net63),
    .Z(read_data1[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net64),
    .Z(read_data1[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net65),
    .Z(read_data1[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net66),
    .Z(read_data1[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(read_data1[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(read_data1[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(read_data1[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(read_data1[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net71),
    .Z(read_data1[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net72),
    .Z(read_data1[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net73),
    .Z(read_data1[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net74),
    .Z(read_data1[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net75),
    .Z(read_data1[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net76),
    .Z(read_data1[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net77),
    .Z(read_data1[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net78),
    .Z(read_data1[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net79),
    .Z(read_data1[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net80),
    .Z(read_data2[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net81),
    .Z(read_data2[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net82),
    .Z(read_data2[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net83),
    .Z(read_data2[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net84),
    .Z(read_data2[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net85),
    .Z(read_data2[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net86),
    .Z(read_data2[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net87),
    .Z(read_data2[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net88),
    .Z(read_data2[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net89),
    .Z(read_data2[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net90),
    .Z(read_data2[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net91),
    .Z(read_data2[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net92),
    .Z(read_data2[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net93),
    .Z(read_data2[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net94),
    .Z(read_data2[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net95),
    .Z(read_data2[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net96),
    .Z(read_data2[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net97),
    .Z(read_data2[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net98),
    .Z(read_data2[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net99),
    .Z(read_data2[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net100),
    .Z(read_data2[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net101),
    .Z(read_data2[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net102),
    .Z(read_data2[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net103),
    .Z(read_data2[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net104),
    .Z(read_data2[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net105),
    .Z(read_data2[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net106),
    .Z(read_data2[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net107),
    .Z(read_data2[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net108),
    .Z(read_data2[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net109),
    .Z(read_data2[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net110),
    .Z(read_data2[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net111),
    .Z(read_data2[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_30_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_31_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_32_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_33_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_34_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_35_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_36_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_37_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_38_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_39_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_40_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_41_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload0 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload1 (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload2 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload3 (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload4 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload5 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload6 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload7 (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload8 (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload9 (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload10 (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload11 (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload12 (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload13 (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload14 (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload15 (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload16 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload17 (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload18 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload19 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload20 (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload21 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload22 (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload23 (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload24 (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload25 (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload26 (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload27 (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload28 (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload29 (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload30 (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload31 (.I(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload32 (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload33 (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload34 (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload35 (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload36 (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload37 (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload38 (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload39 (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold1 (.I(write_data[5]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(write_data[4]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(read_addr1[4]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold4 (.I(write_data[0]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold5 (.I(write_data[11]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold6 (.I(write_data[13]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold7 (.I(write_data[30]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold8 (.I(write_data[18]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold9 (.I(write_data[20]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold10 (.I(write_data[19]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold11 (.I(write_data[16]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold12 (.I(write_data[28]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold13 (.I(write_data[14]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold14 (.I(write_data[15]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold15 (.I(write_data[10]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold16 (.I(write_data[7]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold17 (.I(write_data[2]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold18 (.I(write_data[12]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold19 (.I(write_data[9]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold20 (.I(write_data[1]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold21 (.I(write_data[29]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold22 (.I(write_data[31]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold23 (.I(write_data[27]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold24 (.I(write_data[6]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold25 (.I(write_data[24]),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold26 (.I(write_data[17]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold27 (.I(write_data[3]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold28 (.I(write_data[8]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold29 (.I(write_data[22]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold30 (.I(write_data[25]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold31 (.I(write_data[23]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold32 (.I(write_data[26]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold33 (.I(write_data[21]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net56));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net104));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net109));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1434 ();
endmodule
