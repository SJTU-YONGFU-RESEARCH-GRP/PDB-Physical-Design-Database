module dma_controller (clk,
    debug_has_active_channels,
    rst_n,
    channel_busy,
    channel_done,
    channel_dst_addr,
    channel_enable,
    channel_error,
    channel_length,
    channel_mode,
    channel_src_addr,
    channel_start,
    debug_active_channels,
    debug_channel_state,
    debug_transfer_count,
    dst_addr,
    dst_wdata,
    dst_wready,
    dst_write,
    dst_wstrb,
    src_addr,
    src_rdata,
    src_read,
    src_rready,
    src_rvalid);
 input clk;
 output debug_has_active_channels;
 input rst_n;
 output [3:0] channel_busy;
 output [3:0] channel_done;
 input [127:0] channel_dst_addr;
 input [3:0] channel_enable;
 output [3:0] channel_error;
 input [127:0] channel_length;
 input [7:0] channel_mode;
 input [127:0] channel_src_addr;
 input [3:0] channel_start;
 output [3:0] debug_active_channels;
 output [11:0] debug_channel_state;
 output [127:0] debug_transfer_count;
 output [127:0] dst_addr;
 output [127:0] dst_wdata;
 input [3:0] dst_wready;
 output [3:0] dst_write;
 output [15:0] dst_wstrb;
 output [127:0] src_addr;
 input [127:0] src_rdata;
 output [3:0] src_read;
 output [3:0] src_rready;
 input [3:0] src_rvalid;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire net221;
 wire _1453_;
 wire _1454_;
 wire net219;
 wire net217;
 wire net216;
 wire _1458_;
 wire _1459_;
 wire net214;
 wire net213;
 wire net212;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire net210;
 wire net209;
 wire net208;
 wire _1469_;
 wire _1470_;
 wire net207;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire net206;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire net205;
 wire _1481_;
 wire net204;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire net203;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire net202;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire net201;
 wire net200;
 wire _1505_;
 wire net199;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire net198;
 wire _1515_;
 wire _1516_;
 wire net197;
 wire _1518_;
 wire net196;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire net195;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire net194;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire net193;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire net192;
 wire net191;
 wire _1607_;
 wire net190;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire net189;
 wire _1613_;
 wire net188;
 wire _1615_;
 wire net187;
 wire _1617_;
 wire _1618_;
 wire net186;
 wire _1620_;
 wire _1621_;
 wire net185;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire net184;
 wire _1629_;
 wire net183;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire net182;
 wire _1641_;
 wire net181;
 wire _1643_;
 wire net180;
 wire _1645_;
 wire net179;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire net178;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire net177;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire net176;
 wire net175;
 wire _1736_;
 wire net174;
 wire _1738_;
 wire net173;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire net172;
 wire _1744_;
 wire net171;
 wire net170;
 wire _1747_;
 wire _1748_;
 wire net169;
 wire net168;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire net167;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire net166;
 wire _1768_;
 wire _1769_;
 wire net165;
 wire _1771_;
 wire _1772_;
 wire net164;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire net163;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire net162;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire net161;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire net160;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire net159;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire net158;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire net157;
 wire net156;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire net155;
 wire _1874_;
 wire net154;
 wire _1876_;
 wire net153;
 wire net152;
 wire _1879_;
 wire _1880_;
 wire net151;
 wire net150;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire net149;
 wire _1889_;
 wire _1890_;
 wire net148;
 wire net147;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire net146;
 wire _1905_;
 wire net145;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire net144;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire net143;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire net142;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire net141;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire net140;
 wire _1980_;
 wire net139;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire net138;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire net137;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire net136;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire net135;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire net134;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire net133;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire net132;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire net131;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire net130;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire net129;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire net128;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire net127;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire net126;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire net125;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire net124;
 wire _2249_;
 wire _2250_;
 wire net123;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire net122;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire net121;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire net120;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire net119;
 wire _2393_;
 wire net118;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire net117;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire net116;
 wire _2468_;
 wire net115;
 wire _2470_;
 wire net114;
 wire _2472_;
 wire net113;
 wire _2474_;
 wire net112;
 wire _2476_;
 wire net111;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire net110;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire net109;
 wire _2513_;
 wire net108;
 wire _2515_;
 wire _2516_;
 wire net107;
 wire _2518_;
 wire net106;
 wire _2520_;
 wire _2521_;
 wire net105;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire net104;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire net103;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire net102;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire net101;
 wire net100;
 wire _2610_;
 wire net99;
 wire _2612_;
 wire net98;
 wire _2614_;
 wire net97;
 wire _2616_;
 wire _2617_;
 wire net96;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire net95;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire net94;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire net93;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire net92;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire net91;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire net90;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire net89;
 wire net88;
 wire _2745_;
 wire net87;
 wire _2747_;
 wire net86;
 wire _2749_;
 wire net85;
 wire _2751_;
 wire net84;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire net83;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire net82;
 wire _2773_;
 wire net81;
 wire _2775_;
 wire _2776_;
 wire net80;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire net79;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire net78;
 wire _2792_;
 wire net77;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire net76;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire net75;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire net74;
 wire net73;
 wire _2896_;
 wire net72;
 wire _2898_;
 wire net71;
 wire _2900_;
 wire net70;
 wire _2902_;
 wire net69;
 wire net68;
 wire _2905_;
 wire net67;
 wire _2907_;
 wire _2908_;
 wire net66;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire net65;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire net64;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire net63;
 wire _2932_;
 wire net62;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire net61;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire net60;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire net59;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire net58;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire net57;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire net56;
 wire net55;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire net54;
 wire net53;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire net52;
 wire net51;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire net50;
 wire net49;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire net48;
 wire net47;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire net46;
 wire net45;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire net44;
 wire net43;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire _3372_;
 wire net34;
 wire net33;
 wire _3375_;
 wire net32;
 wire net31;
 wire _3378_;
 wire net30;
 wire net29;
 wire _3381_;
 wire net28;
 wire net27;
 wire _3384_;
 wire net26;
 wire net25;
 wire _3387_;
 wire _3388_;
 wire net24;
 wire net23;
 wire net22;
 wire _3392_;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire _3406_;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire net220;
 wire _3425_;
 wire _3426_;
 wire net211;
 wire _3428_;
 wire net215;
 wire net218;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire \active_channel_count[0] ;
 wire \active_channel_count[1] ;
 wire \active_channel_count[2] ;
 wire \active_channel_count[3] ;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire \current_dst_addr[0][0] ;
 wire \current_dst_addr[0][10] ;
 wire \current_dst_addr[0][11] ;
 wire \current_dst_addr[0][12] ;
 wire \current_dst_addr[0][13] ;
 wire \current_dst_addr[0][14] ;
 wire \current_dst_addr[0][15] ;
 wire \current_dst_addr[0][16] ;
 wire \current_dst_addr[0][17] ;
 wire \current_dst_addr[0][18] ;
 wire \current_dst_addr[0][19] ;
 wire \current_dst_addr[0][1] ;
 wire \current_dst_addr[0][20] ;
 wire \current_dst_addr[0][21] ;
 wire \current_dst_addr[0][22] ;
 wire \current_dst_addr[0][23] ;
 wire \current_dst_addr[0][24] ;
 wire \current_dst_addr[0][25] ;
 wire \current_dst_addr[0][26] ;
 wire \current_dst_addr[0][27] ;
 wire \current_dst_addr[0][28] ;
 wire \current_dst_addr[0][29] ;
 wire \current_dst_addr[0][2] ;
 wire \current_dst_addr[0][30] ;
 wire \current_dst_addr[0][31] ;
 wire \current_dst_addr[0][3] ;
 wire \current_dst_addr[0][4] ;
 wire \current_dst_addr[0][5] ;
 wire \current_dst_addr[0][6] ;
 wire \current_dst_addr[0][7] ;
 wire \current_dst_addr[0][8] ;
 wire \current_dst_addr[0][9] ;
 wire \current_dst_addr[1][0] ;
 wire \current_dst_addr[1][10] ;
 wire \current_dst_addr[1][11] ;
 wire \current_dst_addr[1][12] ;
 wire \current_dst_addr[1][13] ;
 wire \current_dst_addr[1][14] ;
 wire \current_dst_addr[1][15] ;
 wire \current_dst_addr[1][16] ;
 wire \current_dst_addr[1][17] ;
 wire \current_dst_addr[1][18] ;
 wire \current_dst_addr[1][19] ;
 wire \current_dst_addr[1][1] ;
 wire \current_dst_addr[1][20] ;
 wire \current_dst_addr[1][21] ;
 wire \current_dst_addr[1][22] ;
 wire \current_dst_addr[1][23] ;
 wire \current_dst_addr[1][24] ;
 wire \current_dst_addr[1][25] ;
 wire \current_dst_addr[1][26] ;
 wire \current_dst_addr[1][27] ;
 wire \current_dst_addr[1][28] ;
 wire \current_dst_addr[1][29] ;
 wire \current_dst_addr[1][2] ;
 wire \current_dst_addr[1][30] ;
 wire \current_dst_addr[1][31] ;
 wire \current_dst_addr[1][3] ;
 wire \current_dst_addr[1][4] ;
 wire \current_dst_addr[1][5] ;
 wire \current_dst_addr[1][6] ;
 wire \current_dst_addr[1][7] ;
 wire \current_dst_addr[1][8] ;
 wire \current_dst_addr[1][9] ;
 wire \current_dst_addr[2][0] ;
 wire \current_dst_addr[2][10] ;
 wire \current_dst_addr[2][11] ;
 wire \current_dst_addr[2][12] ;
 wire \current_dst_addr[2][13] ;
 wire \current_dst_addr[2][14] ;
 wire \current_dst_addr[2][15] ;
 wire \current_dst_addr[2][16] ;
 wire \current_dst_addr[2][17] ;
 wire \current_dst_addr[2][18] ;
 wire \current_dst_addr[2][19] ;
 wire \current_dst_addr[2][1] ;
 wire \current_dst_addr[2][20] ;
 wire \current_dst_addr[2][21] ;
 wire \current_dst_addr[2][22] ;
 wire \current_dst_addr[2][23] ;
 wire \current_dst_addr[2][24] ;
 wire \current_dst_addr[2][25] ;
 wire \current_dst_addr[2][26] ;
 wire \current_dst_addr[2][27] ;
 wire \current_dst_addr[2][28] ;
 wire \current_dst_addr[2][29] ;
 wire \current_dst_addr[2][2] ;
 wire \current_dst_addr[2][30] ;
 wire \current_dst_addr[2][31] ;
 wire \current_dst_addr[2][3] ;
 wire \current_dst_addr[2][4] ;
 wire \current_dst_addr[2][5] ;
 wire \current_dst_addr[2][6] ;
 wire \current_dst_addr[2][7] ;
 wire \current_dst_addr[2][8] ;
 wire \current_dst_addr[2][9] ;
 wire \current_dst_addr[3][0] ;
 wire \current_dst_addr[3][10] ;
 wire \current_dst_addr[3][11] ;
 wire \current_dst_addr[3][12] ;
 wire \current_dst_addr[3][13] ;
 wire \current_dst_addr[3][14] ;
 wire \current_dst_addr[3][15] ;
 wire \current_dst_addr[3][16] ;
 wire \current_dst_addr[3][17] ;
 wire \current_dst_addr[3][18] ;
 wire \current_dst_addr[3][19] ;
 wire \current_dst_addr[3][1] ;
 wire \current_dst_addr[3][20] ;
 wire \current_dst_addr[3][21] ;
 wire \current_dst_addr[3][22] ;
 wire \current_dst_addr[3][23] ;
 wire \current_dst_addr[3][24] ;
 wire \current_dst_addr[3][25] ;
 wire \current_dst_addr[3][26] ;
 wire \current_dst_addr[3][27] ;
 wire \current_dst_addr[3][28] ;
 wire \current_dst_addr[3][29] ;
 wire \current_dst_addr[3][2] ;
 wire \current_dst_addr[3][30] ;
 wire \current_dst_addr[3][31] ;
 wire \current_dst_addr[3][3] ;
 wire \current_dst_addr[3][4] ;
 wire \current_dst_addr[3][5] ;
 wire \current_dst_addr[3][6] ;
 wire \current_dst_addr[3][7] ;
 wire \current_dst_addr[3][8] ;
 wire \current_dst_addr[3][9] ;
 wire \current_src_addr[0][0] ;
 wire \current_src_addr[0][10] ;
 wire \current_src_addr[0][11] ;
 wire \current_src_addr[0][12] ;
 wire \current_src_addr[0][13] ;
 wire \current_src_addr[0][14] ;
 wire \current_src_addr[0][15] ;
 wire \current_src_addr[0][16] ;
 wire \current_src_addr[0][17] ;
 wire \current_src_addr[0][18] ;
 wire \current_src_addr[0][19] ;
 wire \current_src_addr[0][1] ;
 wire \current_src_addr[0][20] ;
 wire \current_src_addr[0][21] ;
 wire \current_src_addr[0][22] ;
 wire \current_src_addr[0][23] ;
 wire \current_src_addr[0][24] ;
 wire \current_src_addr[0][25] ;
 wire \current_src_addr[0][26] ;
 wire \current_src_addr[0][27] ;
 wire \current_src_addr[0][28] ;
 wire \current_src_addr[0][29] ;
 wire \current_src_addr[0][2] ;
 wire \current_src_addr[0][30] ;
 wire \current_src_addr[0][31] ;
 wire \current_src_addr[0][3] ;
 wire \current_src_addr[0][4] ;
 wire \current_src_addr[0][5] ;
 wire \current_src_addr[0][6] ;
 wire \current_src_addr[0][7] ;
 wire \current_src_addr[0][8] ;
 wire \current_src_addr[0][9] ;
 wire \current_src_addr[1][0] ;
 wire \current_src_addr[1][10] ;
 wire \current_src_addr[1][11] ;
 wire \current_src_addr[1][12] ;
 wire \current_src_addr[1][13] ;
 wire \current_src_addr[1][14] ;
 wire \current_src_addr[1][15] ;
 wire \current_src_addr[1][16] ;
 wire \current_src_addr[1][17] ;
 wire \current_src_addr[1][18] ;
 wire \current_src_addr[1][19] ;
 wire \current_src_addr[1][1] ;
 wire \current_src_addr[1][20] ;
 wire \current_src_addr[1][21] ;
 wire \current_src_addr[1][22] ;
 wire \current_src_addr[1][23] ;
 wire \current_src_addr[1][24] ;
 wire \current_src_addr[1][25] ;
 wire \current_src_addr[1][26] ;
 wire \current_src_addr[1][27] ;
 wire \current_src_addr[1][28] ;
 wire \current_src_addr[1][29] ;
 wire \current_src_addr[1][2] ;
 wire \current_src_addr[1][30] ;
 wire \current_src_addr[1][31] ;
 wire \current_src_addr[1][3] ;
 wire \current_src_addr[1][4] ;
 wire \current_src_addr[1][5] ;
 wire \current_src_addr[1][6] ;
 wire \current_src_addr[1][7] ;
 wire \current_src_addr[1][8] ;
 wire \current_src_addr[1][9] ;
 wire \current_src_addr[2][0] ;
 wire \current_src_addr[2][10] ;
 wire \current_src_addr[2][11] ;
 wire \current_src_addr[2][12] ;
 wire \current_src_addr[2][13] ;
 wire \current_src_addr[2][14] ;
 wire \current_src_addr[2][15] ;
 wire \current_src_addr[2][16] ;
 wire \current_src_addr[2][17] ;
 wire \current_src_addr[2][18] ;
 wire \current_src_addr[2][19] ;
 wire \current_src_addr[2][1] ;
 wire \current_src_addr[2][20] ;
 wire \current_src_addr[2][21] ;
 wire \current_src_addr[2][22] ;
 wire \current_src_addr[2][23] ;
 wire \current_src_addr[2][24] ;
 wire \current_src_addr[2][25] ;
 wire \current_src_addr[2][26] ;
 wire \current_src_addr[2][27] ;
 wire \current_src_addr[2][28] ;
 wire \current_src_addr[2][29] ;
 wire \current_src_addr[2][2] ;
 wire \current_src_addr[2][30] ;
 wire \current_src_addr[2][31] ;
 wire \current_src_addr[2][3] ;
 wire \current_src_addr[2][4] ;
 wire \current_src_addr[2][5] ;
 wire \current_src_addr[2][6] ;
 wire \current_src_addr[2][7] ;
 wire \current_src_addr[2][8] ;
 wire \current_src_addr[2][9] ;
 wire \current_src_addr[3][0] ;
 wire \current_src_addr[3][10] ;
 wire \current_src_addr[3][11] ;
 wire \current_src_addr[3][12] ;
 wire \current_src_addr[3][13] ;
 wire \current_src_addr[3][14] ;
 wire \current_src_addr[3][15] ;
 wire \current_src_addr[3][16] ;
 wire \current_src_addr[3][17] ;
 wire \current_src_addr[3][18] ;
 wire \current_src_addr[3][19] ;
 wire \current_src_addr[3][1] ;
 wire \current_src_addr[3][20] ;
 wire \current_src_addr[3][21] ;
 wire \current_src_addr[3][22] ;
 wire \current_src_addr[3][23] ;
 wire \current_src_addr[3][24] ;
 wire \current_src_addr[3][25] ;
 wire \current_src_addr[3][26] ;
 wire \current_src_addr[3][27] ;
 wire \current_src_addr[3][28] ;
 wire \current_src_addr[3][29] ;
 wire \current_src_addr[3][2] ;
 wire \current_src_addr[3][30] ;
 wire \current_src_addr[3][31] ;
 wire \current_src_addr[3][3] ;
 wire \current_src_addr[3][4] ;
 wire \current_src_addr[3][5] ;
 wire \current_src_addr[3][6] ;
 wire \current_src_addr[3][7] ;
 wire \current_src_addr[3][8] ;
 wire \current_src_addr[3][9] ;
 wire \data_buffer[0][0] ;
 wire \data_buffer[0][10] ;
 wire \data_buffer[0][11] ;
 wire \data_buffer[0][12] ;
 wire \data_buffer[0][13] ;
 wire \data_buffer[0][14] ;
 wire \data_buffer[0][15] ;
 wire \data_buffer[0][16] ;
 wire \data_buffer[0][17] ;
 wire \data_buffer[0][18] ;
 wire \data_buffer[0][19] ;
 wire \data_buffer[0][1] ;
 wire \data_buffer[0][20] ;
 wire \data_buffer[0][21] ;
 wire \data_buffer[0][22] ;
 wire \data_buffer[0][23] ;
 wire \data_buffer[0][24] ;
 wire \data_buffer[0][25] ;
 wire \data_buffer[0][26] ;
 wire \data_buffer[0][27] ;
 wire \data_buffer[0][28] ;
 wire \data_buffer[0][29] ;
 wire \data_buffer[0][2] ;
 wire \data_buffer[0][30] ;
 wire \data_buffer[0][31] ;
 wire \data_buffer[0][3] ;
 wire \data_buffer[0][4] ;
 wire \data_buffer[0][5] ;
 wire \data_buffer[0][6] ;
 wire \data_buffer[0][7] ;
 wire \data_buffer[0][8] ;
 wire \data_buffer[0][9] ;
 wire \data_buffer[1][0] ;
 wire \data_buffer[1][10] ;
 wire \data_buffer[1][11] ;
 wire \data_buffer[1][12] ;
 wire \data_buffer[1][13] ;
 wire \data_buffer[1][14] ;
 wire \data_buffer[1][15] ;
 wire \data_buffer[1][16] ;
 wire \data_buffer[1][17] ;
 wire \data_buffer[1][18] ;
 wire \data_buffer[1][19] ;
 wire \data_buffer[1][1] ;
 wire \data_buffer[1][20] ;
 wire \data_buffer[1][21] ;
 wire \data_buffer[1][22] ;
 wire \data_buffer[1][23] ;
 wire \data_buffer[1][24] ;
 wire \data_buffer[1][25] ;
 wire \data_buffer[1][26] ;
 wire \data_buffer[1][27] ;
 wire \data_buffer[1][28] ;
 wire \data_buffer[1][29] ;
 wire \data_buffer[1][2] ;
 wire \data_buffer[1][30] ;
 wire \data_buffer[1][31] ;
 wire \data_buffer[1][3] ;
 wire \data_buffer[1][4] ;
 wire \data_buffer[1][5] ;
 wire \data_buffer[1][6] ;
 wire \data_buffer[1][7] ;
 wire \data_buffer[1][8] ;
 wire \data_buffer[1][9] ;
 wire \data_buffer[2][0] ;
 wire \data_buffer[2][10] ;
 wire \data_buffer[2][11] ;
 wire \data_buffer[2][12] ;
 wire \data_buffer[2][13] ;
 wire \data_buffer[2][14] ;
 wire \data_buffer[2][15] ;
 wire \data_buffer[2][16] ;
 wire \data_buffer[2][17] ;
 wire \data_buffer[2][18] ;
 wire \data_buffer[2][19] ;
 wire \data_buffer[2][1] ;
 wire \data_buffer[2][20] ;
 wire \data_buffer[2][21] ;
 wire \data_buffer[2][22] ;
 wire \data_buffer[2][23] ;
 wire \data_buffer[2][24] ;
 wire \data_buffer[2][25] ;
 wire \data_buffer[2][26] ;
 wire \data_buffer[2][27] ;
 wire \data_buffer[2][28] ;
 wire \data_buffer[2][29] ;
 wire \data_buffer[2][2] ;
 wire \data_buffer[2][30] ;
 wire \data_buffer[2][31] ;
 wire \data_buffer[2][3] ;
 wire \data_buffer[2][4] ;
 wire \data_buffer[2][5] ;
 wire \data_buffer[2][6] ;
 wire \data_buffer[2][7] ;
 wire \data_buffer[2][8] ;
 wire \data_buffer[2][9] ;
 wire \data_buffer[3][0] ;
 wire \data_buffer[3][10] ;
 wire \data_buffer[3][11] ;
 wire \data_buffer[3][12] ;
 wire \data_buffer[3][13] ;
 wire \data_buffer[3][14] ;
 wire \data_buffer[3][15] ;
 wire \data_buffer[3][16] ;
 wire \data_buffer[3][17] ;
 wire \data_buffer[3][18] ;
 wire \data_buffer[3][19] ;
 wire \data_buffer[3][1] ;
 wire \data_buffer[3][20] ;
 wire \data_buffer[3][21] ;
 wire \data_buffer[3][22] ;
 wire \data_buffer[3][23] ;
 wire \data_buffer[3][24] ;
 wire \data_buffer[3][25] ;
 wire \data_buffer[3][26] ;
 wire \data_buffer[3][27] ;
 wire \data_buffer[3][28] ;
 wire \data_buffer[3][29] ;
 wire \data_buffer[3][2] ;
 wire \data_buffer[3][30] ;
 wire \data_buffer[3][31] ;
 wire \data_buffer[3][3] ;
 wire \data_buffer[3][4] ;
 wire \data_buffer[3][5] ;
 wire \data_buffer[3][6] ;
 wire \data_buffer[3][7] ;
 wire \data_buffer[3][8] ;
 wire \data_buffer[3][9] ;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire clknet_leaf_10_clk;
 wire net1271;
 wire net957;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire net961;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire net964;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire net968;
 wire clknet_leaf_9_clk;
 wire net1274;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net1283;
 wire net1239;
 wire net1237;
 wire net1238;
 wire net1259;
 wire net1258;
 wire net1247;
 wire net1249;
 wire net1252;
 wire net1254;
 wire net1262;
 wire net1260;
 wire net1272;
 wire net1273;
 wire net1261;
 wire net1275;
 wire net1263;
 wire net1268;
 wire net1264;
 wire net1279;
 wire net1265;
 wire net1267;
 wire net1278;
 wire net1266;
 wire net1269;
 wire net1270;
 wire net1277;
 wire net1276;
 wire net1227;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire net1292;
 wire net1291;
 wire net1228;
 wire net1290;
 wire net1289;
 wire net1288;
 wire net1287;
 wire net1286;
 wire net1229;
 wire net1285;
 wire net1230;
 wire net1284;
 wire net1282;
 wire net1231;
 wire net1281;
 wire net1232;
 wire net1280;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1240;
 wire net1241;
 wire net1243;
 wire net1242;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1248;
 wire net1250;
 wire net1251;
 wire net1253;
 wire net1256;
 wire net1255;
 wire net1257;
 wire clknet_leaf_0_clk;
 wire net1293;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;

 sky130_fd_sc_hd__nor2_1 _3444_ (.A(net564),
    .B(net563),
    .Y(_1450_));
 sky130_fd_sc_hd__and2_1 _3445_ (.A(net562),
    .B(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input221 (.A(channel_length[64]),
    .X(net221));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input220 (.A(channel_length[63]),
    .X(net220));
 sky130_fd_sc_hd__nor2_1 _3448_ (.A(net556),
    .B(net555),
    .Y(_1453_));
 sky130_fd_sc_hd__and2_1 _3449_ (.A(net565),
    .B(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input219 (.A(channel_length[62]),
    .X(net219));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input218 (.A(channel_length[61]),
    .X(net218));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input217 (.A(channel_length[60]),
    .X(net217));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input216 (.A(channel_length[5]),
    .X(net216));
 sky130_fd_sc_hd__nand2b_1 _3454_ (.A_N(net557),
    .B(net554),
    .Y(_1458_));
 sky130_fd_sc_hd__nor2_4 _3455_ (.A(net558),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input215 (.A(channel_length[59]),
    .X(net215));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input214 (.A(channel_length[58]),
    .X(net214));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input213 (.A(channel_length[57]),
    .X(net213));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input212 (.A(channel_length[56]),
    .X(net212));
 sky130_fd_sc_hd__nor3b_2 _3460_ (.A(net1271),
    .B(net1272),
    .C_N(net1273),
    .Y(_1463_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input211 (.A(channel_length[55]),
    .X(net211));
 sky130_fd_sc_hd__nor2b_1 _3462_ (.A(net565),
    .B_N(net400),
    .Y(_1464_));
 sky130_fd_sc_hd__and3_1 _3463_ (.A(net132),
    .B(_1453_),
    .C(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input210 (.A(channel_length[54]),
    .X(net210));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input209 (.A(channel_length[53]),
    .X(net209));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input208 (.A(channel_length[52]),
    .X(net208));
 sky130_fd_sc_hd__nand2_1 _3467_ (.A(net126),
    .B(net1251),
    .Y(_1469_));
 sky130_fd_sc_hd__nand4bb_2 _3468_ (.A_N(net555),
    .B_N(net565),
    .C(net404),
    .D(net556),
    .Y(_1470_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input207 (.A(channel_length[51]),
    .X(net207));
 sky130_fd_sc_hd__nor2_1 _3470_ (.A(net267),
    .B(net1268),
    .Y(_1472_));
 sky130_fd_sc_hd__nand3_2 _3471_ (.A(net132),
    .B(_1453_),
    .C(_1464_),
    .Y(_1473_));
 sky130_fd_sc_hd__nor4bb_4 _3472_ (.A(net555),
    .B(net565),
    .C_N(net404),
    .D_N(net556),
    .Y(_1474_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input206 (.A(channel_length[50]),
    .X(net206));
 sky130_fd_sc_hd__nand2b_1 _3474_ (.A_N(net267),
    .B(net1267),
    .Y(_1476_));
 sky130_fd_sc_hd__nand2_1 _3475_ (.A(net1250),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__nand2_1 _3476_ (.A(\current_dst_addr[3][2] ),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__o21ai_0 _3477_ (.A1(\current_dst_addr[3][2] ),
    .A2(_1472_),
    .B1(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__nand2_1 _3478_ (.A(_1469_),
    .B(_1479_),
    .Y(_0122_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input205 (.A(channel_length[4]),
    .X(net205));
 sky130_fd_sc_hd__nand2_1 _3480_ (.A(net127),
    .B(net1251),
    .Y(_1481_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input204 (.A(channel_length[49]),
    .X(net204));
 sky130_fd_sc_hd__nand2_1 _3482_ (.A(\current_dst_addr[3][3] ),
    .B(net1250),
    .Y(_1483_));
 sky130_fd_sc_hd__nor2_1 _3483_ (.A(_0382_),
    .B(_1476_),
    .Y(_1484_));
 sky130_fd_sc_hd__a31oi_1 _3484_ (.A1(_1476_),
    .A2(_1481_),
    .A3(_1483_),
    .B1(_1484_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _3485_ (.A(\current_dst_addr[3][4] ),
    .Y(_1485_));
 sky130_fd_sc_hd__o21ai_0 _3486_ (.A1(_0381_),
    .A2(_1476_),
    .B1(_1477_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_1 _3487_ (.A(\current_dst_addr[3][4] ),
    .B(_0381_),
    .Y(_1487_));
 sky130_fd_sc_hd__or3_1 _3488_ (.A(net267),
    .B(net1268),
    .C(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__o21ai_0 _3489_ (.A1(net2),
    .A2(net1250),
    .B1(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__a21oi_1 _3490_ (.A1(_1485_),
    .A2(_1486_),
    .B1(_1489_),
    .Y(_0126_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input203 (.A(channel_length[48]),
    .X(net203));
 sky130_fd_sc_hd__nand3_1 _3492_ (.A(\current_dst_addr[3][2] ),
    .B(\current_dst_addr[3][3] ),
    .C(\current_dst_addr[3][4] ),
    .Y(_1491_));
 sky130_fd_sc_hd__nor2_1 _3493_ (.A(_1476_),
    .B(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_1 _3494_ (.A(_1472_),
    .B(_1491_),
    .Y(_1493_));
 sky130_fd_sc_hd__a21oi_1 _3495_ (.A1(_1477_),
    .A2(_1493_),
    .B1(\current_dst_addr[3][5] ),
    .Y(_1494_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input202 (.A(channel_length[47]),
    .X(net202));
 sky130_fd_sc_hd__nor2_1 _3497_ (.A(net3),
    .B(net1250),
    .Y(_1496_));
 sky130_fd_sc_hd__a211oi_1 _3498_ (.A1(\current_dst_addr[3][5] ),
    .A2(_1492_),
    .B1(_1494_),
    .C1(_1496_),
    .Y(_0127_));
 sky130_fd_sc_hd__nor2_1 _3499_ (.A(_1476_),
    .B(_1487_),
    .Y(_1497_));
 sky130_fd_sc_hd__nand3_1 _3500_ (.A(\current_dst_addr[3][4] ),
    .B(_0381_),
    .C(\current_dst_addr[3][5] ),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_1 _3501_ (.A(_1472_),
    .B(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__a21oi_1 _3502_ (.A1(_1477_),
    .A2(_1499_),
    .B1(\current_dst_addr[3][6] ),
    .Y(_1500_));
 sky130_fd_sc_hd__nor2_1 _3503_ (.A(net4),
    .B(net1250),
    .Y(_1501_));
 sky130_fd_sc_hd__a311oi_1 _3504_ (.A1(\current_dst_addr[3][5] ),
    .A2(\current_dst_addr[3][6] ),
    .A3(_1497_),
    .B1(_1500_),
    .C1(_1501_),
    .Y(_0128_));
 sky130_fd_sc_hd__a311oi_1 _3505_ (.A1(\current_dst_addr[3][5] ),
    .A2(\current_dst_addr[3][6] ),
    .A3(_1492_),
    .B1(net1251),
    .C1(\current_dst_addr[3][7] ),
    .Y(_1502_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input201 (.A(channel_length[46]),
    .X(net201));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input200 (.A(channel_length[45]),
    .X(net200));
 sky130_fd_sc_hd__or3_1 _3508_ (.A(net267),
    .B(net1268),
    .C(_1491_),
    .X(_1505_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input199 (.A(channel_length[44]),
    .X(net199));
 sky130_fd_sc_hd__nand3_1 _3510_ (.A(\current_dst_addr[3][5] ),
    .B(\current_dst_addr[3][6] ),
    .C(\current_dst_addr[3][7] ),
    .Y(_1507_));
 sky130_fd_sc_hd__o22ai_1 _3511_ (.A1(net5),
    .A2(net1250),
    .B1(_1505_),
    .B2(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__nor2_1 _3512_ (.A(_1502_),
    .B(_1508_),
    .Y(_0129_));
 sky130_fd_sc_hd__and3_1 _3513_ (.A(\current_dst_addr[3][5] ),
    .B(\current_dst_addr[3][6] ),
    .C(\current_dst_addr[3][7] ),
    .X(_1509_));
 sky130_fd_sc_hd__o21ai_0 _3514_ (.A1(_1487_),
    .A2(_1507_),
    .B1(_1472_),
    .Y(_1510_));
 sky130_fd_sc_hd__a21oi_1 _3515_ (.A1(_1477_),
    .A2(_1510_),
    .B1(\current_dst_addr[3][8] ),
    .Y(_1511_));
 sky130_fd_sc_hd__nor2_1 _3516_ (.A(net6),
    .B(net1250),
    .Y(_1512_));
 sky130_fd_sc_hd__a311oi_1 _3517_ (.A1(\current_dst_addr[3][8] ),
    .A2(_1497_),
    .A3(_1509_),
    .B1(_1511_),
    .C1(_1512_),
    .Y(_0130_));
 sky130_fd_sc_hd__and3_1 _3518_ (.A(\current_dst_addr[3][8] ),
    .B(\current_dst_addr[3][9] ),
    .C(_1509_),
    .X(_1513_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input198 (.A(channel_length[43]),
    .X(net198));
 sky130_fd_sc_hd__a311oi_1 _3520_ (.A1(\current_dst_addr[3][8] ),
    .A2(_1492_),
    .A3(_1509_),
    .B1(\current_dst_addr[3][9] ),
    .C1(net1251),
    .Y(_1515_));
 sky130_fd_sc_hd__nor2_1 _3521_ (.A(net7),
    .B(net1250),
    .Y(_1516_));
 sky130_fd_sc_hd__a211oi_1 _3522_ (.A1(_1492_),
    .A2(_1513_),
    .B1(_1515_),
    .C1(_1516_),
    .Y(_0131_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input197 (.A(channel_length[42]),
    .X(net197));
 sky130_fd_sc_hd__nor2_1 _3524_ (.A(net8),
    .B(net1250),
    .Y(_1518_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input196 (.A(channel_length[41]),
    .X(net196));
 sky130_fd_sc_hd__a211oi_1 _3526_ (.A1(_1497_),
    .A2(_1513_),
    .B1(\current_dst_addr[3][10] ),
    .C1(net1251),
    .Y(_1520_));
 sky130_fd_sc_hd__a311oi_1 _3527_ (.A1(\current_dst_addr[3][10] ),
    .A2(_1497_),
    .A3(_1513_),
    .B1(_1518_),
    .C1(_1520_),
    .Y(_0102_));
 sky130_fd_sc_hd__a311oi_1 _3528_ (.A1(\current_dst_addr[3][10] ),
    .A2(_1492_),
    .A3(_1513_),
    .B1(\current_dst_addr[3][11] ),
    .C1(net1251),
    .Y(_1521_));
 sky130_fd_sc_hd__and3_1 _3529_ (.A(\current_dst_addr[3][8] ),
    .B(\current_dst_addr[3][9] ),
    .C(\current_dst_addr[3][10] ),
    .X(_1522_));
 sky130_fd_sc_hd__nand3_1 _3530_ (.A(\current_dst_addr[3][11] ),
    .B(_1509_),
    .C(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__o22ai_1 _3531_ (.A1(net9),
    .A2(net1250),
    .B1(_1505_),
    .B2(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__nor2_1 _3532_ (.A(_1521_),
    .B(_1524_),
    .Y(_0103_));
 sky130_fd_sc_hd__nor2_1 _3533_ (.A(_1488_),
    .B(_1523_),
    .Y(_1525_));
 sky130_fd_sc_hd__nor3_1 _3534_ (.A(\current_dst_addr[3][12] ),
    .B(net1251),
    .C(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__nor2_1 _3535_ (.A(net10),
    .B(net1250),
    .Y(_1527_));
 sky130_fd_sc_hd__a211oi_1 _3536_ (.A1(\current_dst_addr[3][12] ),
    .A2(_1525_),
    .B1(_1526_),
    .C1(_1527_),
    .Y(_0104_));
 sky130_fd_sc_hd__and3_1 _3537_ (.A(\current_dst_addr[3][11] ),
    .B(_1509_),
    .C(_1522_),
    .X(_1528_));
 sky130_fd_sc_hd__a311oi_1 _3538_ (.A1(\current_dst_addr[3][12] ),
    .A2(_1492_),
    .A3(_1528_),
    .B1(\current_dst_addr[3][13] ),
    .C1(net1251),
    .Y(_1529_));
 sky130_fd_sc_hd__nand4_1 _3539_ (.A(\current_dst_addr[3][12] ),
    .B(\current_dst_addr[3][13] ),
    .C(_1492_),
    .D(_1528_),
    .Y(_1530_));
 sky130_fd_sc_hd__o21ai_0 _3540_ (.A1(net11),
    .A2(net1250),
    .B1(_1530_),
    .Y(_1531_));
 sky130_fd_sc_hd__nor2_1 _3541_ (.A(_1529_),
    .B(_1531_),
    .Y(_0105_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input195 (.A(channel_length[40]),
    .X(net195));
 sky130_fd_sc_hd__and3_1 _3543_ (.A(\current_dst_addr[3][11] ),
    .B(\current_dst_addr[3][12] ),
    .C(\current_dst_addr[3][13] ),
    .X(_1533_));
 sky130_fd_sc_hd__nand3_1 _3544_ (.A(_1509_),
    .B(_1522_),
    .C(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__nor2_1 _3545_ (.A(_1488_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__o21ai_0 _3546_ (.A1(_1487_),
    .A2(_1534_),
    .B1(_1472_),
    .Y(_1536_));
 sky130_fd_sc_hd__a21oi_1 _3547_ (.A1(_1477_),
    .A2(_1536_),
    .B1(\current_dst_addr[3][14] ),
    .Y(_1537_));
 sky130_fd_sc_hd__nor2_1 _3548_ (.A(net13),
    .B(net1250),
    .Y(_1538_));
 sky130_fd_sc_hd__a211oi_1 _3549_ (.A1(\current_dst_addr[3][14] ),
    .A2(_1535_),
    .B1(_1537_),
    .C1(_1538_),
    .Y(_0106_));
 sky130_fd_sc_hd__nor2_1 _3550_ (.A(_1505_),
    .B(_1534_),
    .Y(_1539_));
 sky130_fd_sc_hd__a211oi_1 _3551_ (.A1(\current_dst_addr[3][14] ),
    .A2(_1539_),
    .B1(net1251),
    .C1(\current_dst_addr[3][15] ),
    .Y(_1540_));
 sky130_fd_sc_hd__nor2_1 _3552_ (.A(net14),
    .B(net1250),
    .Y(_1541_));
 sky130_fd_sc_hd__a311oi_1 _3553_ (.A1(\current_dst_addr[3][14] ),
    .A2(\current_dst_addr[3][15] ),
    .A3(_1539_),
    .B1(_1540_),
    .C1(_1541_),
    .Y(_0107_));
 sky130_fd_sc_hd__a311oi_1 _3554_ (.A1(\current_dst_addr[3][14] ),
    .A2(\current_dst_addr[3][15] ),
    .A3(_1535_),
    .B1(net1251),
    .C1(\current_dst_addr[3][16] ),
    .Y(_1542_));
 sky130_fd_sc_hd__nand4_1 _3555_ (.A(\current_dst_addr[3][14] ),
    .B(\current_dst_addr[3][15] ),
    .C(\current_dst_addr[3][16] ),
    .D(_1535_),
    .Y(_1543_));
 sky130_fd_sc_hd__o21ai_0 _3556_ (.A1(net15),
    .A2(net1250),
    .B1(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__nor2_1 _3557_ (.A(_1542_),
    .B(_1544_),
    .Y(_0108_));
 sky130_fd_sc_hd__and4_1 _3558_ (.A(\current_dst_addr[3][14] ),
    .B(\current_dst_addr[3][15] ),
    .C(\current_dst_addr[3][16] ),
    .D(_1539_),
    .X(_1545_));
 sky130_fd_sc_hd__nor3_1 _3559_ (.A(\current_dst_addr[3][17] ),
    .B(net1251),
    .C(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__nor2_1 _3560_ (.A(net16),
    .B(net1250),
    .Y(_1547_));
 sky130_fd_sc_hd__a211oi_1 _3561_ (.A1(\current_dst_addr[3][17] ),
    .A2(_1545_),
    .B1(_1546_),
    .C1(_1547_),
    .Y(_0109_));
 sky130_fd_sc_hd__and4_1 _3562_ (.A(\current_dst_addr[3][14] ),
    .B(\current_dst_addr[3][15] ),
    .C(\current_dst_addr[3][16] ),
    .D(\current_dst_addr[3][17] ),
    .X(_1548_));
 sky130_fd_sc_hd__nand4_1 _3563_ (.A(\current_dst_addr[3][14] ),
    .B(\current_dst_addr[3][15] ),
    .C(\current_dst_addr[3][16] ),
    .D(\current_dst_addr[3][17] ),
    .Y(_1549_));
 sky130_fd_sc_hd__o31ai_1 _3564_ (.A1(_1487_),
    .A2(_1534_),
    .A3(_1549_),
    .B1(_1472_),
    .Y(_1550_));
 sky130_fd_sc_hd__a21oi_1 _3565_ (.A1(_1477_),
    .A2(_1550_),
    .B1(\current_dst_addr[3][18] ),
    .Y(_1551_));
 sky130_fd_sc_hd__nor2_1 _3566_ (.A(net17),
    .B(net1250),
    .Y(_1552_));
 sky130_fd_sc_hd__a311oi_1 _3567_ (.A1(\current_dst_addr[3][18] ),
    .A2(_1535_),
    .A3(_1548_),
    .B1(_1551_),
    .C1(_1552_),
    .Y(_0110_));
 sky130_fd_sc_hd__nor3_2 _3568_ (.A(_1505_),
    .B(_1534_),
    .C(_1549_),
    .Y(_1553_));
 sky130_fd_sc_hd__a211oi_1 _3569_ (.A1(\current_dst_addr[3][18] ),
    .A2(_1553_),
    .B1(net1251),
    .C1(\current_dst_addr[3][19] ),
    .Y(_1554_));
 sky130_fd_sc_hd__nor2_1 _3570_ (.A(net18),
    .B(net1250),
    .Y(_1555_));
 sky130_fd_sc_hd__a311oi_1 _3571_ (.A1(\current_dst_addr[3][18] ),
    .A2(\current_dst_addr[3][19] ),
    .A3(_1553_),
    .B1(_1554_),
    .C1(_1555_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_1 _3572_ (.A(\current_dst_addr[3][20] ),
    .Y(_1556_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input194 (.A(channel_length[3]),
    .X(net194));
 sky130_fd_sc_hd__nand4_1 _3574_ (.A(\current_dst_addr[3][18] ),
    .B(\current_dst_addr[3][19] ),
    .C(_1535_),
    .D(_1548_),
    .Y(_1558_));
 sky130_fd_sc_hd__o22ai_1 _3575_ (.A1(net19),
    .A2(net1250),
    .B1(_1558_),
    .B2(_1556_),
    .Y(_1559_));
 sky130_fd_sc_hd__a31oi_1 _3576_ (.A1(_1556_),
    .A2(net1250),
    .A3(_1558_),
    .B1(_1559_),
    .Y(_0112_));
 sky130_fd_sc_hd__nand4_1 _3577_ (.A(\current_dst_addr[3][18] ),
    .B(\current_dst_addr[3][19] ),
    .C(\current_dst_addr[3][20] ),
    .D(_1553_),
    .Y(_1560_));
 sky130_fd_sc_hd__nor2_1 _3578_ (.A(\current_dst_addr[3][21] ),
    .B(net1251),
    .Y(_1561_));
 sky130_fd_sc_hd__and4_1 _3579_ (.A(\current_dst_addr[3][18] ),
    .B(\current_dst_addr[3][19] ),
    .C(\current_dst_addr[3][20] ),
    .D(\current_dst_addr[3][21] ),
    .X(_1562_));
 sky130_fd_sc_hd__nand2_1 _3580_ (.A(_1553_),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__o21ai_0 _3581_ (.A1(net20),
    .A2(net1250),
    .B1(_1563_),
    .Y(_1564_));
 sky130_fd_sc_hd__a21oi_1 _3582_ (.A1(_1560_),
    .A2(_1561_),
    .B1(_1564_),
    .Y(_0113_));
 sky130_fd_sc_hd__a311oi_1 _3583_ (.A1(_1535_),
    .A2(_1548_),
    .A3(_1562_),
    .B1(net1251),
    .C1(\current_dst_addr[3][22] ),
    .Y(_1565_));
 sky130_fd_sc_hd__nand4_1 _3584_ (.A(\current_dst_addr[3][22] ),
    .B(_1535_),
    .C(_1548_),
    .D(_1562_),
    .Y(_1566_));
 sky130_fd_sc_hd__o21ai_0 _3585_ (.A1(net21),
    .A2(net1250),
    .B1(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__nor2_1 _3586_ (.A(_1565_),
    .B(_1567_),
    .Y(_0114_));
 sky130_fd_sc_hd__nand3_1 _3587_ (.A(\current_dst_addr[3][22] ),
    .B(_1548_),
    .C(_1562_),
    .Y(_1568_));
 sky130_fd_sc_hd__nor3_4 _3588_ (.A(_1505_),
    .B(_1534_),
    .C(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__nor3_1 _3589_ (.A(\current_dst_addr[3][23] ),
    .B(net1251),
    .C(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nor2_1 _3590_ (.A(_1534_),
    .B(_1568_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_1 _3591_ (.A(\current_dst_addr[3][23] ),
    .B(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__o22ai_1 _3592_ (.A1(net22),
    .A2(net1250),
    .B1(_1505_),
    .B2(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__nor2_1 _3593_ (.A(_1570_),
    .B(_1573_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand2_1 _3594_ (.A(\current_dst_addr[3][12] ),
    .B(\current_dst_addr[3][13] ),
    .Y(_1574_));
 sky130_fd_sc_hd__nor3_1 _3595_ (.A(_1523_),
    .B(_1574_),
    .C(_1568_),
    .Y(_1575_));
 sky130_fd_sc_hd__nand4_1 _3596_ (.A(\current_dst_addr[3][4] ),
    .B(_0381_),
    .C(\current_dst_addr[3][23] ),
    .D(_1575_),
    .Y(_1576_));
 sky130_fd_sc_hd__xor2_1 _3597_ (.A(\current_dst_addr[3][24] ),
    .B(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__o22ai_1 _3598_ (.A1(net24),
    .A2(net1250),
    .B1(_1477_),
    .B2(\current_dst_addr[3][24] ),
    .Y(_1578_));
 sky130_fd_sc_hd__a21oi_1 _3599_ (.A1(_1472_),
    .A2(_1577_),
    .B1(_1578_),
    .Y(_0116_));
 sky130_fd_sc_hd__a311oi_1 _3600_ (.A1(\current_dst_addr[3][23] ),
    .A2(\current_dst_addr[3][24] ),
    .A3(_1569_),
    .B1(net1251),
    .C1(\current_dst_addr[3][25] ),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_1 _3601_ (.A(_1492_),
    .B(_1571_),
    .Y(_1580_));
 sky130_fd_sc_hd__nand3_1 _3602_ (.A(\current_dst_addr[3][23] ),
    .B(\current_dst_addr[3][24] ),
    .C(\current_dst_addr[3][25] ),
    .Y(_1581_));
 sky130_fd_sc_hd__o22ai_1 _3603_ (.A1(net25),
    .A2(net1250),
    .B1(_1580_),
    .B2(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__nor2_1 _3604_ (.A(_1579_),
    .B(_1582_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_1 _3605_ (.A(\current_dst_addr[3][26] ),
    .Y(_1583_));
 sky130_fd_sc_hd__nor3_2 _3606_ (.A(_1488_),
    .B(_1534_),
    .C(_1568_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand2b_1 _3607_ (.A_N(_1581_),
    .B(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__o22ai_1 _3608_ (.A1(net26),
    .A2(net1250),
    .B1(_1585_),
    .B2(_1583_),
    .Y(_1586_));
 sky130_fd_sc_hd__a31oi_1 _3609_ (.A1(_1583_),
    .A2(net1250),
    .A3(_1585_),
    .B1(_1586_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_1 _3610_ (.A(_1583_),
    .B(_1581_),
    .Y(_1587_));
 sky130_fd_sc_hd__nor2_1 _3611_ (.A(net27),
    .B(net1250),
    .Y(_1588_));
 sky130_fd_sc_hd__a211oi_1 _3612_ (.A1(_1569_),
    .A2(_1587_),
    .B1(\current_dst_addr[3][27] ),
    .C1(net1251),
    .Y(_1589_));
 sky130_fd_sc_hd__a311oi_1 _3613_ (.A1(\current_dst_addr[3][27] ),
    .A2(_1569_),
    .A3(_1587_),
    .B1(_1588_),
    .C1(_1589_),
    .Y(_0119_));
 sky130_fd_sc_hd__and3_1 _3614_ (.A(\current_dst_addr[3][27] ),
    .B(\current_dst_addr[3][28] ),
    .C(_1587_),
    .X(_1590_));
 sky130_fd_sc_hd__a311oi_1 _3615_ (.A1(\current_dst_addr[3][27] ),
    .A2(_1584_),
    .A3(_1587_),
    .B1(\current_dst_addr[3][28] ),
    .C1(net1251),
    .Y(_1591_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input193 (.A(channel_length[39]),
    .X(net193));
 sky130_fd_sc_hd__nor2_1 _3617_ (.A(net28),
    .B(net1250),
    .Y(_1593_));
 sky130_fd_sc_hd__a211oi_1 _3618_ (.A1(_1584_),
    .A2(_1590_),
    .B1(_1591_),
    .C1(_1593_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand2_1 _3619_ (.A(\current_dst_addr[3][29] ),
    .B(net1250),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_1 _3620_ (.A(_1569_),
    .B(_1590_),
    .Y(_1595_));
 sky130_fd_sc_hd__mux2i_1 _3621_ (.A0(\current_dst_addr[3][29] ),
    .A1(_1594_),
    .S(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__a21o_1 _3622_ (.A1(net29),
    .A2(net1251),
    .B1(_1596_),
    .X(_0121_));
 sky130_fd_sc_hd__a311oi_1 _3623_ (.A1(\current_dst_addr[3][29] ),
    .A2(_1584_),
    .A3(_1590_),
    .B1(\current_dst_addr[3][30] ),
    .C1(net1251),
    .Y(_1597_));
 sky130_fd_sc_hd__nand4_1 _3624_ (.A(\current_dst_addr[3][29] ),
    .B(\current_dst_addr[3][30] ),
    .C(_1584_),
    .D(_1590_),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_0 _3625_ (.A1(net30),
    .A2(net1250),
    .B1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_1597_),
    .B(_1599_),
    .Y(_0123_));
 sky130_fd_sc_hd__nand4_1 _3627_ (.A(\current_dst_addr[3][29] ),
    .B(\current_dst_addr[3][30] ),
    .C(_1569_),
    .D(_1590_),
    .Y(_1600_));
 sky130_fd_sc_hd__nand3_1 _3628_ (.A(\current_dst_addr[3][31] ),
    .B(net1250),
    .C(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__nand2_1 _3629_ (.A(net31),
    .B(net1251),
    .Y(_1602_));
 sky130_fd_sc_hd__o211ai_1 _3630_ (.A1(\current_dst_addr[3][31] ),
    .A2(_1600_),
    .B1(_1601_),
    .C1(_1602_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor2b_1 _3631_ (.A(net562),
    .B_N(net399),
    .Y(_1603_));
 sky130_fd_sc_hd__and3_2 _3632_ (.A(net131),
    .B(_1450_),
    .C(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input192 (.A(channel_length[38]),
    .X(net192));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input191 (.A(channel_length[37]),
    .X(net191));
 sky130_fd_sc_hd__nand4bb_4 _3635_ (.A_N(net563),
    .B_N(net562),
    .C(net403),
    .D(net564),
    .Y(_1607_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input190 (.A(channel_length[36]),
    .X(net190));
 sky130_fd_sc_hd__nor2_1 _3637_ (.A(net265),
    .B(net1266),
    .Y(_1609_));
 sky130_fd_sc_hd__nor2_1 _3638_ (.A(_1604_),
    .B(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__and4bb_2 _3639_ (.A_N(net563),
    .B_N(net562),
    .C(net403),
    .D(net564),
    .X(_1611_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input189 (.A(channel_length[35]),
    .X(net189));
 sky130_fd_sc_hd__nand2b_1 _3641_ (.A_N(net265),
    .B(_1611_),
    .Y(_1613_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input188 (.A(channel_length[34]),
    .X(net188));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(\current_dst_addr[2][2] ),
    .B(_1613_),
    .Y(_1615_));
 sky130_fd_sc_hd__a221o_1 _3644_ (.A1(net91),
    .A2(_1604_),
    .B1(_1610_),
    .B2(\current_dst_addr[2][2] ),
    .C1(_1615_),
    .X(_0092_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input187 (.A(channel_length[33]),
    .X(net187));
 sky130_fd_sc_hd__nand2_1 _3646_ (.A(net92),
    .B(_1604_),
    .Y(_1617_));
 sky130_fd_sc_hd__nand3_4 _3647_ (.A(net131),
    .B(_1450_),
    .C(_1603_),
    .Y(_1618_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input186 (.A(channel_length[32]),
    .X(net186));
 sky130_fd_sc_hd__nand2_1 _3649_ (.A(\current_dst_addr[2][3] ),
    .B(net1248),
    .Y(_1620_));
 sky130_fd_sc_hd__nor2_1 _3650_ (.A(_0384_),
    .B(_1613_),
    .Y(_1621_));
 sky130_fd_sc_hd__a31oi_1 _3651_ (.A1(_1613_),
    .A2(_1617_),
    .A3(_1620_),
    .B1(_1621_),
    .Y(_0095_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input185 (.A(channel_length[31]),
    .X(net185));
 sky130_fd_sc_hd__nand2_1 _3653_ (.A(net1248),
    .B(_1613_),
    .Y(_1623_));
 sky130_fd_sc_hd__or3_1 _3654_ (.A(net265),
    .B(_0383_),
    .C(net1266),
    .X(_1624_));
 sky130_fd_sc_hd__a21oi_1 _3655_ (.A1(_1623_),
    .A2(_1624_),
    .B1(\current_dst_addr[2][4] ),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _3656_ (.A(\current_dst_addr[2][4] ),
    .B(_0383_),
    .Y(_1626_));
 sky130_fd_sc_hd__nor3_2 _3657_ (.A(net265),
    .B(_1607_),
    .C(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input184 (.A(channel_length[30]),
    .X(net184));
 sky130_fd_sc_hd__nor2_1 _3659_ (.A(net93),
    .B(net1248),
    .Y(_1629_));
 sky130_fd_sc_hd__nor3_1 _3660_ (.A(_1625_),
    .B(_1627_),
    .C(_1629_),
    .Y(_0096_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input183 (.A(channel_length[2]),
    .X(net183));
 sky130_fd_sc_hd__nand3_1 _3662_ (.A(\current_dst_addr[2][2] ),
    .B(\current_dst_addr[2][3] ),
    .C(\current_dst_addr[2][4] ),
    .Y(_1631_));
 sky130_fd_sc_hd__a21oi_1 _3663_ (.A1(_1609_),
    .A2(_1631_),
    .B1(_1610_),
    .Y(_1632_));
 sky130_fd_sc_hd__nor2_1 _3664_ (.A(_1613_),
    .B(_1631_),
    .Y(_1633_));
 sky130_fd_sc_hd__nand2_1 _3665_ (.A(\current_dst_addr[2][5] ),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__o221a_2 _3666_ (.A1(net94),
    .A2(net1248),
    .B1(_1632_),
    .B2(\current_dst_addr[2][5] ),
    .C1(_1634_),
    .X(_0097_));
 sky130_fd_sc_hd__nor2_1 _3667_ (.A(net96),
    .B(net1248),
    .Y(_1635_));
 sky130_fd_sc_hd__nand3_1 _3668_ (.A(\current_dst_addr[2][4] ),
    .B(_0383_),
    .C(\current_dst_addr[2][5] ),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _3669_ (.A(_1609_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__a21oi_1 _3670_ (.A1(_1623_),
    .A2(_1637_),
    .B1(\current_dst_addr[2][6] ),
    .Y(_1638_));
 sky130_fd_sc_hd__a311oi_1 _3671_ (.A1(\current_dst_addr[2][5] ),
    .A2(\current_dst_addr[2][6] ),
    .A3(_1627_),
    .B1(_1635_),
    .C1(_1638_),
    .Y(_0098_));
 sky130_fd_sc_hd__and3_1 _3672_ (.A(\current_dst_addr[2][5] ),
    .B(\current_dst_addr[2][6] ),
    .C(\current_dst_addr[2][7] ),
    .X(_1639_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input182 (.A(channel_length[29]),
    .X(net182));
 sky130_fd_sc_hd__a311oi_1 _3674_ (.A1(\current_dst_addr[2][5] ),
    .A2(\current_dst_addr[2][6] ),
    .A3(_1633_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][7] ),
    .Y(_1641_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input181 (.A(channel_length[28]),
    .X(net181));
 sky130_fd_sc_hd__nor2_1 _3676_ (.A(net97),
    .B(net1248),
    .Y(_1643_));
 sky130_fd_sc_hd__a211oi_1 _3677_ (.A1(_1633_),
    .A2(_1639_),
    .B1(_1641_),
    .C1(_1643_),
    .Y(_0099_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input180 (.A(channel_length[27]),
    .X(net180));
 sky130_fd_sc_hd__a211oi_1 _3679_ (.A1(_1627_),
    .A2(_1639_),
    .B1(\current_dst_addr[2][8] ),
    .C1(_1604_),
    .Y(_1645_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input179 (.A(channel_length[26]),
    .X(net179));
 sky130_fd_sc_hd__nor2_1 _3681_ (.A(net98),
    .B(net1248),
    .Y(_1647_));
 sky130_fd_sc_hd__a311oi_1 _3682_ (.A1(\current_dst_addr[2][8] ),
    .A2(_1627_),
    .A3(_1639_),
    .B1(_1645_),
    .C1(_1647_),
    .Y(_0100_));
 sky130_fd_sc_hd__and3_1 _3683_ (.A(\current_dst_addr[2][2] ),
    .B(\current_dst_addr[2][3] ),
    .C(\current_dst_addr[2][4] ),
    .X(_1648_));
 sky130_fd_sc_hd__nand3_1 _3684_ (.A(\current_dst_addr[2][8] ),
    .B(_1648_),
    .C(_1639_),
    .Y(_1649_));
 sky130_fd_sc_hd__a21oi_1 _3685_ (.A1(_1609_),
    .A2(_1649_),
    .B1(_1610_),
    .Y(_1650_));
 sky130_fd_sc_hd__and3_1 _3686_ (.A(\current_dst_addr[2][8] ),
    .B(\current_dst_addr[2][9] ),
    .C(_1639_),
    .X(_1651_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input178 (.A(channel_length[25]),
    .X(net178));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(_1633_),
    .B(_1651_),
    .Y(_1653_));
 sky130_fd_sc_hd__o221a_2 _3689_ (.A1(net99),
    .A2(net1248),
    .B1(_1650_),
    .B2(\current_dst_addr[2][9] ),
    .C1(_1653_),
    .X(_0101_));
 sky130_fd_sc_hd__nand3_1 _3690_ (.A(\current_dst_addr[2][4] ),
    .B(_0383_),
    .C(_1651_),
    .Y(_1654_));
 sky130_fd_sc_hd__a21oi_1 _3691_ (.A1(_1609_),
    .A2(_1654_),
    .B1(_1610_),
    .Y(_1655_));
 sky130_fd_sc_hd__and2_1 _3692_ (.A(_1627_),
    .B(_1651_),
    .X(_1656_));
 sky130_fd_sc_hd__nand2_1 _3693_ (.A(\current_dst_addr[2][10] ),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__o221a_2 _3694_ (.A1(net100),
    .A2(net1248),
    .B1(_1655_),
    .B2(\current_dst_addr[2][10] ),
    .C1(_1657_),
    .X(_0072_));
 sky130_fd_sc_hd__nand3_1 _3695_ (.A(\current_dst_addr[2][10] ),
    .B(_1648_),
    .C(_1651_),
    .Y(_1658_));
 sky130_fd_sc_hd__a21oi_1 _3696_ (.A1(_1609_),
    .A2(_1658_),
    .B1(_1610_),
    .Y(_1659_));
 sky130_fd_sc_hd__nor2_1 _3697_ (.A(\current_dst_addr[2][11] ),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _3698_ (.A(\current_dst_addr[2][10] ),
    .B(\current_dst_addr[2][11] ),
    .Y(_1661_));
 sky130_fd_sc_hd__o22ai_1 _3699_ (.A1(net101),
    .A2(net1248),
    .B1(_1653_),
    .B2(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__nor2_1 _3700_ (.A(_1660_),
    .B(_1662_),
    .Y(_0073_));
 sky130_fd_sc_hd__nor2_1 _3701_ (.A(net102),
    .B(net1248),
    .Y(_1663_));
 sky130_fd_sc_hd__a311oi_1 _3702_ (.A1(\current_dst_addr[2][10] ),
    .A2(\current_dst_addr[2][11] ),
    .A3(_1656_),
    .B1(net1249),
    .C1(\current_dst_addr[2][12] ),
    .Y(_1664_));
 sky130_fd_sc_hd__and4_1 _3703_ (.A(\current_dst_addr[2][10] ),
    .B(\current_dst_addr[2][11] ),
    .C(\current_dst_addr[2][12] ),
    .D(_1656_),
    .X(_1665_));
 sky130_fd_sc_hd__nor3_1 _3704_ (.A(_1663_),
    .B(_1664_),
    .C(_1665_),
    .Y(_0074_));
 sky130_fd_sc_hd__and3_1 _3705_ (.A(\current_dst_addr[2][10] ),
    .B(\current_dst_addr[2][11] ),
    .C(\current_dst_addr[2][12] ),
    .X(_1666_));
 sky130_fd_sc_hd__a311oi_1 _3706_ (.A1(_1633_),
    .A2(_1651_),
    .A3(_1666_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][13] ),
    .Y(_1667_));
 sky130_fd_sc_hd__and2_1 _3707_ (.A(\current_dst_addr[2][13] ),
    .B(_1666_),
    .X(_1668_));
 sky130_fd_sc_hd__nand3_1 _3708_ (.A(_1633_),
    .B(_1651_),
    .C(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__o21ai_0 _3709_ (.A1(net103),
    .A2(net1248),
    .B1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__nor2_1 _3710_ (.A(_1667_),
    .B(_1670_),
    .Y(_0075_));
 sky130_fd_sc_hd__nor2_1 _3711_ (.A(net104),
    .B(net1248),
    .Y(_1671_));
 sky130_fd_sc_hd__a211oi_1 _3712_ (.A1(_1656_),
    .A2(_1668_),
    .B1(\current_dst_addr[2][14] ),
    .C1(net1249),
    .Y(_1672_));
 sky130_fd_sc_hd__a311oi_1 _3713_ (.A1(\current_dst_addr[2][14] ),
    .A2(_1656_),
    .A3(_1668_),
    .B1(_1671_),
    .C1(_1672_),
    .Y(_0076_));
 sky130_fd_sc_hd__and3_1 _3714_ (.A(\current_dst_addr[2][13] ),
    .B(\current_dst_addr[2][14] ),
    .C(_1666_),
    .X(_1673_));
 sky130_fd_sc_hd__nand3_1 _3715_ (.A(_1648_),
    .B(_1651_),
    .C(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__nor2_1 _3716_ (.A(_1613_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__a21oi_1 _3717_ (.A1(_1609_),
    .A2(_1674_),
    .B1(_1610_),
    .Y(_1676_));
 sky130_fd_sc_hd__nor2_1 _3718_ (.A(\current_dst_addr[2][15] ),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input177 (.A(channel_length[24]),
    .X(net177));
 sky130_fd_sc_hd__nor2_1 _3720_ (.A(net105),
    .B(net1248),
    .Y(_1679_));
 sky130_fd_sc_hd__a211oi_1 _3721_ (.A1(\current_dst_addr[2][15] ),
    .A2(_1675_),
    .B1(_1677_),
    .C1(_1679_),
    .Y(_0077_));
 sky130_fd_sc_hd__and3_1 _3722_ (.A(_1627_),
    .B(_1651_),
    .C(_1673_),
    .X(_1680_));
 sky130_fd_sc_hd__a211oi_1 _3723_ (.A1(\current_dst_addr[2][15] ),
    .A2(_1680_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][16] ),
    .Y(_1681_));
 sky130_fd_sc_hd__nor2_1 _3724_ (.A(net107),
    .B(net1248),
    .Y(_1682_));
 sky130_fd_sc_hd__a311oi_1 _3725_ (.A1(\current_dst_addr[2][15] ),
    .A2(\current_dst_addr[2][16] ),
    .A3(_1680_),
    .B1(_1681_),
    .C1(_1682_),
    .Y(_0078_));
 sky130_fd_sc_hd__and3_1 _3726_ (.A(\current_dst_addr[2][15] ),
    .B(\current_dst_addr[2][16] ),
    .C(\current_dst_addr[2][17] ),
    .X(_1683_));
 sky130_fd_sc_hd__a311oi_1 _3727_ (.A1(\current_dst_addr[2][15] ),
    .A2(\current_dst_addr[2][16] ),
    .A3(_1675_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][17] ),
    .Y(_1684_));
 sky130_fd_sc_hd__nor2_1 _3728_ (.A(net108),
    .B(net1248),
    .Y(_1685_));
 sky130_fd_sc_hd__a211oi_1 _3729_ (.A1(_1675_),
    .A2(_1683_),
    .B1(_1684_),
    .C1(_1685_),
    .Y(_0079_));
 sky130_fd_sc_hd__nor2_1 _3730_ (.A(net109),
    .B(net1248),
    .Y(_1686_));
 sky130_fd_sc_hd__a211oi_1 _3731_ (.A1(_1680_),
    .A2(_1683_),
    .B1(\current_dst_addr[2][18] ),
    .C1(_1604_),
    .Y(_1687_));
 sky130_fd_sc_hd__and3_1 _3732_ (.A(\current_dst_addr[2][18] ),
    .B(_1680_),
    .C(_1683_),
    .X(_1688_));
 sky130_fd_sc_hd__nor3_1 _3733_ (.A(_1686_),
    .B(_1687_),
    .C(_1688_),
    .Y(_0080_));
 sky130_fd_sc_hd__and3_1 _3734_ (.A(\current_dst_addr[2][18] ),
    .B(\current_dst_addr[2][19] ),
    .C(_1683_),
    .X(_1689_));
 sky130_fd_sc_hd__a311oi_1 _3735_ (.A1(\current_dst_addr[2][18] ),
    .A2(_1675_),
    .A3(_1683_),
    .B1(\current_dst_addr[2][19] ),
    .C1(_1604_),
    .Y(_1690_));
 sky130_fd_sc_hd__nor2_1 _3736_ (.A(net110),
    .B(net1248),
    .Y(_1691_));
 sky130_fd_sc_hd__a211oi_1 _3737_ (.A1(_1675_),
    .A2(_1689_),
    .B1(_1690_),
    .C1(_1691_),
    .Y(_0081_));
 sky130_fd_sc_hd__nor2_1 _3738_ (.A(net111),
    .B(net1248),
    .Y(_1692_));
 sky130_fd_sc_hd__a211oi_1 _3739_ (.A1(\current_dst_addr[2][19] ),
    .A2(_1688_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][20] ),
    .Y(_1693_));
 sky130_fd_sc_hd__a311oi_1 _3740_ (.A1(\current_dst_addr[2][19] ),
    .A2(\current_dst_addr[2][20] ),
    .A3(_1688_),
    .B1(_1692_),
    .C1(_1693_),
    .Y(_0082_));
 sky130_fd_sc_hd__a311oi_1 _3741_ (.A1(\current_dst_addr[2][20] ),
    .A2(_1675_),
    .A3(_1689_),
    .B1(\current_dst_addr[2][21] ),
    .C1(_1604_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand3_1 _3742_ (.A(\current_dst_addr[2][20] ),
    .B(\current_dst_addr[2][21] ),
    .C(_1689_),
    .Y(_1695_));
 sky130_fd_sc_hd__o32ai_1 _3743_ (.A1(_1613_),
    .A2(_1674_),
    .A3(_1695_),
    .B1(net1248),
    .B2(net112),
    .Y(_1696_));
 sky130_fd_sc_hd__nor2_1 _3744_ (.A(_1694_),
    .B(_1696_),
    .Y(_0083_));
 sky130_fd_sc_hd__nand3_1 _3745_ (.A(_1627_),
    .B(_1651_),
    .C(_1673_),
    .Y(_1697_));
 sky130_fd_sc_hd__nor2_1 _3746_ (.A(_1697_),
    .B(_1695_),
    .Y(_1698_));
 sky130_fd_sc_hd__nor3_1 _3747_ (.A(\current_dst_addr[2][22] ),
    .B(net1249),
    .C(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_1 _3748_ (.A(net113),
    .B(net1248),
    .Y(_1700_));
 sky130_fd_sc_hd__a211oi_1 _3749_ (.A1(\current_dst_addr[2][22] ),
    .A2(_1698_),
    .B1(_1699_),
    .C1(_1700_),
    .Y(_0084_));
 sky130_fd_sc_hd__nand4_1 _3750_ (.A(\current_dst_addr[2][20] ),
    .B(\current_dst_addr[2][21] ),
    .C(\current_dst_addr[2][22] ),
    .D(_1689_),
    .Y(_1701_));
 sky130_fd_sc_hd__nor3_2 _3751_ (.A(_1613_),
    .B(_1674_),
    .C(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__nor3_1 _3752_ (.A(\current_dst_addr[2][23] ),
    .B(_1604_),
    .C(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__nor2_1 _3753_ (.A(net114),
    .B(net1248),
    .Y(_1704_));
 sky130_fd_sc_hd__a211oi_1 _3754_ (.A1(\current_dst_addr[2][23] ),
    .A2(_1702_),
    .B1(_1703_),
    .C1(_1704_),
    .Y(_0085_));
 sky130_fd_sc_hd__nor2_1 _3755_ (.A(net115),
    .B(net1248),
    .Y(_1705_));
 sky130_fd_sc_hd__nor2_1 _3756_ (.A(_1697_),
    .B(_1701_),
    .Y(_1706_));
 sky130_fd_sc_hd__a211oi_1 _3757_ (.A1(\current_dst_addr[2][23] ),
    .A2(_1706_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][24] ),
    .Y(_1707_));
 sky130_fd_sc_hd__and3_1 _3758_ (.A(\current_dst_addr[2][23] ),
    .B(\current_dst_addr[2][24] ),
    .C(_1706_),
    .X(_1708_));
 sky130_fd_sc_hd__nor3_1 _3759_ (.A(_1705_),
    .B(_1707_),
    .C(_1708_),
    .Y(_0086_));
 sky130_fd_sc_hd__and3_1 _3760_ (.A(\current_dst_addr[2][23] ),
    .B(\current_dst_addr[2][24] ),
    .C(\current_dst_addr[2][25] ),
    .X(_1709_));
 sky130_fd_sc_hd__a311oi_1 _3761_ (.A1(\current_dst_addr[2][23] ),
    .A2(\current_dst_addr[2][24] ),
    .A3(_1702_),
    .B1(_1604_),
    .C1(\current_dst_addr[2][25] ),
    .Y(_1710_));
 sky130_fd_sc_hd__nor2_1 _3762_ (.A(net116),
    .B(net1248),
    .Y(_1711_));
 sky130_fd_sc_hd__a211oi_1 _3763_ (.A1(_1702_),
    .A2(_1709_),
    .B1(_1710_),
    .C1(_1711_),
    .Y(_0087_));
 sky130_fd_sc_hd__and4_1 _3764_ (.A(\current_dst_addr[2][23] ),
    .B(\current_dst_addr[2][24] ),
    .C(\current_dst_addr[2][25] ),
    .D(\current_dst_addr[2][26] ),
    .X(_1712_));
 sky130_fd_sc_hd__a211oi_1 _3765_ (.A1(_1706_),
    .A2(_1709_),
    .B1(\current_dst_addr[2][26] ),
    .C1(_1604_),
    .Y(_1713_));
 sky130_fd_sc_hd__nor2_1 _3766_ (.A(net118),
    .B(net1248),
    .Y(_1714_));
 sky130_fd_sc_hd__a211oi_1 _3767_ (.A1(_1706_),
    .A2(_1712_),
    .B1(_1713_),
    .C1(_1714_),
    .Y(_0088_));
 sky130_fd_sc_hd__and2_1 _3768_ (.A(\current_dst_addr[2][27] ),
    .B(_1712_),
    .X(_1715_));
 sky130_fd_sc_hd__a211oi_1 _3769_ (.A1(_1702_),
    .A2(_1712_),
    .B1(\current_dst_addr[2][27] ),
    .C1(_1604_),
    .Y(_1716_));
 sky130_fd_sc_hd__nor2_1 _3770_ (.A(net119),
    .B(net1248),
    .Y(_1717_));
 sky130_fd_sc_hd__a211oi_1 _3771_ (.A1(_1702_),
    .A2(_1715_),
    .B1(_1716_),
    .C1(_1717_),
    .Y(_0089_));
 sky130_fd_sc_hd__nor2_1 _3772_ (.A(net120),
    .B(net1248),
    .Y(_1718_));
 sky130_fd_sc_hd__a211oi_1 _3773_ (.A1(_1706_),
    .A2(_1715_),
    .B1(\current_dst_addr[2][28] ),
    .C1(_1604_),
    .Y(_1719_));
 sky130_fd_sc_hd__a311oi_1 _3774_ (.A1(\current_dst_addr[2][28] ),
    .A2(_1706_),
    .A3(_1715_),
    .B1(_1718_),
    .C1(_1719_),
    .Y(_0090_));
 sky130_fd_sc_hd__and4_1 _3775_ (.A(\current_dst_addr[2][27] ),
    .B(\current_dst_addr[2][28] ),
    .C(\current_dst_addr[2][29] ),
    .D(_1712_),
    .X(_1720_));
 sky130_fd_sc_hd__a311oi_1 _3776_ (.A1(\current_dst_addr[2][28] ),
    .A2(_1702_),
    .A3(_1715_),
    .B1(\current_dst_addr[2][29] ),
    .C1(_1604_),
    .Y(_1721_));
 sky130_fd_sc_hd__nor2_1 _3777_ (.A(net121),
    .B(net1248),
    .Y(_1722_));
 sky130_fd_sc_hd__a211oi_1 _3778_ (.A1(_1702_),
    .A2(_1720_),
    .B1(_1721_),
    .C1(_1722_),
    .Y(_0091_));
 sky130_fd_sc_hd__nor2_1 _3779_ (.A(net122),
    .B(net1248),
    .Y(_1723_));
 sky130_fd_sc_hd__a211oi_1 _3780_ (.A1(_1706_),
    .A2(_1720_),
    .B1(\current_dst_addr[2][30] ),
    .C1(_1604_),
    .Y(_1724_));
 sky130_fd_sc_hd__a311oi_1 _3781_ (.A1(\current_dst_addr[2][30] ),
    .A2(_1706_),
    .A3(_1720_),
    .B1(_1723_),
    .C1(_1724_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_1 _3782_ (.A(\current_dst_addr[2][31] ),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _3783_ (.A(\current_dst_addr[2][30] ),
    .B(_1720_),
    .Y(_1726_));
 sky130_fd_sc_hd__nor3_1 _3784_ (.A(_1674_),
    .B(_1701_),
    .C(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__o21ai_0 _3785_ (.A1(_1613_),
    .A2(_1727_),
    .B1(_1623_),
    .Y(_1728_));
 sky130_fd_sc_hd__nor2_1 _3786_ (.A(net123),
    .B(net1248),
    .Y(_1729_));
 sky130_fd_sc_hd__a31oi_1 _3787_ (.A1(\current_dst_addr[2][31] ),
    .A2(_1609_),
    .A3(_1727_),
    .B1(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__a21boi_0 _3788_ (.A1(_1725_),
    .A2(_1728_),
    .B1_N(_1730_),
    .Y(_0094_));
 sky130_fd_sc_hd__nor2b_1 _3789_ (.A(net1272),
    .B_N(net398),
    .Y(_1731_));
 sky130_fd_sc_hd__nor2_1 _3790_ (.A(net1271),
    .B(net1273),
    .Y(_1732_));
 sky130_fd_sc_hd__and3_2 _3791_ (.A(net130),
    .B(_1731_),
    .C(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input176 (.A(channel_length[23]),
    .X(net176));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input175 (.A(channel_length[22]),
    .X(net175));
 sky130_fd_sc_hd__nand4bb_2 _3794_ (.A_N(net1273),
    .B_N(net1272),
    .C(net1293),
    .D(net1271),
    .Y(_1736_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input174 (.A(channel_length[21]),
    .X(net174));
 sky130_fd_sc_hd__nor2_1 _3796_ (.A(net263),
    .B(_1736_),
    .Y(_1738_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input173 (.A(channel_length[20]),
    .X(net173));
 sky130_fd_sc_hd__nor2_1 _3798_ (.A(net1247),
    .B(_1738_),
    .Y(_1740_));
 sky130_fd_sc_hd__nor4bb_4 _3799_ (.A(net1273),
    .B(net1272),
    .C_N(net1293),
    .D_N(net561),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2b_1 _3800_ (.A_N(net263),
    .B(net1264),
    .Y(_1742_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input172 (.A(channel_length[1]),
    .X(net172));
 sky130_fd_sc_hd__nor2_1 _3802_ (.A(\current_dst_addr[1][2] ),
    .B(_1742_),
    .Y(_1744_));
 sky130_fd_sc_hd__a221o_1 _3803_ (.A1(net56),
    .A2(net1246),
    .B1(_1740_),
    .B2(\current_dst_addr[1][2] ),
    .C1(_1744_),
    .X(_0062_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input171 (.A(channel_length[19]),
    .X(net171));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input170 (.A(channel_length[18]),
    .X(net170));
 sky130_fd_sc_hd__nand2_1 _3806_ (.A(net57),
    .B(net1247),
    .Y(_1747_));
 sky130_fd_sc_hd__nand3_4 _3807_ (.A(net130),
    .B(_1731_),
    .C(_1732_),
    .Y(_1748_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input169 (.A(channel_length[17]),
    .X(net169));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input168 (.A(channel_length[16]),
    .X(net168));
 sky130_fd_sc_hd__nand2_1 _3810_ (.A(\current_dst_addr[1][3] ),
    .B(net1245),
    .Y(_1751_));
 sky130_fd_sc_hd__nor2_1 _3811_ (.A(_0386_),
    .B(_1742_),
    .Y(_1752_));
 sky130_fd_sc_hd__a31oi_1 _3812_ (.A1(_1742_),
    .A2(_1747_),
    .A3(_1751_),
    .B1(_1752_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_1 _3813_ (.A(\current_dst_addr[1][4] ),
    .Y(_1753_));
 sky130_fd_sc_hd__nand2_1 _3814_ (.A(_1748_),
    .B(_1742_),
    .Y(_1754_));
 sky130_fd_sc_hd__o21ai_0 _3815_ (.A1(_0385_),
    .A2(_1742_),
    .B1(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__nand2_1 _3816_ (.A(\current_dst_addr[1][4] ),
    .B(_0385_),
    .Y(_1756_));
 sky130_fd_sc_hd__o22ai_1 _3817_ (.A1(net58),
    .A2(net1245),
    .B1(_1742_),
    .B2(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__a21oi_1 _3818_ (.A1(_1753_),
    .A2(_1755_),
    .B1(_1757_),
    .Y(_0066_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input167 (.A(channel_length[15]),
    .X(net167));
 sky130_fd_sc_hd__nand3_1 _3820_ (.A(\current_dst_addr[1][2] ),
    .B(\current_dst_addr[1][3] ),
    .C(\current_dst_addr[1][4] ),
    .Y(_1759_));
 sky130_fd_sc_hd__a21oi_1 _3821_ (.A1(_1738_),
    .A2(_1759_),
    .B1(_1740_),
    .Y(_1760_));
 sky130_fd_sc_hd__nor2_1 _3822_ (.A(_1742_),
    .B(_1759_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _3823_ (.A(\current_dst_addr[1][5] ),
    .B(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__o221a_2 _3824_ (.A1(net59),
    .A2(net1245),
    .B1(_1760_),
    .B2(\current_dst_addr[1][5] ),
    .C1(_1762_),
    .X(_0067_));
 sky130_fd_sc_hd__nand3_1 _3825_ (.A(\current_dst_addr[1][4] ),
    .B(_0385_),
    .C(\current_dst_addr[1][5] ),
    .Y(_1763_));
 sky130_fd_sc_hd__a21oi_1 _3826_ (.A1(_1738_),
    .A2(_1763_),
    .B1(_1740_),
    .Y(_1764_));
 sky130_fd_sc_hd__nor2_1 _3827_ (.A(_1742_),
    .B(_1756_),
    .Y(_1765_));
 sky130_fd_sc_hd__nand3_1 _3828_ (.A(\current_dst_addr[1][5] ),
    .B(\current_dst_addr[1][6] ),
    .C(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__o221a_2 _3829_ (.A1(net60),
    .A2(net1245),
    .B1(_1764_),
    .B2(\current_dst_addr[1][6] ),
    .C1(_1766_),
    .X(_0068_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input166 (.A(channel_length[14]),
    .X(net166));
 sky130_fd_sc_hd__a311oi_1 _3831_ (.A1(\current_dst_addr[1][5] ),
    .A2(\current_dst_addr[1][6] ),
    .A3(_1761_),
    .B1(net1247),
    .C1(\current_dst_addr[1][7] ),
    .Y(_1768_));
 sky130_fd_sc_hd__nand3_1 _3832_ (.A(\current_dst_addr[1][5] ),
    .B(\current_dst_addr[1][6] ),
    .C(\current_dst_addr[1][7] ),
    .Y(_1769_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input165 (.A(channel_length[13]),
    .X(net165));
 sky130_fd_sc_hd__o32ai_1 _3834_ (.A1(_1742_),
    .A2(_1759_),
    .A3(_1769_),
    .B1(net1245),
    .B2(net61),
    .Y(_1771_));
 sky130_fd_sc_hd__nor2_1 _3835_ (.A(_1768_),
    .B(_1771_),
    .Y(_0069_));
 sky130_fd_sc_hd__nor2_1 _3836_ (.A(_1756_),
    .B(_1769_),
    .Y(_1772_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input164 (.A(channel_length[12]),
    .X(net164));
 sky130_fd_sc_hd__nor2_1 _3838_ (.A(net63),
    .B(net1245),
    .Y(_1774_));
 sky130_fd_sc_hd__o21ai_0 _3839_ (.A1(_1756_),
    .A2(_1769_),
    .B1(_1738_),
    .Y(_1775_));
 sky130_fd_sc_hd__a21oi_1 _3840_ (.A1(_1754_),
    .A2(_1775_),
    .B1(\current_dst_addr[1][8] ),
    .Y(_1776_));
 sky130_fd_sc_hd__a311oi_1 _3841_ (.A1(\current_dst_addr[1][8] ),
    .A2(_1738_),
    .A3(_1772_),
    .B1(_1774_),
    .C1(_1776_),
    .Y(_0070_));
 sky130_fd_sc_hd__nor2_1 _3842_ (.A(_1759_),
    .B(_1769_),
    .Y(_1777_));
 sky130_fd_sc_hd__a21oi_1 _3843_ (.A1(\current_dst_addr[1][8] ),
    .A2(_1777_),
    .B1(_1742_),
    .Y(_1778_));
 sky130_fd_sc_hd__nor2_1 _3844_ (.A(_1740_),
    .B(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_1 _3845_ (.A(\current_dst_addr[1][8] ),
    .B(\current_dst_addr[1][9] ),
    .Y(_1780_));
 sky130_fd_sc_hd__nor3_1 _3846_ (.A(_1759_),
    .B(_1769_),
    .C(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _3847_ (.A(_1738_),
    .B(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__o221a_2 _3848_ (.A1(net64),
    .A2(net1245),
    .B1(_1779_),
    .B2(\current_dst_addr[1][9] ),
    .C1(_1782_),
    .X(_0071_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input163 (.A(channel_length[127]),
    .X(net163));
 sky130_fd_sc_hd__nand3_1 _3850_ (.A(\current_dst_addr[1][8] ),
    .B(\current_dst_addr[1][9] ),
    .C(_1772_),
    .Y(_1784_));
 sky130_fd_sc_hd__nor2_1 _3851_ (.A(_1742_),
    .B(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__a21oi_1 _3852_ (.A1(_1738_),
    .A2(_1784_),
    .B1(_1740_),
    .Y(_1786_));
 sky130_fd_sc_hd__nor2_1 _3853_ (.A(\current_dst_addr[1][10] ),
    .B(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input162 (.A(channel_length[126]),
    .X(net162));
 sky130_fd_sc_hd__nor2_1 _3855_ (.A(net65),
    .B(_1748_),
    .Y(_1789_));
 sky130_fd_sc_hd__a211oi_1 _3856_ (.A1(\current_dst_addr[1][10] ),
    .A2(_1785_),
    .B1(_1787_),
    .C1(_1789_),
    .Y(_0042_));
 sky130_fd_sc_hd__and2_1 _3857_ (.A(_1738_),
    .B(_1781_),
    .X(_1790_));
 sky130_fd_sc_hd__nor2_1 _3858_ (.A(net66),
    .B(_1748_),
    .Y(_1791_));
 sky130_fd_sc_hd__a211oi_1 _3859_ (.A1(\current_dst_addr[1][10] ),
    .A2(_1790_),
    .B1(net1246),
    .C1(\current_dst_addr[1][11] ),
    .Y(_1792_));
 sky130_fd_sc_hd__a311oi_1 _3860_ (.A1(\current_dst_addr[1][10] ),
    .A2(\current_dst_addr[1][11] ),
    .A3(_1790_),
    .B1(_1791_),
    .C1(_1792_),
    .Y(_0043_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input161 (.A(channel_length[125]),
    .X(net161));
 sky130_fd_sc_hd__nor2_1 _3862_ (.A(net67),
    .B(_1748_),
    .Y(_1794_));
 sky130_fd_sc_hd__a311oi_1 _3863_ (.A1(\current_dst_addr[1][10] ),
    .A2(\current_dst_addr[1][11] ),
    .A3(_1785_),
    .B1(net1246),
    .C1(\current_dst_addr[1][12] ),
    .Y(_1795_));
 sky130_fd_sc_hd__and4_1 _3864_ (.A(\current_dst_addr[1][10] ),
    .B(\current_dst_addr[1][11] ),
    .C(\current_dst_addr[1][12] ),
    .D(_1785_),
    .X(_1796_));
 sky130_fd_sc_hd__nor3_1 _3865_ (.A(_1794_),
    .B(_1795_),
    .C(_1796_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand4_1 _3866_ (.A(\current_dst_addr[1][10] ),
    .B(\current_dst_addr[1][11] ),
    .C(\current_dst_addr[1][12] ),
    .D(_1790_),
    .Y(_1797_));
 sky130_fd_sc_hd__nor2_1 _3867_ (.A(\current_dst_addr[1][13] ),
    .B(net1246),
    .Y(_1798_));
 sky130_fd_sc_hd__nand4_1 _3868_ (.A(\current_dst_addr[1][10] ),
    .B(\current_dst_addr[1][11] ),
    .C(\current_dst_addr[1][12] ),
    .D(\current_dst_addr[1][13] ),
    .Y(_1799_));
 sky130_fd_sc_hd__o22ai_1 _3869_ (.A1(net68),
    .A2(_1748_),
    .B1(_1782_),
    .B2(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__a21oi_1 _3870_ (.A1(_1797_),
    .A2(_1798_),
    .B1(_1800_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_1 _3871_ (.A(\current_dst_addr[1][14] ),
    .Y(_1801_));
 sky130_fd_sc_hd__nor2_1 _3872_ (.A(_1801_),
    .B(_1799_),
    .Y(_1802_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input160 (.A(channel_length[124]),
    .X(net160));
 sky130_fd_sc_hd__nor3_1 _3874_ (.A(_1742_),
    .B(_1784_),
    .C(_1799_),
    .Y(_1804_));
 sky130_fd_sc_hd__nor3_1 _3875_ (.A(\current_dst_addr[1][14] ),
    .B(net1246),
    .C(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__nor2_1 _3876_ (.A(net69),
    .B(_1748_),
    .Y(_1806_));
 sky130_fd_sc_hd__a211oi_1 _3877_ (.A1(_1785_),
    .A2(_1802_),
    .B1(_1805_),
    .C1(_1806_),
    .Y(_0046_));
 sky130_fd_sc_hd__a21oi_1 _3878_ (.A1(_1781_),
    .A2(_1802_),
    .B1(_1742_),
    .Y(_1807_));
 sky130_fd_sc_hd__nor2_1 _3879_ (.A(_1740_),
    .B(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__nor2_1 _3880_ (.A(\current_dst_addr[1][15] ),
    .B(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__nand2_1 _3881_ (.A(\current_dst_addr[1][15] ),
    .B(_1802_),
    .Y(_1810_));
 sky130_fd_sc_hd__o22ai_1 _3882_ (.A1(net70),
    .A2(_1748_),
    .B1(_1782_),
    .B2(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__nor2_1 _3883_ (.A(_1809_),
    .B(_1811_),
    .Y(_0047_));
 sky130_fd_sc_hd__and2_1 _3884_ (.A(\current_dst_addr[1][15] ),
    .B(_1802_),
    .X(_1812_));
 sky130_fd_sc_hd__o21ai_0 _3885_ (.A1(_1784_),
    .A2(_1810_),
    .B1(_1738_),
    .Y(_1813_));
 sky130_fd_sc_hd__a21oi_1 _3886_ (.A1(_1754_),
    .A2(_1813_),
    .B1(\current_dst_addr[1][16] ),
    .Y(_1814_));
 sky130_fd_sc_hd__nor2_1 _3887_ (.A(net71),
    .B(_1748_),
    .Y(_1815_));
 sky130_fd_sc_hd__a311oi_1 _3888_ (.A1(\current_dst_addr[1][16] ),
    .A2(_1785_),
    .A3(_1812_),
    .B1(_1814_),
    .C1(_1815_),
    .Y(_0048_));
 sky130_fd_sc_hd__a311oi_1 _3889_ (.A1(\current_dst_addr[1][16] ),
    .A2(_1790_),
    .A3(_1812_),
    .B1(\current_dst_addr[1][17] ),
    .C1(net1246),
    .Y(_1816_));
 sky130_fd_sc_hd__nand4_1 _3890_ (.A(\current_dst_addr[1][16] ),
    .B(\current_dst_addr[1][17] ),
    .C(_1790_),
    .D(_1812_),
    .Y(_1817_));
 sky130_fd_sc_hd__o21ai_0 _3891_ (.A1(net72),
    .A2(_1748_),
    .B1(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__nor2_1 _3892_ (.A(_1816_),
    .B(_1818_),
    .Y(_0049_));
 sky130_fd_sc_hd__nor3_1 _3893_ (.A(_1756_),
    .B(_1769_),
    .C(_1780_),
    .Y(_1819_));
 sky130_fd_sc_hd__nand4_1 _3894_ (.A(\current_dst_addr[1][14] ),
    .B(\current_dst_addr[1][15] ),
    .C(\current_dst_addr[1][16] ),
    .D(\current_dst_addr[1][17] ),
    .Y(_1820_));
 sky130_fd_sc_hd__nor2_1 _3895_ (.A(_1799_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__and3_1 _3896_ (.A(_1738_),
    .B(_1819_),
    .C(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__nor3_1 _3897_ (.A(\current_dst_addr[1][18] ),
    .B(net1246),
    .C(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__nor2_1 _3898_ (.A(net74),
    .B(net1245),
    .Y(_1824_));
 sky130_fd_sc_hd__a211oi_1 _3899_ (.A1(\current_dst_addr[1][18] ),
    .A2(_1822_),
    .B1(_1823_),
    .C1(_1824_),
    .Y(_0050_));
 sky130_fd_sc_hd__nor3_1 _3900_ (.A(_1782_),
    .B(_1799_),
    .C(_1820_),
    .Y(_1825_));
 sky130_fd_sc_hd__a211oi_1 _3901_ (.A1(\current_dst_addr[1][18] ),
    .A2(_1825_),
    .B1(net1246),
    .C1(\current_dst_addr[1][19] ),
    .Y(_1826_));
 sky130_fd_sc_hd__nor2_1 _3902_ (.A(net75),
    .B(net1245),
    .Y(_1827_));
 sky130_fd_sc_hd__a311oi_1 _3903_ (.A1(\current_dst_addr[1][18] ),
    .A2(\current_dst_addr[1][19] ),
    .A3(_1825_),
    .B1(_1826_),
    .C1(_1827_),
    .Y(_0051_));
 sky130_fd_sc_hd__and3_1 _3904_ (.A(\current_dst_addr[1][18] ),
    .B(\current_dst_addr[1][19] ),
    .C(\current_dst_addr[1][20] ),
    .X(_1828_));
 sky130_fd_sc_hd__a311oi_1 _3905_ (.A1(\current_dst_addr[1][18] ),
    .A2(\current_dst_addr[1][19] ),
    .A3(_1822_),
    .B1(net1246),
    .C1(\current_dst_addr[1][20] ),
    .Y(_1829_));
 sky130_fd_sc_hd__nor2_1 _3906_ (.A(net76),
    .B(net1245),
    .Y(_1830_));
 sky130_fd_sc_hd__a211oi_1 _3907_ (.A1(_1822_),
    .A2(_1828_),
    .B1(_1829_),
    .C1(_1830_),
    .Y(_0052_));
 sky130_fd_sc_hd__nor2_1 _3908_ (.A(net77),
    .B(net1245),
    .Y(_1831_));
 sky130_fd_sc_hd__a211oi_1 _3909_ (.A1(_1825_),
    .A2(_1828_),
    .B1(\current_dst_addr[1][21] ),
    .C1(net1246),
    .Y(_1832_));
 sky130_fd_sc_hd__a311oi_1 _3910_ (.A1(\current_dst_addr[1][21] ),
    .A2(_1825_),
    .A3(_1828_),
    .B1(_1831_),
    .C1(_1832_),
    .Y(_0053_));
 sky130_fd_sc_hd__nor2_1 _3911_ (.A(net78),
    .B(net1245),
    .Y(_1833_));
 sky130_fd_sc_hd__a311oi_1 _3912_ (.A1(\current_dst_addr[1][21] ),
    .A2(_1822_),
    .A3(_1828_),
    .B1(\current_dst_addr[1][22] ),
    .C1(net1246),
    .Y(_1834_));
 sky130_fd_sc_hd__and3_1 _3913_ (.A(\current_dst_addr[1][21] ),
    .B(\current_dst_addr[1][22] ),
    .C(_1828_),
    .X(_1835_));
 sky130_fd_sc_hd__and4_1 _3914_ (.A(_1738_),
    .B(_1819_),
    .C(_1821_),
    .D(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input159 (.A(channel_length[123]),
    .X(net159));
 sky130_fd_sc_hd__nor3_1 _3916_ (.A(_1833_),
    .B(_1834_),
    .C(_1836_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand3_1 _3917_ (.A(_1781_),
    .B(_1821_),
    .C(_1835_),
    .Y(_1838_));
 sky130_fd_sc_hd__a21oi_1 _3918_ (.A1(_1738_),
    .A2(_1838_),
    .B1(_1740_),
    .Y(_1839_));
 sky130_fd_sc_hd__and4_1 _3919_ (.A(_1738_),
    .B(_1781_),
    .C(_1821_),
    .D(_1835_),
    .X(_1840_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input158 (.A(channel_length[122]),
    .X(net158));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(\current_dst_addr[1][23] ),
    .B(_1840_),
    .Y(_1842_));
 sky130_fd_sc_hd__o221a_2 _3922_ (.A1(net79),
    .A2(_1748_),
    .B1(_1839_),
    .B2(\current_dst_addr[1][23] ),
    .C1(_1842_),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_1 _3923_ (.A(net80),
    .B(_1748_),
    .Y(_1843_));
 sky130_fd_sc_hd__a211oi_1 _3924_ (.A1(\current_dst_addr[1][23] ),
    .A2(_1836_),
    .B1(net1246),
    .C1(\current_dst_addr[1][24] ),
    .Y(_1844_));
 sky130_fd_sc_hd__a311oi_1 _3925_ (.A1(\current_dst_addr[1][23] ),
    .A2(\current_dst_addr[1][24] ),
    .A3(_1836_),
    .B1(_1843_),
    .C1(_1844_),
    .Y(_0056_));
 sky130_fd_sc_hd__and3_1 _3926_ (.A(\current_dst_addr[1][23] ),
    .B(\current_dst_addr[1][24] ),
    .C(\current_dst_addr[1][25] ),
    .X(_1845_));
 sky130_fd_sc_hd__nor2_1 _3927_ (.A(net81),
    .B(_1748_),
    .Y(_1846_));
 sky130_fd_sc_hd__a311oi_1 _3928_ (.A1(\current_dst_addr[1][23] ),
    .A2(\current_dst_addr[1][24] ),
    .A3(_1840_),
    .B1(net1246),
    .C1(\current_dst_addr[1][25] ),
    .Y(_1847_));
 sky130_fd_sc_hd__a211oi_1 _3929_ (.A1(_1840_),
    .A2(_1845_),
    .B1(_1846_),
    .C1(_1847_),
    .Y(_0057_));
 sky130_fd_sc_hd__nor2_1 _3930_ (.A(net82),
    .B(_1748_),
    .Y(_1848_));
 sky130_fd_sc_hd__a211oi_1 _3931_ (.A1(_1836_),
    .A2(_1845_),
    .B1(\current_dst_addr[1][26] ),
    .C1(net1246),
    .Y(_1849_));
 sky130_fd_sc_hd__a311oi_1 _3932_ (.A1(\current_dst_addr[1][26] ),
    .A2(_1836_),
    .A3(_1845_),
    .B1(_1848_),
    .C1(_1849_),
    .Y(_0058_));
 sky130_fd_sc_hd__and3_1 _3933_ (.A(\current_dst_addr[1][26] ),
    .B(\current_dst_addr[1][27] ),
    .C(_1845_),
    .X(_1850_));
 sky130_fd_sc_hd__a311oi_1 _3934_ (.A1(\current_dst_addr[1][26] ),
    .A2(_1840_),
    .A3(_1845_),
    .B1(\current_dst_addr[1][27] ),
    .C1(net1246),
    .Y(_1851_));
 sky130_fd_sc_hd__nor2_1 _3935_ (.A(net83),
    .B(_1748_),
    .Y(_1852_));
 sky130_fd_sc_hd__a211oi_1 _3936_ (.A1(_1840_),
    .A2(_1850_),
    .B1(_1851_),
    .C1(_1852_),
    .Y(_0059_));
 sky130_fd_sc_hd__and2_0 _3937_ (.A(\current_dst_addr[1][28] ),
    .B(_1850_),
    .X(_1853_));
 sky130_fd_sc_hd__a211oi_1 _3938_ (.A1(_1836_),
    .A2(_1850_),
    .B1(\current_dst_addr[1][28] ),
    .C1(net1246),
    .Y(_1854_));
 sky130_fd_sc_hd__nor2_1 _3939_ (.A(net85),
    .B(_1748_),
    .Y(_1855_));
 sky130_fd_sc_hd__a211oi_1 _3940_ (.A1(_1836_),
    .A2(_1853_),
    .B1(_1854_),
    .C1(_1855_),
    .Y(_0060_));
 sky130_fd_sc_hd__nor2_1 _3941_ (.A(net86),
    .B(net1245),
    .Y(_1856_));
 sky130_fd_sc_hd__a211oi_1 _3942_ (.A1(_1840_),
    .A2(_1853_),
    .B1(\current_dst_addr[1][29] ),
    .C1(net1246),
    .Y(_1857_));
 sky130_fd_sc_hd__a311oi_1 _3943_ (.A1(\current_dst_addr[1][29] ),
    .A2(_1840_),
    .A3(_1853_),
    .B1(_1856_),
    .C1(_1857_),
    .Y(_0061_));
 sky130_fd_sc_hd__a311oi_1 _3944_ (.A1(\current_dst_addr[1][29] ),
    .A2(_1836_),
    .A3(_1853_),
    .B1(\current_dst_addr[1][30] ),
    .C1(net1246),
    .Y(_1858_));
 sky130_fd_sc_hd__nand4_1 _3945_ (.A(\current_dst_addr[1][29] ),
    .B(\current_dst_addr[1][30] ),
    .C(_1836_),
    .D(_1853_),
    .Y(_1859_));
 sky130_fd_sc_hd__o21ai_0 _3946_ (.A1(net87),
    .A2(net1245),
    .B1(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nor2_1 _3947_ (.A(_1858_),
    .B(_1860_),
    .Y(_0063_));
 sky130_fd_sc_hd__and4_1 _3948_ (.A(\current_dst_addr[1][29] ),
    .B(\current_dst_addr[1][30] ),
    .C(_1840_),
    .D(_1853_),
    .X(_1861_));
 sky130_fd_sc_hd__nor3_1 _3949_ (.A(\current_dst_addr[1][31] ),
    .B(net1246),
    .C(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__nor2_1 _3950_ (.A(net88),
    .B(_1748_),
    .Y(_1863_));
 sky130_fd_sc_hd__a211oi_1 _3951_ (.A1(\current_dst_addr[1][31] ),
    .A2(_1861_),
    .B1(_1862_),
    .C1(_1863_),
    .Y(_0064_));
 sky130_fd_sc_hd__nor2b_1 _3952_ (.A(net557),
    .B_N(net397),
    .Y(_1864_));
 sky130_fd_sc_hd__nor2_1 _3953_ (.A(net558),
    .B(net554),
    .Y(_1865_));
 sky130_fd_sc_hd__and3_2 _3954_ (.A(net129),
    .B(_1864_),
    .C(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input157 (.A(channel_length[121]),
    .X(net157));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input156 (.A(channel_length[120]),
    .X(net156));
 sky130_fd_sc_hd__nand4bb_4 _3957_ (.A_N(net554),
    .B_N(net557),
    .C(net401),
    .D(net558),
    .Y(_1869_));
 sky130_fd_sc_hd__nor2_1 _3958_ (.A(net261),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__nor2_1 _3959_ (.A(_1866_),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__nor4bb_4 _3960_ (.A(net554),
    .B(net557),
    .C_N(net401),
    .D_N(net558),
    .Y(_1872_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input155 (.A(channel_length[11]),
    .X(net155));
 sky130_fd_sc_hd__nand2b_1 _3962_ (.A_N(net261),
    .B(_1872_),
    .Y(_1874_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input154 (.A(channel_length[119]),
    .X(net154));
 sky130_fd_sc_hd__nor2_1 _3964_ (.A(\current_dst_addr[0][2] ),
    .B(_1874_),
    .Y(_1876_));
 sky130_fd_sc_hd__a221o_1 _3965_ (.A1(net51),
    .A2(_1866_),
    .B1(_1871_),
    .B2(\current_dst_addr[0][2] ),
    .C1(_1876_),
    .X(_0032_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input153 (.A(channel_length[118]),
    .X(net153));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input152 (.A(channel_length[117]),
    .X(net152));
 sky130_fd_sc_hd__nand2_1 _3968_ (.A(net62),
    .B(_1866_),
    .Y(_1879_));
 sky130_fd_sc_hd__nand3_4 _3969_ (.A(net129),
    .B(_1864_),
    .C(_1865_),
    .Y(_1880_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input151 (.A(channel_length[116]),
    .X(net151));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input150 (.A(channel_length[115]),
    .X(net150));
 sky130_fd_sc_hd__nand2_1 _3972_ (.A(\current_dst_addr[0][3] ),
    .B(_1880_),
    .Y(_1883_));
 sky130_fd_sc_hd__nor2_1 _3973_ (.A(_0388_),
    .B(_1874_),
    .Y(_1884_));
 sky130_fd_sc_hd__a31oi_1 _3974_ (.A1(_1874_),
    .A2(_1879_),
    .A3(_1883_),
    .B1(_1884_),
    .Y(_0035_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_0387_),
    .B(_1874_),
    .Y(_1885_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_1871_),
    .B(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__nor2_1 _3977_ (.A(\current_dst_addr[0][4] ),
    .B(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input149 (.A(channel_length[114]),
    .X(net149));
 sky130_fd_sc_hd__nand2_1 _3979_ (.A(\current_dst_addr[0][4] ),
    .B(_0387_),
    .Y(_1889_));
 sky130_fd_sc_hd__o22ai_1 _3980_ (.A1(net73),
    .A2(_1880_),
    .B1(_1874_),
    .B2(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__nor2_1 _3981_ (.A(_1887_),
    .B(_1890_),
    .Y(_0036_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input148 (.A(channel_length[113]),
    .X(net148));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input147 (.A(channel_length[112]),
    .X(net147));
 sky130_fd_sc_hd__nand3_1 _3984_ (.A(\current_dst_addr[0][2] ),
    .B(\current_dst_addr[0][3] ),
    .C(\current_dst_addr[0][4] ),
    .Y(_1893_));
 sky130_fd_sc_hd__a21oi_1 _3985_ (.A1(_1870_),
    .A2(_1893_),
    .B1(_1871_),
    .Y(_1894_));
 sky130_fd_sc_hd__nor2_1 _3986_ (.A(_1874_),
    .B(_1893_),
    .Y(_1895_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(\current_dst_addr[0][5] ),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__o221a_2 _3988_ (.A1(net84),
    .A2(_1880_),
    .B1(_1894_),
    .B2(\current_dst_addr[0][5] ),
    .C1(_1896_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _3989_ (.A(_1880_),
    .B(_1874_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand3_1 _3990_ (.A(\current_dst_addr[0][4] ),
    .B(_0387_),
    .C(\current_dst_addr[0][5] ),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(_1870_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__a21oi_1 _3992_ (.A1(_1897_),
    .A2(_1899_),
    .B1(\current_dst_addr[0][6] ),
    .Y(_1900_));
 sky130_fd_sc_hd__nand2_1 _3993_ (.A(\current_dst_addr[0][5] ),
    .B(\current_dst_addr[0][6] ),
    .Y(_1901_));
 sky130_fd_sc_hd__o32ai_1 _3994_ (.A1(_1874_),
    .A2(_1889_),
    .A3(_1901_),
    .B1(_1880_),
    .B2(net95),
    .Y(_1902_));
 sky130_fd_sc_hd__nor2_1 _3995_ (.A(_1900_),
    .B(_1902_),
    .Y(_0038_));
 sky130_fd_sc_hd__and3_1 _3996_ (.A(\current_dst_addr[0][5] ),
    .B(\current_dst_addr[0][6] ),
    .C(\current_dst_addr[0][7] ),
    .X(_1903_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input146 (.A(channel_length[111]),
    .X(net146));
 sky130_fd_sc_hd__nor2_1 _3998_ (.A(net106),
    .B(_1880_),
    .Y(_1905_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input145 (.A(channel_length[110]),
    .X(net145));
 sky130_fd_sc_hd__a311oi_1 _4000_ (.A1(\current_dst_addr[0][5] ),
    .A2(\current_dst_addr[0][6] ),
    .A3(_1895_),
    .B1(_1866_),
    .C1(\current_dst_addr[0][7] ),
    .Y(_1907_));
 sky130_fd_sc_hd__a211oi_1 _4001_ (.A1(_1895_),
    .A2(_1903_),
    .B1(_1905_),
    .C1(_1907_),
    .Y(_0039_));
 sky130_fd_sc_hd__nand3_1 _4002_ (.A(\current_dst_addr[0][4] ),
    .B(_0387_),
    .C(_1903_),
    .Y(_1908_));
 sky130_fd_sc_hd__a21oi_1 _4003_ (.A1(_1870_),
    .A2(_1908_),
    .B1(_1871_),
    .Y(_1909_));
 sky130_fd_sc_hd__nand3_1 _4004_ (.A(\current_dst_addr[0][5] ),
    .B(\current_dst_addr[0][6] ),
    .C(\current_dst_addr[0][7] ),
    .Y(_1910_));
 sky130_fd_sc_hd__nor2_1 _4005_ (.A(_1889_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nand3_1 _4006_ (.A(\current_dst_addr[0][8] ),
    .B(_1870_),
    .C(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__o221a_2 _4007_ (.A1(net117),
    .A2(_1880_),
    .B1(_1909_),
    .B2(\current_dst_addr[0][8] ),
    .C1(_1912_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_1 _4008_ (.A(net128),
    .B(_1880_),
    .Y(_1913_));
 sky130_fd_sc_hd__nor2_1 _4009_ (.A(_1893_),
    .B(_1910_),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(\current_dst_addr[0][8] ),
    .B(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__a21oi_1 _4011_ (.A1(_1870_),
    .A2(_1915_),
    .B1(_1871_),
    .Y(_1916_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(\current_dst_addr[0][9] ),
    .B(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__nand2b_1 _4013_ (.A_N(_1893_),
    .B(_1903_),
    .Y(_1918_));
 sky130_fd_sc_hd__nand2_1 _4014_ (.A(\current_dst_addr[0][8] ),
    .B(\current_dst_addr[0][9] ),
    .Y(_1919_));
 sky130_fd_sc_hd__nor3_1 _4015_ (.A(_1874_),
    .B(_1918_),
    .C(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__nor3_1 _4016_ (.A(_1913_),
    .B(_1917_),
    .C(_1920_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand3_1 _4017_ (.A(\current_dst_addr[0][8] ),
    .B(\current_dst_addr[0][9] ),
    .C(_1911_),
    .Y(_1921_));
 sky130_fd_sc_hd__nor2_1 _4018_ (.A(_1874_),
    .B(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__a21oi_1 _4019_ (.A1(_1870_),
    .A2(_1921_),
    .B1(_1871_),
    .Y(_1923_));
 sky130_fd_sc_hd__nor2_1 _4020_ (.A(\current_dst_addr[0][10] ),
    .B(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__nor2_1 _4021_ (.A(net12),
    .B(_1880_),
    .Y(_1925_));
 sky130_fd_sc_hd__a211oi_1 _4022_ (.A1(\current_dst_addr[0][10] ),
    .A2(_1922_),
    .B1(_1924_),
    .C1(_1925_),
    .Y(_0012_));
 sky130_fd_sc_hd__nor2_1 _4023_ (.A(net23),
    .B(_1880_),
    .Y(_1926_));
 sky130_fd_sc_hd__a211oi_1 _4024_ (.A1(\current_dst_addr[0][10] ),
    .A2(_1920_),
    .B1(_1866_),
    .C1(\current_dst_addr[0][11] ),
    .Y(_1927_));
 sky130_fd_sc_hd__a311oi_1 _4025_ (.A1(\current_dst_addr[0][10] ),
    .A2(\current_dst_addr[0][11] ),
    .A3(_1920_),
    .B1(_1926_),
    .C1(_1927_),
    .Y(_0013_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input144 (.A(channel_length[10]),
    .X(net144));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(\current_dst_addr[0][10] ),
    .B(\current_dst_addr[0][11] ),
    .Y(_1929_));
 sky130_fd_sc_hd__nor3_1 _4028_ (.A(_1874_),
    .B(_1921_),
    .C(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__nor2_1 _4029_ (.A(net32),
    .B(_1880_),
    .Y(_1931_));
 sky130_fd_sc_hd__a21oi_1 _4030_ (.A1(\current_dst_addr[0][12] ),
    .A2(_1930_),
    .B1(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__o31a_1 _4031_ (.A1(\current_dst_addr[0][12] ),
    .A2(_1866_),
    .A3(_1930_),
    .B1(_1932_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_1 _4032_ (.A(\current_dst_addr[0][10] ),
    .B(\current_dst_addr[0][11] ),
    .C(\current_dst_addr[0][12] ),
    .X(_1933_));
 sky130_fd_sc_hd__a211oi_1 _4033_ (.A1(_1920_),
    .A2(_1933_),
    .B1(\current_dst_addr[0][13] ),
    .C1(_1866_),
    .Y(_1934_));
 sky130_fd_sc_hd__nor2_1 _4034_ (.A(net33),
    .B(net1243),
    .Y(_1935_));
 sky130_fd_sc_hd__a311oi_1 _4035_ (.A1(\current_dst_addr[0][13] ),
    .A2(_1920_),
    .A3(_1933_),
    .B1(_1934_),
    .C1(_1935_),
    .Y(_0015_));
 sky130_fd_sc_hd__and4_1 _4036_ (.A(\current_dst_addr[0][10] ),
    .B(\current_dst_addr[0][11] ),
    .C(\current_dst_addr[0][12] ),
    .D(\current_dst_addr[0][13] ),
    .X(_1936_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input143 (.A(channel_length[109]),
    .X(net143));
 sky130_fd_sc_hd__a211oi_1 _4038_ (.A1(_1922_),
    .A2(_1936_),
    .B1(\current_dst_addr[0][14] ),
    .C1(_1866_),
    .Y(_1938_));
 sky130_fd_sc_hd__nor2_1 _4039_ (.A(net34),
    .B(_1880_),
    .Y(_1939_));
 sky130_fd_sc_hd__a311oi_1 _4040_ (.A1(\current_dst_addr[0][14] ),
    .A2(_1922_),
    .A3(_1936_),
    .B1(_1938_),
    .C1(_1939_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_1 _4041_ (.A(\current_dst_addr[0][15] ),
    .Y(_1940_));
 sky130_fd_sc_hd__nand2_1 _4042_ (.A(\current_dst_addr[0][14] ),
    .B(_1936_),
    .Y(_1941_));
 sky130_fd_sc_hd__nor3_1 _4043_ (.A(_1918_),
    .B(_1919_),
    .C(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__o21ai_0 _4044_ (.A1(_1874_),
    .A2(_1942_),
    .B1(_1897_),
    .Y(_1943_));
 sky130_fd_sc_hd__nand3_1 _4045_ (.A(\current_dst_addr[0][15] ),
    .B(_1870_),
    .C(_1942_),
    .Y(_1944_));
 sky130_fd_sc_hd__o21ai_0 _4046_ (.A1(net35),
    .A2(_1880_),
    .B1(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__a21oi_1 _4047_ (.A1(_1940_),
    .A2(_1943_),
    .B1(_1945_),
    .Y(_0017_));
 sky130_fd_sc_hd__and3_1 _4048_ (.A(\current_dst_addr[0][14] ),
    .B(\current_dst_addr[0][15] ),
    .C(_1936_),
    .X(_1946_));
 sky130_fd_sc_hd__nand3_1 _4049_ (.A(\current_dst_addr[0][14] ),
    .B(\current_dst_addr[0][15] ),
    .C(_1936_),
    .Y(_1947_));
 sky130_fd_sc_hd__o21ai_0 _4050_ (.A1(_1921_),
    .A2(_1947_),
    .B1(_1870_),
    .Y(_1948_));
 sky130_fd_sc_hd__a21oi_1 _4051_ (.A1(_1897_),
    .A2(_1948_),
    .B1(\current_dst_addr[0][16] ),
    .Y(_1949_));
 sky130_fd_sc_hd__nor2_1 _4052_ (.A(net36),
    .B(_1880_),
    .Y(_1950_));
 sky130_fd_sc_hd__a311oi_1 _4053_ (.A1(\current_dst_addr[0][16] ),
    .A2(_1922_),
    .A3(_1946_),
    .B1(_1949_),
    .C1(_1950_),
    .Y(_0018_));
 sky130_fd_sc_hd__a311oi_1 _4054_ (.A1(\current_dst_addr[0][16] ),
    .A2(_1920_),
    .A3(_1946_),
    .B1(\current_dst_addr[0][17] ),
    .C1(_1866_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand4_1 _4055_ (.A(\current_dst_addr[0][16] ),
    .B(\current_dst_addr[0][17] ),
    .C(_1920_),
    .D(_1946_),
    .Y(_1952_));
 sky130_fd_sc_hd__o21ai_0 _4056_ (.A1(net37),
    .A2(_1880_),
    .B1(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__nor2_1 _4057_ (.A(_1951_),
    .B(_1953_),
    .Y(_0019_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input142 (.A(channel_length[108]),
    .X(net142));
 sky130_fd_sc_hd__and4_1 _4059_ (.A(\current_dst_addr[0][8] ),
    .B(\current_dst_addr[0][9] ),
    .C(\current_dst_addr[0][16] ),
    .D(\current_dst_addr[0][17] ),
    .X(_1955_));
 sky130_fd_sc_hd__nand4_1 _4060_ (.A(\current_dst_addr[0][14] ),
    .B(\current_dst_addr[0][15] ),
    .C(_1936_),
    .D(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__nor2_1 _4061_ (.A(_1908_),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__o21ai_0 _4062_ (.A1(_1908_),
    .A2(_1956_),
    .B1(_1870_),
    .Y(_1958_));
 sky130_fd_sc_hd__a21oi_1 _4063_ (.A1(_1897_),
    .A2(_1958_),
    .B1(\current_dst_addr[0][18] ),
    .Y(_1959_));
 sky130_fd_sc_hd__nor2_1 _4064_ (.A(net38),
    .B(_1880_),
    .Y(_1960_));
 sky130_fd_sc_hd__a311oi_1 _4065_ (.A1(\current_dst_addr[0][18] ),
    .A2(_1870_),
    .A3(_1957_),
    .B1(_1959_),
    .C1(_1960_),
    .Y(_0020_));
 sky130_fd_sc_hd__nor2_1 _4066_ (.A(_1918_),
    .B(_1956_),
    .Y(_1961_));
 sky130_fd_sc_hd__a311oi_1 _4067_ (.A1(\current_dst_addr[0][18] ),
    .A2(_1870_),
    .A3(_1961_),
    .B1(\current_dst_addr[0][19] ),
    .C1(_1866_),
    .Y(_1962_));
 sky130_fd_sc_hd__nand4_1 _4068_ (.A(\current_dst_addr[0][18] ),
    .B(\current_dst_addr[0][19] ),
    .C(_1870_),
    .D(_1961_),
    .Y(_1963_));
 sky130_fd_sc_hd__o21ai_0 _4069_ (.A1(net39),
    .A2(_1880_),
    .B1(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__nor2_1 _4070_ (.A(_1962_),
    .B(_1964_),
    .Y(_0021_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input141 (.A(channel_length[107]),
    .X(net141));
 sky130_fd_sc_hd__nor2_1 _4072_ (.A(\current_dst_addr[0][20] ),
    .B(_1866_),
    .Y(_1966_));
 sky130_fd_sc_hd__nand4_1 _4073_ (.A(\current_dst_addr[0][18] ),
    .B(\current_dst_addr[0][19] ),
    .C(_1870_),
    .D(_1957_),
    .Y(_1967_));
 sky130_fd_sc_hd__mux2i_1 _4074_ (.A0(\current_dst_addr[0][20] ),
    .A1(_1966_),
    .S(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__o21a_1 _4075_ (.A1(net41),
    .A2(_1880_),
    .B1(_1968_),
    .X(_0022_));
 sky130_fd_sc_hd__nand3_1 _4076_ (.A(\current_dst_addr[0][18] ),
    .B(\current_dst_addr[0][19] ),
    .C(\current_dst_addr[0][20] ),
    .Y(_1969_));
 sky130_fd_sc_hd__nor2_1 _4077_ (.A(_1874_),
    .B(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__a211oi_1 _4078_ (.A1(_1961_),
    .A2(_1970_),
    .B1(\current_dst_addr[0][21] ),
    .C1(_1866_),
    .Y(_1971_));
 sky130_fd_sc_hd__nor2_1 _4079_ (.A(net42),
    .B(_1880_),
    .Y(_1972_));
 sky130_fd_sc_hd__a311oi_1 _4080_ (.A1(\current_dst_addr[0][21] ),
    .A2(_1961_),
    .A3(_1970_),
    .B1(_1971_),
    .C1(_1972_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_1 _4081_ (.A(\current_dst_addr[0][22] ),
    .Y(_1973_));
 sky130_fd_sc_hd__nand3_1 _4082_ (.A(\current_dst_addr[0][21] ),
    .B(_1957_),
    .C(_1970_),
    .Y(_1974_));
 sky130_fd_sc_hd__o22ai_1 _4083_ (.A1(net43),
    .A2(_1880_),
    .B1(_1974_),
    .B2(_1973_),
    .Y(_1975_));
 sky130_fd_sc_hd__a31oi_1 _4084_ (.A1(_1973_),
    .A2(_1880_),
    .A3(_1974_),
    .B1(_1975_),
    .Y(_0024_));
 sky130_fd_sc_hd__nand4_1 _4085_ (.A(\current_dst_addr[0][18] ),
    .B(\current_dst_addr[0][19] ),
    .C(\current_dst_addr[0][20] ),
    .D(\current_dst_addr[0][21] ),
    .Y(_1976_));
 sky130_fd_sc_hd__nor3_1 _4086_ (.A(_1973_),
    .B(_1874_),
    .C(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__and2_0 _4087_ (.A(_1961_),
    .B(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input140 (.A(channel_length[106]),
    .X(net140));
 sky130_fd_sc_hd__nor3_1 _4089_ (.A(\current_dst_addr[0][23] ),
    .B(_1866_),
    .C(_1978_),
    .Y(_1980_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input139 (.A(channel_length[105]),
    .X(net139));
 sky130_fd_sc_hd__nor2_1 _4091_ (.A(net44),
    .B(_1880_),
    .Y(_1982_));
 sky130_fd_sc_hd__a211oi_1 _4092_ (.A1(\current_dst_addr[0][23] ),
    .A2(_1978_),
    .B1(_1980_),
    .C1(_1982_),
    .Y(_0025_));
 sky130_fd_sc_hd__and2_1 _4093_ (.A(_1957_),
    .B(_1977_),
    .X(_1983_));
 sky130_fd_sc_hd__a211oi_1 _4094_ (.A1(\current_dst_addr[0][23] ),
    .A2(_1983_),
    .B1(_1866_),
    .C1(\current_dst_addr[0][24] ),
    .Y(_1984_));
 sky130_fd_sc_hd__nor2_1 _4095_ (.A(net45),
    .B(_1880_),
    .Y(_1985_));
 sky130_fd_sc_hd__a311oi_1 _4096_ (.A1(\current_dst_addr[0][23] ),
    .A2(\current_dst_addr[0][24] ),
    .A3(_1983_),
    .B1(_1984_),
    .C1(_1985_),
    .Y(_0026_));
 sky130_fd_sc_hd__and3_1 _4097_ (.A(\current_dst_addr[0][23] ),
    .B(\current_dst_addr[0][24] ),
    .C(\current_dst_addr[0][25] ),
    .X(_1986_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input138 (.A(channel_length[104]),
    .X(net138));
 sky130_fd_sc_hd__a311oi_1 _4099_ (.A1(\current_dst_addr[0][23] ),
    .A2(\current_dst_addr[0][24] ),
    .A3(_1978_),
    .B1(_1866_),
    .C1(\current_dst_addr[0][25] ),
    .Y(_1988_));
 sky130_fd_sc_hd__nor2_1 _4100_ (.A(net46),
    .B(_1880_),
    .Y(_1989_));
 sky130_fd_sc_hd__a211oi_1 _4101_ (.A1(_1978_),
    .A2(_1986_),
    .B1(_1988_),
    .C1(_1989_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_1 _4102_ (.A(net47),
    .B(_1880_),
    .Y(_1990_));
 sky130_fd_sc_hd__a211oi_1 _4103_ (.A1(_1983_),
    .A2(_1986_),
    .B1(\current_dst_addr[0][26] ),
    .C1(_1866_),
    .Y(_1991_));
 sky130_fd_sc_hd__a311oi_1 _4104_ (.A1(\current_dst_addr[0][26] ),
    .A2(_1983_),
    .A3(_1986_),
    .B1(_1990_),
    .C1(_1991_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand3_1 _4105_ (.A(\current_dst_addr[0][26] ),
    .B(\current_dst_addr[0][27] ),
    .C(_1986_),
    .Y(_1992_));
 sky130_fd_sc_hd__inv_1 _4106_ (.A(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__a311oi_1 _4107_ (.A1(\current_dst_addr[0][26] ),
    .A2(_1978_),
    .A3(_1986_),
    .B1(\current_dst_addr[0][27] ),
    .C1(_1866_),
    .Y(_1994_));
 sky130_fd_sc_hd__nor2_1 _4108_ (.A(net48),
    .B(_1880_),
    .Y(_1995_));
 sky130_fd_sc_hd__a211oi_1 _4109_ (.A1(_1978_),
    .A2(_1993_),
    .B1(_1994_),
    .C1(_1995_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand4_1 _4110_ (.A(\current_dst_addr[0][26] ),
    .B(\current_dst_addr[0][27] ),
    .C(\current_dst_addr[0][28] ),
    .D(_1986_),
    .Y(_1996_));
 sky130_fd_sc_hd__nor4_2 _4111_ (.A(_1973_),
    .B(_1874_),
    .C(_1976_),
    .D(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__a211oi_1 _4112_ (.A1(_1983_),
    .A2(_1993_),
    .B1(\current_dst_addr[0][28] ),
    .C1(_1866_),
    .Y(_1998_));
 sky130_fd_sc_hd__nor2_1 _4113_ (.A(net49),
    .B(_1880_),
    .Y(_1999_));
 sky130_fd_sc_hd__a211oi_1 _4114_ (.A1(_1957_),
    .A2(_1997_),
    .B1(_1998_),
    .C1(_1999_),
    .Y(_0030_));
 sky130_fd_sc_hd__nor2_1 _4115_ (.A(net50),
    .B(_1880_),
    .Y(_2000_));
 sky130_fd_sc_hd__a211oi_1 _4116_ (.A1(_1961_),
    .A2(_1997_),
    .B1(\current_dst_addr[0][29] ),
    .C1(_1866_),
    .Y(_2001_));
 sky130_fd_sc_hd__a311oi_1 _4117_ (.A1(\current_dst_addr[0][29] ),
    .A2(_1961_),
    .A3(_1997_),
    .B1(_2000_),
    .C1(_2001_),
    .Y(_0031_));
 sky130_fd_sc_hd__a311oi_1 _4118_ (.A1(\current_dst_addr[0][29] ),
    .A2(_1957_),
    .A3(_1997_),
    .B1(\current_dst_addr[0][30] ),
    .C1(_1866_),
    .Y(_2002_));
 sky130_fd_sc_hd__nand4_1 _4119_ (.A(\current_dst_addr[0][29] ),
    .B(\current_dst_addr[0][30] ),
    .C(_1957_),
    .D(_1997_),
    .Y(_2003_));
 sky130_fd_sc_hd__o21ai_0 _4120_ (.A1(net52),
    .A2(_1880_),
    .B1(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__nor2_1 _4121_ (.A(_2002_),
    .B(_2004_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_1 _4122_ (.A(\current_dst_addr[0][31] ),
    .Y(_2005_));
 sky130_fd_sc_hd__nand4_1 _4123_ (.A(\current_dst_addr[0][29] ),
    .B(\current_dst_addr[0][30] ),
    .C(_1961_),
    .D(_1997_),
    .Y(_2006_));
 sky130_fd_sc_hd__o22ai_1 _4124_ (.A1(net53),
    .A2(_1880_),
    .B1(_2006_),
    .B2(_2005_),
    .Y(_2007_));
 sky130_fd_sc_hd__a31oi_1 _4125_ (.A1(_2005_),
    .A2(_1880_),
    .A3(_2006_),
    .B1(_2007_),
    .Y(_0034_));
 sky130_fd_sc_hd__nor2_1 _4126_ (.A(net268),
    .B(_1470_),
    .Y(_2008_));
 sky130_fd_sc_hd__nor2_1 _4127_ (.A(net1251),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__nand2b_1 _4128_ (.A_N(net268),
    .B(_1474_),
    .Y(_2010_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input137 (.A(channel_length[103]),
    .X(net137));
 sky130_fd_sc_hd__nor2_1 _4130_ (.A(\current_src_addr[3][2] ),
    .B(_2010_),
    .Y(_2012_));
 sky130_fd_sc_hd__a221o_1 _4131_ (.A1(net394),
    .A2(net1251),
    .B1(_2009_),
    .B2(\current_src_addr[3][2] ),
    .C1(_2012_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _4132_ (.A(net395),
    .B(net1251),
    .Y(_2013_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(\current_src_addr[3][3] ),
    .B(net1250),
    .Y(_2014_));
 sky130_fd_sc_hd__nor2_1 _4134_ (.A(_0390_),
    .B(_2010_),
    .Y(_2015_));
 sky130_fd_sc_hd__a31oi_1 _4135_ (.A1(_2010_),
    .A2(_2013_),
    .A3(_2014_),
    .B1(_2015_),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_1 _4136_ (.A(\current_src_addr[3][4] ),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _4137_ (.A(net1250),
    .B(_2010_),
    .Y(_2017_));
 sky130_fd_sc_hd__o21ai_0 _4138_ (.A1(_0389_),
    .A2(_2010_),
    .B1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_1 _4139_ (.A(\current_src_addr[3][4] ),
    .B(_0389_),
    .Y(_2019_));
 sky130_fd_sc_hd__o22ai_1 _4140_ (.A1(net270),
    .A2(net1250),
    .B1(_2010_),
    .B2(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__a21oi_1 _4141_ (.A1(_2016_),
    .A2(_2018_),
    .B1(_2020_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand3_1 _4142_ (.A(\current_src_addr[3][2] ),
    .B(\current_src_addr[3][3] ),
    .C(\current_src_addr[3][4] ),
    .Y(_2021_));
 sky130_fd_sc_hd__a21oi_1 _4143_ (.A1(_2008_),
    .A2(_2021_),
    .B1(_2009_),
    .Y(_2022_));
 sky130_fd_sc_hd__nor2_1 _4144_ (.A(_2010_),
    .B(_2021_),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _4145_ (.A(\current_src_addr[3][5] ),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__o221a_2 _4146_ (.A1(net271),
    .A2(net1250),
    .B1(_2022_),
    .B2(\current_src_addr[3][5] ),
    .C1(_2024_),
    .X(_0247_));
 sky130_fd_sc_hd__nand3_1 _4147_ (.A(\current_src_addr[3][4] ),
    .B(_0389_),
    .C(\current_src_addr[3][5] ),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _4148_ (.A(_2008_),
    .B(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__a21oi_1 _4149_ (.A1(_2017_),
    .A2(_2026_),
    .B1(\current_src_addr[3][6] ),
    .Y(_2027_));
 sky130_fd_sc_hd__nand2_1 _4150_ (.A(\current_src_addr[3][5] ),
    .B(\current_src_addr[3][6] ),
    .Y(_2028_));
 sky130_fd_sc_hd__o32ai_1 _4151_ (.A1(_2010_),
    .A2(_2019_),
    .A3(_2028_),
    .B1(net1250),
    .B2(net272),
    .Y(_2029_));
 sky130_fd_sc_hd__nor2_1 _4152_ (.A(_2027_),
    .B(_2029_),
    .Y(_0248_));
 sky130_fd_sc_hd__o21ai_0 _4153_ (.A1(_2021_),
    .A2(_2028_),
    .B1(_2008_),
    .Y(_2030_));
 sky130_fd_sc_hd__a21oi_1 _4154_ (.A1(_2017_),
    .A2(_2030_),
    .B1(\current_src_addr[3][7] ),
    .Y(_2031_));
 sky130_fd_sc_hd__nand3_1 _4155_ (.A(\current_src_addr[3][5] ),
    .B(\current_src_addr[3][6] ),
    .C(\current_src_addr[3][7] ),
    .Y(_2032_));
 sky130_fd_sc_hd__or3_1 _4156_ (.A(_2010_),
    .B(_2021_),
    .C(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__o21ai_0 _4157_ (.A1(net273),
    .A2(net1250),
    .B1(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__nor2_1 _4158_ (.A(_2031_),
    .B(_2034_),
    .Y(_0249_));
 sky130_fd_sc_hd__or2_2 _4159_ (.A(_2019_),
    .B(_2032_),
    .X(_2035_));
 sky130_fd_sc_hd__a21oi_1 _4160_ (.A1(_2008_),
    .A2(_2035_),
    .B1(_2009_),
    .Y(_2036_));
 sky130_fd_sc_hd__nor2_1 _4161_ (.A(_2010_),
    .B(_2035_),
    .Y(_2037_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input136 (.A(channel_length[102]),
    .X(net136));
 sky130_fd_sc_hd__nand2_1 _4163_ (.A(\current_src_addr[3][8] ),
    .B(_2037_),
    .Y(_2039_));
 sky130_fd_sc_hd__o221a_2 _4164_ (.A1(net274),
    .A2(net1250),
    .B1(_2036_),
    .B2(\current_src_addr[3][8] ),
    .C1(_2039_),
    .X(_0250_));
 sky130_fd_sc_hd__nor4_4 _4165_ (.A(net268),
    .B(_1470_),
    .C(_2021_),
    .D(_2032_),
    .Y(_2040_));
 sky130_fd_sc_hd__nor2_1 _4166_ (.A(net275),
    .B(net1250),
    .Y(_2041_));
 sky130_fd_sc_hd__a211oi_1 _4167_ (.A1(\current_src_addr[3][8] ),
    .A2(_2040_),
    .B1(net1251),
    .C1(\current_src_addr[3][9] ),
    .Y(_2042_));
 sky130_fd_sc_hd__a311oi_1 _4168_ (.A1(\current_src_addr[3][8] ),
    .A2(\current_src_addr[3][9] ),
    .A3(_2040_),
    .B1(_2041_),
    .C1(_2042_),
    .Y(_0251_));
 sky130_fd_sc_hd__and3_1 _4169_ (.A(\current_src_addr[3][8] ),
    .B(\current_src_addr[3][9] ),
    .C(\current_src_addr[3][10] ),
    .X(_2043_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input135 (.A(channel_length[101]),
    .X(net135));
 sky130_fd_sc_hd__a311oi_1 _4171_ (.A1(\current_src_addr[3][8] ),
    .A2(\current_src_addr[3][9] ),
    .A3(_2037_),
    .B1(net1251),
    .C1(\current_src_addr[3][10] ),
    .Y(_2045_));
 sky130_fd_sc_hd__nor2_1 _4172_ (.A(net276),
    .B(net1250),
    .Y(_2046_));
 sky130_fd_sc_hd__a211oi_1 _4173_ (.A1(_2037_),
    .A2(_2043_),
    .B1(_2045_),
    .C1(_2046_),
    .Y(_0222_));
 sky130_fd_sc_hd__nor2_1 _4174_ (.A(net277),
    .B(net1250),
    .Y(_2047_));
 sky130_fd_sc_hd__a211oi_1 _4175_ (.A1(_2040_),
    .A2(_2043_),
    .B1(\current_src_addr[3][11] ),
    .C1(net1251),
    .Y(_2048_));
 sky130_fd_sc_hd__a311oi_1 _4176_ (.A1(\current_src_addr[3][11] ),
    .A2(_2040_),
    .A3(_2043_),
    .B1(_2047_),
    .C1(_2048_),
    .Y(_0223_));
 sky130_fd_sc_hd__and3_1 _4177_ (.A(\current_src_addr[3][11] ),
    .B(\current_src_addr[3][12] ),
    .C(_2043_),
    .X(_2049_));
 sky130_fd_sc_hd__a311oi_1 _4178_ (.A1(\current_src_addr[3][11] ),
    .A2(_2037_),
    .A3(_2043_),
    .B1(\current_src_addr[3][12] ),
    .C1(net1251),
    .Y(_2050_));
 sky130_fd_sc_hd__nor2_1 _4179_ (.A(net278),
    .B(net1250),
    .Y(_2051_));
 sky130_fd_sc_hd__a211oi_1 _4180_ (.A1(_2037_),
    .A2(_2049_),
    .B1(_2050_),
    .C1(_2051_),
    .Y(_0224_));
 sky130_fd_sc_hd__a211oi_1 _4181_ (.A1(_2040_),
    .A2(_2049_),
    .B1(\current_src_addr[3][13] ),
    .C1(net1251),
    .Y(_2052_));
 sky130_fd_sc_hd__nor2_1 _4182_ (.A(net279),
    .B(net1250),
    .Y(_2053_));
 sky130_fd_sc_hd__and3_1 _4183_ (.A(\current_src_addr[3][13] ),
    .B(_2040_),
    .C(_2049_),
    .X(_2054_));
 sky130_fd_sc_hd__nor3_1 _4184_ (.A(_2052_),
    .B(_2053_),
    .C(_2054_),
    .Y(_0225_));
 sky130_fd_sc_hd__and3_1 _4185_ (.A(\current_src_addr[3][11] ),
    .B(\current_src_addr[3][12] ),
    .C(\current_src_addr[3][13] ),
    .X(_2055_));
 sky130_fd_sc_hd__nand2_1 _4186_ (.A(_2043_),
    .B(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__o21ai_0 _4187_ (.A1(_2035_),
    .A2(_2056_),
    .B1(_2008_),
    .Y(_2057_));
 sky130_fd_sc_hd__a21oi_1 _4188_ (.A1(_2017_),
    .A2(_2057_),
    .B1(\current_src_addr[3][14] ),
    .Y(_2058_));
 sky130_fd_sc_hd__nand3_1 _4189_ (.A(\current_src_addr[3][14] ),
    .B(_2043_),
    .C(_2055_),
    .Y(_2059_));
 sky130_fd_sc_hd__o32ai_1 _4190_ (.A1(_2010_),
    .A2(_2035_),
    .A3(_2059_),
    .B1(net1250),
    .B2(net281),
    .Y(_2060_));
 sky130_fd_sc_hd__nor2_1 _4191_ (.A(_2058_),
    .B(_2060_),
    .Y(_0226_));
 sky130_fd_sc_hd__and4_1 _4192_ (.A(\current_src_addr[3][14] ),
    .B(\current_src_addr[3][15] ),
    .C(_2043_),
    .D(_2055_),
    .X(_2061_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input134 (.A(channel_length[100]),
    .X(net134));
 sky130_fd_sc_hd__nor2_1 _4194_ (.A(_2033_),
    .B(_2059_),
    .Y(_2063_));
 sky130_fd_sc_hd__nor3_1 _4195_ (.A(\current_src_addr[3][15] ),
    .B(net1251),
    .C(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__nor2_1 _4196_ (.A(net282),
    .B(net1250),
    .Y(_2065_));
 sky130_fd_sc_hd__a211oi_1 _4197_ (.A1(_2040_),
    .A2(_2061_),
    .B1(_2064_),
    .C1(_2065_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_1 _4198_ (.A(net283),
    .B(net1250),
    .Y(_2066_));
 sky130_fd_sc_hd__a211oi_1 _4199_ (.A1(_2037_),
    .A2(_2061_),
    .B1(\current_src_addr[3][16] ),
    .C1(net1251),
    .Y(_2067_));
 sky130_fd_sc_hd__a311oi_1 _4200_ (.A1(\current_src_addr[3][16] ),
    .A2(_2037_),
    .A3(_2061_),
    .B1(_2066_),
    .C1(_2067_),
    .Y(_0228_));
 sky130_fd_sc_hd__a41oi_1 _4201_ (.A1(\current_src_addr[3][14] ),
    .A2(\current_src_addr[3][15] ),
    .A3(\current_src_addr[3][16] ),
    .A4(_2054_),
    .B1(\current_src_addr[3][17] ),
    .Y(_2068_));
 sky130_fd_sc_hd__nor2_1 _4202_ (.A(net284),
    .B(net1250),
    .Y(_2069_));
 sky130_fd_sc_hd__and2_1 _4203_ (.A(\current_src_addr[3][16] ),
    .B(\current_src_addr[3][17] ),
    .X(_2070_));
 sky130_fd_sc_hd__and3_1 _4204_ (.A(_2040_),
    .B(_2061_),
    .C(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input133 (.A(channel_length[0]),
    .X(net133));
 sky130_fd_sc_hd__a211oi_1 _4206_ (.A1(net1250),
    .A2(_2068_),
    .B1(_2069_),
    .C1(_2071_),
    .Y(_0229_));
 sky130_fd_sc_hd__and2_1 _4207_ (.A(_2061_),
    .B(_2070_),
    .X(_2073_));
 sky130_fd_sc_hd__nand3_1 _4208_ (.A(\current_src_addr[3][18] ),
    .B(_2037_),
    .C(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__o21ai_0 _4209_ (.A1(net285),
    .A2(net1250),
    .B1(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__nor2_1 _4210_ (.A(_2019_),
    .B(_2032_),
    .Y(_2076_));
 sky130_fd_sc_hd__a211oi_1 _4211_ (.A1(_2076_),
    .A2(_2073_),
    .B1(\current_src_addr[3][18] ),
    .C1(_2010_),
    .Y(_2077_));
 sky130_fd_sc_hd__nor2_1 _4212_ (.A(\current_src_addr[3][18] ),
    .B(_2017_),
    .Y(_2078_));
 sky130_fd_sc_hd__nor3_1 _4213_ (.A(_2075_),
    .B(_2077_),
    .C(_2078_),
    .Y(_0230_));
 sky130_fd_sc_hd__nor2_1 _4214_ (.A(net286),
    .B(net1250),
    .Y(_2079_));
 sky130_fd_sc_hd__a211oi_1 _4215_ (.A1(\current_src_addr[3][18] ),
    .A2(_2071_),
    .B1(net1251),
    .C1(\current_src_addr[3][19] ),
    .Y(_2080_));
 sky130_fd_sc_hd__a311oi_1 _4216_ (.A1(\current_src_addr[3][18] ),
    .A2(\current_src_addr[3][19] ),
    .A3(_2071_),
    .B1(_2079_),
    .C1(_2080_),
    .Y(_0231_));
 sky130_fd_sc_hd__and2_1 _4217_ (.A(_2037_),
    .B(_2073_),
    .X(_2081_));
 sky130_fd_sc_hd__and3_1 _4218_ (.A(\current_src_addr[3][18] ),
    .B(\current_src_addr[3][19] ),
    .C(\current_src_addr[3][20] ),
    .X(_2082_));
 sky130_fd_sc_hd__a311oi_1 _4219_ (.A1(\current_src_addr[3][18] ),
    .A2(\current_src_addr[3][19] ),
    .A3(_2081_),
    .B1(net1251),
    .C1(\current_src_addr[3][20] ),
    .Y(_2083_));
 sky130_fd_sc_hd__nor2_1 _4220_ (.A(net287),
    .B(net1250),
    .Y(_2084_));
 sky130_fd_sc_hd__a211oi_1 _4221_ (.A1(_2081_),
    .A2(_2082_),
    .B1(_2083_),
    .C1(_2084_),
    .Y(_0232_));
 sky130_fd_sc_hd__nor2_1 _4222_ (.A(net288),
    .B(net1250),
    .Y(_2085_));
 sky130_fd_sc_hd__a211oi_1 _4223_ (.A1(_2071_),
    .A2(_2082_),
    .B1(\current_src_addr[3][21] ),
    .C1(net1251),
    .Y(_2086_));
 sky130_fd_sc_hd__a311oi_1 _4224_ (.A1(\current_src_addr[3][21] ),
    .A2(_2071_),
    .A3(_2082_),
    .B1(_2085_),
    .C1(_2086_),
    .Y(_0233_));
 sky130_fd_sc_hd__and3_1 _4225_ (.A(\current_src_addr[3][21] ),
    .B(\current_src_addr[3][22] ),
    .C(_2082_),
    .X(_2087_));
 sky130_fd_sc_hd__a311oi_1 _4226_ (.A1(\current_src_addr[3][21] ),
    .A2(_2081_),
    .A3(_2082_),
    .B1(\current_src_addr[3][22] ),
    .C1(net1251),
    .Y(_2088_));
 sky130_fd_sc_hd__nor2_1 _4227_ (.A(net289),
    .B(net1250),
    .Y(_2089_));
 sky130_fd_sc_hd__a211oi_1 _4228_ (.A1(_2081_),
    .A2(_2087_),
    .B1(_2088_),
    .C1(_2089_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand3_1 _4229_ (.A(_2061_),
    .B(_2070_),
    .C(_2087_),
    .Y(_2090_));
 sky130_fd_sc_hd__nor2_2 _4230_ (.A(_2033_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__nor3_1 _4231_ (.A(\current_src_addr[3][23] ),
    .B(net1251),
    .C(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nor2_1 _4232_ (.A(net290),
    .B(net1250),
    .Y(_2093_));
 sky130_fd_sc_hd__a211oi_1 _4233_ (.A1(\current_src_addr[3][23] ),
    .A2(_2091_),
    .B1(_2092_),
    .C1(_2093_),
    .Y(_0235_));
 sky130_fd_sc_hd__and3_1 _4234_ (.A(_2061_),
    .B(_2070_),
    .C(_2087_),
    .X(_2094_));
 sky130_fd_sc_hd__and2_1 _4235_ (.A(_2037_),
    .B(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__a211oi_1 _4236_ (.A1(\current_src_addr[3][23] ),
    .A2(_2095_),
    .B1(net1251),
    .C1(\current_src_addr[3][24] ),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _4237_ (.A(_2037_),
    .B(_2094_),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _4238_ (.A(\current_src_addr[3][23] ),
    .B(\current_src_addr[3][24] ),
    .Y(_2098_));
 sky130_fd_sc_hd__o22ai_1 _4239_ (.A1(net292),
    .A2(net1250),
    .B1(_2097_),
    .B2(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__nor2_1 _4240_ (.A(_2096_),
    .B(_2099_),
    .Y(_0236_));
 sky130_fd_sc_hd__and3_1 _4241_ (.A(\current_src_addr[3][23] ),
    .B(\current_src_addr[3][24] ),
    .C(\current_src_addr[3][25] ),
    .X(_2100_));
 sky130_fd_sc_hd__a311oi_1 _4242_ (.A1(\current_src_addr[3][23] ),
    .A2(\current_src_addr[3][24] ),
    .A3(_2091_),
    .B1(net1251),
    .C1(\current_src_addr[3][25] ),
    .Y(_2101_));
 sky130_fd_sc_hd__nor2_1 _4243_ (.A(net293),
    .B(net1250),
    .Y(_2102_));
 sky130_fd_sc_hd__a211oi_1 _4244_ (.A1(_2091_),
    .A2(_2100_),
    .B1(_2101_),
    .C1(_2102_),
    .Y(_0237_));
 sky130_fd_sc_hd__and2_1 _4245_ (.A(\current_src_addr[3][26] ),
    .B(_2100_),
    .X(_2103_));
 sky130_fd_sc_hd__a211oi_1 _4246_ (.A1(_2095_),
    .A2(_2100_),
    .B1(\current_src_addr[3][26] ),
    .C1(net1251),
    .Y(_2104_));
 sky130_fd_sc_hd__nor2_1 _4247_ (.A(net294),
    .B(net1250),
    .Y(_2105_));
 sky130_fd_sc_hd__a211oi_1 _4248_ (.A1(_2095_),
    .A2(_2103_),
    .B1(_2104_),
    .C1(_2105_),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_1 _4249_ (.A(net295),
    .B(net1250),
    .Y(_2106_));
 sky130_fd_sc_hd__a211oi_1 _4250_ (.A1(_2091_),
    .A2(_2103_),
    .B1(\current_src_addr[3][27] ),
    .C1(net1251),
    .Y(_2107_));
 sky130_fd_sc_hd__and3_1 _4251_ (.A(\current_src_addr[3][27] ),
    .B(_2091_),
    .C(_2103_),
    .X(_2108_));
 sky130_fd_sc_hd__nor3_1 _4252_ (.A(_2106_),
    .B(_2107_),
    .C(_2108_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(\current_src_addr[3][28] ),
    .B(_2008_),
    .Y(_2109_));
 sky130_fd_sc_hd__and3_1 _4254_ (.A(\current_src_addr[3][26] ),
    .B(\current_src_addr[3][27] ),
    .C(_2100_),
    .X(_2110_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(_2076_),
    .B(_2110_),
    .Y(_2111_));
 sky130_fd_sc_hd__o32ai_1 _4256_ (.A1(_2090_),
    .A2(_2109_),
    .A3(_2111_),
    .B1(net1250),
    .B2(net296),
    .Y(_2112_));
 sky130_fd_sc_hd__o21ai_0 _4257_ (.A1(_2090_),
    .A2(_2111_),
    .B1(_2008_),
    .Y(_2113_));
 sky130_fd_sc_hd__a21oi_1 _4258_ (.A1(_2017_),
    .A2(_2113_),
    .B1(\current_src_addr[3][28] ),
    .Y(_2114_));
 sky130_fd_sc_hd__nor2_1 _4259_ (.A(_2112_),
    .B(_2114_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand4_1 _4260_ (.A(\current_src_addr[3][28] ),
    .B(_2071_),
    .C(_2087_),
    .D(_2110_),
    .Y(_2115_));
 sky130_fd_sc_hd__nand2_1 _4261_ (.A(net297),
    .B(net1251),
    .Y(_2116_));
 sky130_fd_sc_hd__o21ai_0 _4262_ (.A1(\current_src_addr[3][29] ),
    .A2(_2115_),
    .B1(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__a31o_2 _4263_ (.A1(\current_src_addr[3][29] ),
    .A2(net1250),
    .A3(_2115_),
    .B1(_2117_),
    .X(_0241_));
 sky130_fd_sc_hd__nor2_1 _4264_ (.A(\current_src_addr[3][30] ),
    .B(net1251),
    .Y(_2118_));
 sky130_fd_sc_hd__nand4_1 _4265_ (.A(\current_src_addr[3][28] ),
    .B(\current_src_addr[3][29] ),
    .C(_2095_),
    .D(_2110_),
    .Y(_2119_));
 sky130_fd_sc_hd__nand4_1 _4266_ (.A(\current_src_addr[3][28] ),
    .B(\current_src_addr[3][29] ),
    .C(\current_src_addr[3][30] ),
    .D(_2110_),
    .Y(_2120_));
 sky130_fd_sc_hd__o22ai_1 _4267_ (.A1(net298),
    .A2(net1250),
    .B1(_2097_),
    .B2(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__a21oi_1 _4268_ (.A1(_2118_),
    .A2(_2119_),
    .B1(_2121_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _4269_ (.A(_2040_),
    .B(_2094_),
    .Y(_2122_));
 sky130_fd_sc_hd__nand2_1 _4270_ (.A(net299),
    .B(net1251),
    .Y(_2123_));
 sky130_fd_sc_hd__o211ai_1 _4271_ (.A1(_2122_),
    .A2(_2120_),
    .B1(\current_src_addr[3][31] ),
    .C1(net1250),
    .Y(_2124_));
 sky130_fd_sc_hd__o311ai_0 _4272_ (.A1(\current_src_addr[3][31] ),
    .A2(_2122_),
    .A3(_2120_),
    .B1(_2123_),
    .C1(_2124_),
    .Y(_0244_));
 sky130_fd_sc_hd__nor2_1 _4273_ (.A(net266),
    .B(net1266),
    .Y(_2125_));
 sky130_fd_sc_hd__nor2_1 _4274_ (.A(_1604_),
    .B(net1242),
    .Y(_2126_));
 sky130_fd_sc_hd__nand2b_1 _4275_ (.A_N(net266),
    .B(_1611_),
    .Y(_2127_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input132 (.A(channel_enable[3]),
    .X(net132));
 sky130_fd_sc_hd__nor2_1 _4277_ (.A(\current_src_addr[2][2] ),
    .B(_2127_),
    .Y(_2129_));
 sky130_fd_sc_hd__a221o_1 _4278_ (.A1(net359),
    .A2(net1249),
    .B1(_2126_),
    .B2(\current_src_addr[2][2] ),
    .C1(_2129_),
    .X(_0212_));
 sky130_fd_sc_hd__nand2_1 _4279_ (.A(net360),
    .B(net1249),
    .Y(_2130_));
 sky130_fd_sc_hd__nand2_1 _4280_ (.A(\current_src_addr[2][3] ),
    .B(net1248),
    .Y(_2131_));
 sky130_fd_sc_hd__nor2_1 _4281_ (.A(_0392_),
    .B(_2127_),
    .Y(_2132_));
 sky130_fd_sc_hd__a31oi_1 _4282_ (.A1(_2127_),
    .A2(_2130_),
    .A3(_2131_),
    .B1(_2132_),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_1 _4283_ (.A(\current_src_addr[2][4] ),
    .Y(_2133_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(net1248),
    .B(_2127_),
    .Y(_2134_));
 sky130_fd_sc_hd__o21ai_0 _4285_ (.A1(_0391_),
    .A2(_2127_),
    .B1(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(\current_src_addr[2][4] ),
    .B(_0391_),
    .Y(_2136_));
 sky130_fd_sc_hd__o22ai_1 _4287_ (.A1(net361),
    .A2(net1248),
    .B1(_2127_),
    .B2(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__a21oi_1 _4288_ (.A1(_2133_),
    .A2(_2135_),
    .B1(_2137_),
    .Y(_0216_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input131 (.A(channel_enable[2]),
    .X(net131));
 sky130_fd_sc_hd__nand3_1 _4290_ (.A(\current_src_addr[2][2] ),
    .B(\current_src_addr[2][3] ),
    .C(\current_src_addr[2][4] ),
    .Y(_2139_));
 sky130_fd_sc_hd__a21oi_1 _4291_ (.A1(net1242),
    .A2(_2139_),
    .B1(_2126_),
    .Y(_2140_));
 sky130_fd_sc_hd__nor2_1 _4292_ (.A(_2127_),
    .B(_2139_),
    .Y(_2141_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(\current_src_addr[2][5] ),
    .B(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__o221a_2 _4294_ (.A1(net362),
    .A2(net1248),
    .B1(_2140_),
    .B2(\current_src_addr[2][5] ),
    .C1(_2142_),
    .X(_0217_));
 sky130_fd_sc_hd__nand3_1 _4295_ (.A(\current_src_addr[2][4] ),
    .B(_0391_),
    .C(\current_src_addr[2][5] ),
    .Y(_2143_));
 sky130_fd_sc_hd__a21oi_1 _4296_ (.A1(net1242),
    .A2(_2143_),
    .B1(_2126_),
    .Y(_2144_));
 sky130_fd_sc_hd__nor2_1 _4297_ (.A(_2127_),
    .B(_2136_),
    .Y(_2145_));
 sky130_fd_sc_hd__nand3_1 _4298_ (.A(\current_src_addr[2][5] ),
    .B(\current_src_addr[2][6] ),
    .C(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__o221a_2 _4299_ (.A1(net364),
    .A2(net1248),
    .B1(_2144_),
    .B2(\current_src_addr[2][6] ),
    .C1(_2146_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _4300_ (.A(\current_src_addr[2][5] ),
    .B(\current_src_addr[2][6] ),
    .C(\current_src_addr[2][7] ),
    .X(_2147_));
 sky130_fd_sc_hd__nor2_1 _4301_ (.A(net365),
    .B(net1248),
    .Y(_2148_));
 sky130_fd_sc_hd__a311oi_1 _4302_ (.A1(\current_src_addr[2][5] ),
    .A2(\current_src_addr[2][6] ),
    .A3(_2141_),
    .B1(net1249),
    .C1(\current_src_addr[2][7] ),
    .Y(_2149_));
 sky130_fd_sc_hd__a211oi_1 _4303_ (.A1(_2141_),
    .A2(_2147_),
    .B1(_2148_),
    .C1(_2149_),
    .Y(_0219_));
 sky130_fd_sc_hd__nand3_1 _4304_ (.A(\current_src_addr[2][4] ),
    .B(_0391_),
    .C(_2147_),
    .Y(_2150_));
 sky130_fd_sc_hd__a21oi_1 _4305_ (.A1(net1242),
    .A2(_2150_),
    .B1(_2126_),
    .Y(_2151_));
 sky130_fd_sc_hd__nor2_1 _4306_ (.A(_2127_),
    .B(_2150_),
    .Y(_2152_));
 sky130_fd_sc_hd__nand2_1 _4307_ (.A(\current_src_addr[2][8] ),
    .B(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__o221a_2 _4308_ (.A1(net366),
    .A2(net1248),
    .B1(_2151_),
    .B2(\current_src_addr[2][8] ),
    .C1(_2153_),
    .X(_0220_));
 sky130_fd_sc_hd__nand3_1 _4309_ (.A(\current_src_addr[2][5] ),
    .B(\current_src_addr[2][6] ),
    .C(\current_src_addr[2][7] ),
    .Y(_2154_));
 sky130_fd_sc_hd__nor2_1 _4310_ (.A(_2139_),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__a21oi_1 _4311_ (.A1(\current_src_addr[2][8] ),
    .A2(_2155_),
    .B1(_2127_),
    .Y(_2156_));
 sky130_fd_sc_hd__nor2_1 _4312_ (.A(_2126_),
    .B(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__nand4_1 _4313_ (.A(\current_src_addr[2][8] ),
    .B(\current_src_addr[2][9] ),
    .C(net1242),
    .D(_2155_),
    .Y(_2158_));
 sky130_fd_sc_hd__o221a_2 _4314_ (.A1(net367),
    .A2(net1248),
    .B1(_2157_),
    .B2(\current_src_addr[2][9] ),
    .C1(_2158_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _4315_ (.A(\current_src_addr[2][8] ),
    .B(\current_src_addr[2][9] ),
    .C(\current_src_addr[2][10] ),
    .X(_2159_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input130 (.A(channel_enable[1]),
    .X(net130));
 sky130_fd_sc_hd__nor2_1 _4317_ (.A(net368),
    .B(net1248),
    .Y(_2161_));
 sky130_fd_sc_hd__a311oi_1 _4318_ (.A1(\current_src_addr[2][8] ),
    .A2(\current_src_addr[2][9] ),
    .A3(_2152_),
    .B1(net1249),
    .C1(\current_src_addr[2][10] ),
    .Y(_2162_));
 sky130_fd_sc_hd__a211oi_1 _4319_ (.A1(_2152_),
    .A2(_2159_),
    .B1(_2161_),
    .C1(_2162_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand2b_1 _4320_ (.A_N(_2139_),
    .B(_2147_),
    .Y(_2163_));
 sky130_fd_sc_hd__nor2_1 _4321_ (.A(_2127_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__a211oi_1 _4322_ (.A1(_2159_),
    .A2(_2164_),
    .B1(\current_src_addr[2][11] ),
    .C1(net1249),
    .Y(_2165_));
 sky130_fd_sc_hd__nor2_1 _4323_ (.A(net369),
    .B(net1248),
    .Y(_2166_));
 sky130_fd_sc_hd__a311oi_1 _4324_ (.A1(\current_src_addr[2][11] ),
    .A2(_2159_),
    .A3(_2164_),
    .B1(_2165_),
    .C1(_2166_),
    .Y(_0193_));
 sky130_fd_sc_hd__and3_1 _4325_ (.A(\current_src_addr[2][11] ),
    .B(\current_src_addr[2][12] ),
    .C(_2159_),
    .X(_2167_));
 sky130_fd_sc_hd__a311oi_1 _4326_ (.A1(\current_src_addr[2][11] ),
    .A2(_2152_),
    .A3(_2159_),
    .B1(\current_src_addr[2][12] ),
    .C1(net1249),
    .Y(_2168_));
 sky130_fd_sc_hd__nor2_1 _4327_ (.A(net370),
    .B(net1248),
    .Y(_2169_));
 sky130_fd_sc_hd__a211oi_1 _4328_ (.A1(_2152_),
    .A2(_2167_),
    .B1(_2168_),
    .C1(_2169_),
    .Y(_0194_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input129 (.A(channel_enable[0]),
    .X(net129));
 sky130_fd_sc_hd__a211oi_1 _4330_ (.A1(_2164_),
    .A2(_2167_),
    .B1(\current_src_addr[2][13] ),
    .C1(net1249),
    .Y(_2171_));
 sky130_fd_sc_hd__nand3_1 _4331_ (.A(\current_src_addr[2][13] ),
    .B(_2164_),
    .C(_2167_),
    .Y(_2172_));
 sky130_fd_sc_hd__o21ai_0 _4332_ (.A1(net371),
    .A2(net1248),
    .B1(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__nor2_1 _4333_ (.A(_2171_),
    .B(_2173_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand4_1 _4334_ (.A(\current_src_addr[2][11] ),
    .B(\current_src_addr[2][12] ),
    .C(\current_src_addr[2][13] ),
    .D(_2159_),
    .Y(_2174_));
 sky130_fd_sc_hd__or2_2 _4335_ (.A(_2150_),
    .B(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__a21oi_1 _4336_ (.A1(net1242),
    .A2(_2175_),
    .B1(_2126_),
    .Y(_2176_));
 sky130_fd_sc_hd__nor3_1 _4337_ (.A(_2127_),
    .B(_2150_),
    .C(_2174_),
    .Y(_2177_));
 sky130_fd_sc_hd__nand2_1 _4338_ (.A(\current_src_addr[2][14] ),
    .B(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__o221a_2 _4339_ (.A1(net372),
    .A2(net1248),
    .B1(_2176_),
    .B2(\current_src_addr[2][14] ),
    .C1(_2178_),
    .X(_0196_));
 sky130_fd_sc_hd__nor3_1 _4340_ (.A(_2127_),
    .B(_2163_),
    .C(_2174_),
    .Y(_2179_));
 sky130_fd_sc_hd__a211oi_1 _4341_ (.A1(\current_src_addr[2][14] ),
    .A2(_2179_),
    .B1(net1249),
    .C1(\current_src_addr[2][15] ),
    .Y(_2180_));
 sky130_fd_sc_hd__nor2_1 _4342_ (.A(net373),
    .B(net1248),
    .Y(_2181_));
 sky130_fd_sc_hd__a311oi_1 _4343_ (.A1(\current_src_addr[2][14] ),
    .A2(\current_src_addr[2][15] ),
    .A3(_2179_),
    .B1(_2180_),
    .C1(_2181_),
    .Y(_0197_));
 sky130_fd_sc_hd__a311oi_1 _4344_ (.A1(\current_src_addr[2][14] ),
    .A2(\current_src_addr[2][15] ),
    .A3(_2177_),
    .B1(net1249),
    .C1(\current_src_addr[2][16] ),
    .Y(_2182_));
 sky130_fd_sc_hd__nand4_1 _4345_ (.A(\current_src_addr[2][14] ),
    .B(\current_src_addr[2][15] ),
    .C(\current_src_addr[2][16] ),
    .D(_2177_),
    .Y(_2183_));
 sky130_fd_sc_hd__o21ai_0 _4346_ (.A1(net375),
    .A2(net1248),
    .B1(_2183_),
    .Y(_2184_));
 sky130_fd_sc_hd__nor2_1 _4347_ (.A(_2182_),
    .B(_2184_),
    .Y(_0198_));
 sky130_fd_sc_hd__and3_1 _4348_ (.A(\current_src_addr[2][14] ),
    .B(\current_src_addr[2][15] ),
    .C(\current_src_addr[2][16] ),
    .X(_2185_));
 sky130_fd_sc_hd__a211oi_1 _4349_ (.A1(_2179_),
    .A2(_2185_),
    .B1(\current_src_addr[2][17] ),
    .C1(net1249),
    .Y(_2186_));
 sky130_fd_sc_hd__nor2_1 _4350_ (.A(net376),
    .B(net1248),
    .Y(_2187_));
 sky130_fd_sc_hd__a311oi_1 _4351_ (.A1(\current_src_addr[2][17] ),
    .A2(_2179_),
    .A3(_2185_),
    .B1(_2186_),
    .C1(_2187_),
    .Y(_0199_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input128 (.A(net1588),
    .X(net128));
 sky130_fd_sc_hd__and2_1 _4353_ (.A(\current_src_addr[2][17] ),
    .B(_2185_),
    .X(_2189_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(\current_src_addr[2][17] ),
    .B(_2185_),
    .Y(_2190_));
 sky130_fd_sc_hd__o21ai_0 _4355_ (.A1(_2175_),
    .A2(_2190_),
    .B1(net1242),
    .Y(_2191_));
 sky130_fd_sc_hd__a21oi_1 _4356_ (.A1(_2134_),
    .A2(_2191_),
    .B1(\current_src_addr[2][18] ),
    .Y(_2192_));
 sky130_fd_sc_hd__nor2_1 _4357_ (.A(net377),
    .B(net1248),
    .Y(_2193_));
 sky130_fd_sc_hd__a311oi_1 _4358_ (.A1(\current_src_addr[2][18] ),
    .A2(_2177_),
    .A3(_2189_),
    .B1(_2192_),
    .C1(_2193_),
    .Y(_0200_));
 sky130_fd_sc_hd__a311oi_1 _4359_ (.A1(\current_src_addr[2][18] ),
    .A2(_2179_),
    .A3(_2189_),
    .B1(\current_src_addr[2][19] ),
    .C1(net1249),
    .Y(_2194_));
 sky130_fd_sc_hd__nand4_1 _4360_ (.A(\current_src_addr[2][18] ),
    .B(\current_src_addr[2][19] ),
    .C(_2179_),
    .D(_2189_),
    .Y(_2195_));
 sky130_fd_sc_hd__o21ai_0 _4361_ (.A1(net378),
    .A2(net1248),
    .B1(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(_2194_),
    .B(_2196_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor2_1 _4363_ (.A(net379),
    .B(net1248),
    .Y(_2197_));
 sky130_fd_sc_hd__nor4_2 _4364_ (.A(_2127_),
    .B(_2150_),
    .C(_2174_),
    .D(_2190_),
    .Y(_2198_));
 sky130_fd_sc_hd__a311oi_1 _4365_ (.A1(\current_src_addr[2][18] ),
    .A2(\current_src_addr[2][19] ),
    .A3(_2198_),
    .B1(net1249),
    .C1(\current_src_addr[2][20] ),
    .Y(_2199_));
 sky130_fd_sc_hd__and4_1 _4366_ (.A(\current_src_addr[2][18] ),
    .B(\current_src_addr[2][19] ),
    .C(\current_src_addr[2][20] ),
    .D(_2198_),
    .X(_2200_));
 sky130_fd_sc_hd__nor3_1 _4367_ (.A(_2197_),
    .B(_2199_),
    .C(_2200_),
    .Y(_0202_));
 sky130_fd_sc_hd__and3_1 _4368_ (.A(\current_src_addr[2][18] ),
    .B(\current_src_addr[2][19] ),
    .C(\current_src_addr[2][20] ),
    .X(_2201_));
 sky130_fd_sc_hd__a311oi_1 _4369_ (.A1(_2179_),
    .A2(_2189_),
    .A3(_2201_),
    .B1(net1249),
    .C1(\current_src_addr[2][21] ),
    .Y(_2202_));
 sky130_fd_sc_hd__nand4_1 _4370_ (.A(\current_src_addr[2][21] ),
    .B(_2179_),
    .C(_2189_),
    .D(_2201_),
    .Y(_2203_));
 sky130_fd_sc_hd__o21ai_0 _4371_ (.A1(net380),
    .A2(net1248),
    .B1(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__nor2_1 _4372_ (.A(_2202_),
    .B(_2204_),
    .Y(_0203_));
 sky130_fd_sc_hd__and4_1 _4373_ (.A(\current_src_addr[2][18] ),
    .B(\current_src_addr[2][19] ),
    .C(\current_src_addr[2][20] ),
    .D(\current_src_addr[2][21] ),
    .X(_2205_));
 sky130_fd_sc_hd__a211oi_1 _4374_ (.A1(_2198_),
    .A2(_2205_),
    .B1(\current_src_addr[2][22] ),
    .C1(net1249),
    .Y(_2206_));
 sky130_fd_sc_hd__nor2_1 _4375_ (.A(net381),
    .B(net1248),
    .Y(_2207_));
 sky130_fd_sc_hd__a311oi_1 _4376_ (.A1(\current_src_addr[2][22] ),
    .A2(_2198_),
    .A3(_2205_),
    .B1(_2206_),
    .C1(_2207_),
    .Y(_0204_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input127 (.A(net1373),
    .X(net127));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(\current_src_addr[2][22] ),
    .B(_2205_),
    .Y(_2209_));
 sky130_fd_sc_hd__nor4_1 _4379_ (.A(_2163_),
    .B(_2174_),
    .C(_2190_),
    .D(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__and2_1 _4380_ (.A(net1242),
    .B(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__or4_1 _4381_ (.A(_2163_),
    .B(_2174_),
    .C(_2190_),
    .D(_2209_),
    .X(_2212_));
 sky130_fd_sc_hd__a21oi_1 _4382_ (.A1(net1242),
    .A2(_2212_),
    .B1(_2126_),
    .Y(_2213_));
 sky130_fd_sc_hd__nor2_1 _4383_ (.A(\current_src_addr[2][23] ),
    .B(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__nor2_1 _4384_ (.A(net382),
    .B(net1248),
    .Y(_2215_));
 sky130_fd_sc_hd__a211oi_1 _4385_ (.A1(\current_src_addr[2][23] ),
    .A2(_2211_),
    .B1(_2214_),
    .C1(_2215_),
    .Y(_0205_));
 sky130_fd_sc_hd__and3_1 _4386_ (.A(\current_src_addr[2][22] ),
    .B(_2198_),
    .C(_2205_),
    .X(_2216_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input126 (.A(net1351),
    .X(net126));
 sky130_fd_sc_hd__a211oi_1 _4388_ (.A1(\current_src_addr[2][23] ),
    .A2(_2216_),
    .B1(net1249),
    .C1(\current_src_addr[2][24] ),
    .Y(_2218_));
 sky130_fd_sc_hd__nor2_1 _4389_ (.A(net383),
    .B(net1248),
    .Y(_2219_));
 sky130_fd_sc_hd__a311oi_1 _4390_ (.A1(\current_src_addr[2][23] ),
    .A2(\current_src_addr[2][24] ),
    .A3(_2216_),
    .B1(_2218_),
    .C1(_2219_),
    .Y(_0206_));
 sky130_fd_sc_hd__a311oi_1 _4391_ (.A1(\current_src_addr[2][23] ),
    .A2(\current_src_addr[2][24] ),
    .A3(_2211_),
    .B1(net1249),
    .C1(\current_src_addr[2][25] ),
    .Y(_2220_));
 sky130_fd_sc_hd__nand2_1 _4392_ (.A(net1242),
    .B(_2210_),
    .Y(_2221_));
 sky130_fd_sc_hd__nand3_1 _4393_ (.A(\current_src_addr[2][23] ),
    .B(\current_src_addr[2][24] ),
    .C(\current_src_addr[2][25] ),
    .Y(_2222_));
 sky130_fd_sc_hd__o22ai_1 _4394_ (.A1(net384),
    .A2(net1248),
    .B1(_2221_),
    .B2(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__nor2_1 _4395_ (.A(_2220_),
    .B(_2223_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand4_1 _4396_ (.A(\current_src_addr[2][23] ),
    .B(\current_src_addr[2][24] ),
    .C(\current_src_addr[2][25] ),
    .D(_2216_),
    .Y(_2224_));
 sky130_fd_sc_hd__nor2_1 _4397_ (.A(\current_src_addr[2][26] ),
    .B(net1249),
    .Y(_2225_));
 sky130_fd_sc_hd__and4_1 _4398_ (.A(\current_src_addr[2][23] ),
    .B(\current_src_addr[2][24] ),
    .C(\current_src_addr[2][25] ),
    .D(\current_src_addr[2][26] ),
    .X(_2226_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input125 (.A(net1348),
    .X(net125));
 sky130_fd_sc_hd__o2bb2ai_1 _4400_ (.A1_N(_2216_),
    .A2_N(_2226_),
    .B1(net386),
    .B2(net1248),
    .Y(_2228_));
 sky130_fd_sc_hd__a21oi_1 _4401_ (.A1(_2224_),
    .A2(_2225_),
    .B1(_2228_),
    .Y(_0208_));
 sky130_fd_sc_hd__a211oi_1 _4402_ (.A1(_2211_),
    .A2(_2226_),
    .B1(\current_src_addr[2][27] ),
    .C1(net1249),
    .Y(_2229_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(\current_src_addr[2][27] ),
    .B(_2226_),
    .Y(_2230_));
 sky130_fd_sc_hd__o22ai_1 _4404_ (.A1(net387),
    .A2(net1248),
    .B1(_2221_),
    .B2(_2230_),
    .Y(_2231_));
 sky130_fd_sc_hd__nor2_1 _4405_ (.A(_2229_),
    .B(_2231_),
    .Y(_0209_));
 sky130_fd_sc_hd__and3_1 _4406_ (.A(\current_src_addr[2][27] ),
    .B(\current_src_addr[2][28] ),
    .C(_2226_),
    .X(_2232_));
 sky130_fd_sc_hd__a311oi_1 _4407_ (.A1(\current_src_addr[2][27] ),
    .A2(_2216_),
    .A3(_2226_),
    .B1(\current_src_addr[2][28] ),
    .C1(net1249),
    .Y(_2233_));
 sky130_fd_sc_hd__nor2_1 _4408_ (.A(net388),
    .B(net1248),
    .Y(_2234_));
 sky130_fd_sc_hd__a211oi_1 _4409_ (.A1(_2216_),
    .A2(_2232_),
    .B1(_2233_),
    .C1(_2234_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand3_1 _4410_ (.A(\current_src_addr[2][27] ),
    .B(\current_src_addr[2][28] ),
    .C(_2226_),
    .Y(_2235_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(net389),
    .B(net1249),
    .Y(_2236_));
 sky130_fd_sc_hd__o211ai_1 _4412_ (.A1(_2221_),
    .A2(_2235_),
    .B1(\current_src_addr[2][29] ),
    .C1(net1248),
    .Y(_2237_));
 sky130_fd_sc_hd__o311ai_0 _4413_ (.A1(\current_src_addr[2][29] ),
    .A2(_2221_),
    .A3(_2235_),
    .B1(_2236_),
    .C1(_2237_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand3_1 _4414_ (.A(\current_src_addr[2][29] ),
    .B(\current_src_addr[2][30] ),
    .C(_2232_),
    .Y(_2238_));
 sky130_fd_sc_hd__inv_1 _4415_ (.A(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__a311oi_1 _4416_ (.A1(\current_src_addr[2][29] ),
    .A2(_2216_),
    .A3(_2232_),
    .B1(\current_src_addr[2][30] ),
    .C1(net1249),
    .Y(_2240_));
 sky130_fd_sc_hd__nor2_1 _4417_ (.A(net390),
    .B(net1248),
    .Y(_2241_));
 sky130_fd_sc_hd__a211oi_1 _4418_ (.A1(_2216_),
    .A2(_2239_),
    .B1(_2240_),
    .C1(_2241_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _4419_ (.A(net391),
    .B(net1248),
    .Y(_2242_));
 sky130_fd_sc_hd__nand2_1 _4420_ (.A(\current_src_addr[2][31] ),
    .B(net1242),
    .Y(_2243_));
 sky130_fd_sc_hd__nor3_1 _4421_ (.A(_2212_),
    .B(_2238_),
    .C(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__o21ai_0 _4422_ (.A1(_2212_),
    .A2(_2238_),
    .B1(net1242),
    .Y(_2245_));
 sky130_fd_sc_hd__a21oi_1 _4423_ (.A1(_2134_),
    .A2(_2245_),
    .B1(\current_src_addr[2][31] ),
    .Y(_2246_));
 sky130_fd_sc_hd__nor3_1 _4424_ (.A(_2242_),
    .B(_2244_),
    .C(_2246_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _4425_ (.A(net264),
    .B(net1265),
    .Y(_2247_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input124 (.A(net1338),
    .X(net124));
 sky130_fd_sc_hd__nor2_1 _4427_ (.A(net1247),
    .B(_2247_),
    .Y(_2249_));
 sky130_fd_sc_hd__nand2b_1 _4428_ (.A_N(net264),
    .B(_1741_),
    .Y(_2250_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input123 (.A(net1554),
    .X(net123));
 sky130_fd_sc_hd__nor2_1 _4430_ (.A(\current_src_addr[1][2] ),
    .B(_2250_),
    .Y(_2252_));
 sky130_fd_sc_hd__a221o_1 _4431_ (.A1(net324),
    .A2(net1247),
    .B1(_2249_),
    .B2(\current_src_addr[1][2] ),
    .C1(_2252_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _4432_ (.A(net325),
    .B(net1247),
    .Y(_2253_));
 sky130_fd_sc_hd__nand2_1 _4433_ (.A(\current_src_addr[1][3] ),
    .B(_1748_),
    .Y(_2254_));
 sky130_fd_sc_hd__nor2_1 _4434_ (.A(_0394_),
    .B(_2250_),
    .Y(_2255_));
 sky130_fd_sc_hd__a31oi_1 _4435_ (.A1(_2250_),
    .A2(_2253_),
    .A3(_2254_),
    .B1(_2255_),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_1 _4436_ (.A(\current_src_addr[1][4] ),
    .Y(_2256_));
 sky130_fd_sc_hd__nand2_1 _4437_ (.A(_1748_),
    .B(_2250_),
    .Y(_2257_));
 sky130_fd_sc_hd__o21ai_0 _4438_ (.A1(_0393_),
    .A2(_2250_),
    .B1(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__nand2_1 _4439_ (.A(\current_src_addr[1][4] ),
    .B(_0393_),
    .Y(_2259_));
 sky130_fd_sc_hd__o22ai_1 _4440_ (.A1(net326),
    .A2(_1748_),
    .B1(_2250_),
    .B2(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__a21oi_1 _4441_ (.A1(_2256_),
    .A2(_2258_),
    .B1(_2260_),
    .Y(_0186_));
 sky130_fd_sc_hd__nand3_1 _4442_ (.A(\current_src_addr[1][2] ),
    .B(\current_src_addr[1][3] ),
    .C(\current_src_addr[1][4] ),
    .Y(_2261_));
 sky130_fd_sc_hd__a21oi_1 _4443_ (.A1(_2247_),
    .A2(_2261_),
    .B1(_2249_),
    .Y(_2262_));
 sky130_fd_sc_hd__nor2_1 _4444_ (.A(_2250_),
    .B(_2261_),
    .Y(_2263_));
 sky130_fd_sc_hd__nand2_1 _4445_ (.A(\current_src_addr[1][5] ),
    .B(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__o221a_2 _4446_ (.A1(net327),
    .A2(_1748_),
    .B1(_2262_),
    .B2(\current_src_addr[1][5] ),
    .C1(_2264_),
    .X(_0187_));
 sky130_fd_sc_hd__nand3_1 _4447_ (.A(\current_src_addr[1][4] ),
    .B(_0393_),
    .C(\current_src_addr[1][5] ),
    .Y(_2265_));
 sky130_fd_sc_hd__a21oi_1 _4448_ (.A1(_2247_),
    .A2(_2265_),
    .B1(_2249_),
    .Y(_2266_));
 sky130_fd_sc_hd__nor2_1 _4449_ (.A(_2250_),
    .B(_2259_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand3_1 _4450_ (.A(\current_src_addr[1][5] ),
    .B(\current_src_addr[1][6] ),
    .C(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__o221a_2 _4451_ (.A1(net328),
    .A2(_1748_),
    .B1(_2266_),
    .B2(\current_src_addr[1][6] ),
    .C1(_2268_),
    .X(_0188_));
 sky130_fd_sc_hd__a311oi_1 _4452_ (.A1(\current_src_addr[1][5] ),
    .A2(\current_src_addr[1][6] ),
    .A3(_2263_),
    .B1(net1247),
    .C1(\current_src_addr[1][7] ),
    .Y(_2269_));
 sky130_fd_sc_hd__nand3_1 _4453_ (.A(\current_src_addr[1][5] ),
    .B(\current_src_addr[1][6] ),
    .C(\current_src_addr[1][7] ),
    .Y(_2270_));
 sky130_fd_sc_hd__o32ai_1 _4454_ (.A1(_2250_),
    .A2(_2261_),
    .A3(_2270_),
    .B1(_1748_),
    .B2(net329),
    .Y(_2271_));
 sky130_fd_sc_hd__nor2_1 _4455_ (.A(_2269_),
    .B(_2271_),
    .Y(_0189_));
 sky130_fd_sc_hd__or2_2 _4456_ (.A(_2259_),
    .B(_2270_),
    .X(_2272_));
 sky130_fd_sc_hd__a21oi_1 _4457_ (.A1(_2247_),
    .A2(_2272_),
    .B1(_2249_),
    .Y(_2273_));
 sky130_fd_sc_hd__nor2_1 _4458_ (.A(_2259_),
    .B(_2270_),
    .Y(_2274_));
 sky130_fd_sc_hd__nand3_1 _4459_ (.A(\current_src_addr[1][8] ),
    .B(_2247_),
    .C(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__o221a_2 _4460_ (.A1(net331),
    .A2(_1748_),
    .B1(_2273_),
    .B2(\current_src_addr[1][8] ),
    .C1(_2275_),
    .X(_0190_));
 sky130_fd_sc_hd__nor2_1 _4461_ (.A(net332),
    .B(_1748_),
    .Y(_2276_));
 sky130_fd_sc_hd__nor2_1 _4462_ (.A(_2261_),
    .B(_2270_),
    .Y(_2277_));
 sky130_fd_sc_hd__a311oi_1 _4463_ (.A1(\current_src_addr[1][8] ),
    .A2(_2247_),
    .A3(_2277_),
    .B1(\current_src_addr[1][9] ),
    .C1(net1247),
    .Y(_2278_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(\current_src_addr[1][8] ),
    .B(\current_src_addr[1][9] ),
    .Y(_2279_));
 sky130_fd_sc_hd__inv_1 _4465_ (.A(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__and3_1 _4466_ (.A(_2247_),
    .B(_2277_),
    .C(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__nor3_1 _4467_ (.A(_2276_),
    .B(_2278_),
    .C(_2281_),
    .Y(_0191_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input122 (.A(net1601),
    .X(net122));
 sky130_fd_sc_hd__nor3_1 _4469_ (.A(_2250_),
    .B(_2272_),
    .C(_2279_),
    .Y(_2283_));
 sky130_fd_sc_hd__o21ai_0 _4470_ (.A1(_2272_),
    .A2(_2279_),
    .B1(_2247_),
    .Y(_2284_));
 sky130_fd_sc_hd__a21oi_1 _4471_ (.A1(_2257_),
    .A2(_2284_),
    .B1(\current_src_addr[1][10] ),
    .Y(_2285_));
 sky130_fd_sc_hd__nor2_1 _4472_ (.A(net333),
    .B(net1245),
    .Y(_2286_));
 sky130_fd_sc_hd__a211oi_1 _4473_ (.A1(\current_src_addr[1][10] ),
    .A2(_2283_),
    .B1(_2285_),
    .C1(_2286_),
    .Y(_0162_));
 sky130_fd_sc_hd__and3_1 _4474_ (.A(_2247_),
    .B(_2277_),
    .C(_2280_),
    .X(_2287_));
 sky130_fd_sc_hd__a211oi_1 _4475_ (.A1(\current_src_addr[1][10] ),
    .A2(_2281_),
    .B1(net1247),
    .C1(\current_src_addr[1][11] ),
    .Y(_2288_));
 sky130_fd_sc_hd__nor2_1 _4476_ (.A(net334),
    .B(net1245),
    .Y(_2289_));
 sky130_fd_sc_hd__a311oi_1 _4477_ (.A1(\current_src_addr[1][10] ),
    .A2(\current_src_addr[1][11] ),
    .A3(_2287_),
    .B1(_2288_),
    .C1(_2289_),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_1 _4478_ (.A(net335),
    .B(net1245),
    .Y(_2290_));
 sky130_fd_sc_hd__a311oi_1 _4479_ (.A1(\current_src_addr[1][10] ),
    .A2(\current_src_addr[1][11] ),
    .A3(_2283_),
    .B1(net1247),
    .C1(\current_src_addr[1][12] ),
    .Y(_2291_));
 sky130_fd_sc_hd__and4_1 _4480_ (.A(\current_src_addr[1][10] ),
    .B(\current_src_addr[1][11] ),
    .C(\current_src_addr[1][12] ),
    .D(_2283_),
    .X(_2292_));
 sky130_fd_sc_hd__nor3_1 _4481_ (.A(_2290_),
    .B(_2291_),
    .C(_2292_),
    .Y(_0164_));
 sky130_fd_sc_hd__and4_1 _4482_ (.A(\current_src_addr[1][10] ),
    .B(\current_src_addr[1][11] ),
    .C(\current_src_addr[1][12] ),
    .D(\current_src_addr[1][13] ),
    .X(_2293_));
 sky130_fd_sc_hd__and3_1 _4483_ (.A(\current_src_addr[1][10] ),
    .B(\current_src_addr[1][11] ),
    .C(\current_src_addr[1][12] ),
    .X(_2294_));
 sky130_fd_sc_hd__a211oi_1 _4484_ (.A1(_2281_),
    .A2(_2294_),
    .B1(\current_src_addr[1][13] ),
    .C1(net1247),
    .Y(_2295_));
 sky130_fd_sc_hd__nor2_1 _4485_ (.A(net336),
    .B(net1245),
    .Y(_2296_));
 sky130_fd_sc_hd__a211oi_1 _4486_ (.A1(_2287_),
    .A2(_2293_),
    .B1(_2295_),
    .C1(_2296_),
    .Y(_0165_));
 sky130_fd_sc_hd__nor2_1 _4487_ (.A(net337),
    .B(net1245),
    .Y(_2297_));
 sky130_fd_sc_hd__a211oi_1 _4488_ (.A1(_2283_),
    .A2(_2293_),
    .B1(\current_src_addr[1][14] ),
    .C1(net1247),
    .Y(_2298_));
 sky130_fd_sc_hd__a311oi_1 _4489_ (.A1(\current_src_addr[1][14] ),
    .A2(_2283_),
    .A3(_2293_),
    .B1(_2297_),
    .C1(_2298_),
    .Y(_0166_));
 sky130_fd_sc_hd__and3_1 _4490_ (.A(\current_src_addr[1][14] ),
    .B(\current_src_addr[1][15] ),
    .C(_2293_),
    .X(_2299_));
 sky130_fd_sc_hd__a311oi_1 _4491_ (.A1(\current_src_addr[1][14] ),
    .A2(_2281_),
    .A3(_2293_),
    .B1(\current_src_addr[1][15] ),
    .C1(net1247),
    .Y(_2300_));
 sky130_fd_sc_hd__nor2_1 _4492_ (.A(net338),
    .B(net1245),
    .Y(_2301_));
 sky130_fd_sc_hd__a211oi_1 _4493_ (.A1(_2287_),
    .A2(_2299_),
    .B1(_2300_),
    .C1(_2301_),
    .Y(_0167_));
 sky130_fd_sc_hd__nor2_1 _4494_ (.A(net339),
    .B(_1748_),
    .Y(_2302_));
 sky130_fd_sc_hd__a211oi_1 _4495_ (.A1(_2283_),
    .A2(_2299_),
    .B1(\current_src_addr[1][16] ),
    .C1(net1247),
    .Y(_2303_));
 sky130_fd_sc_hd__a311oi_1 _4496_ (.A1(\current_src_addr[1][16] ),
    .A2(_2283_),
    .A3(_2299_),
    .B1(_2302_),
    .C1(_2303_),
    .Y(_0168_));
 sky130_fd_sc_hd__nor2_1 _4497_ (.A(_2250_),
    .B(_2279_),
    .Y(_2304_));
 sky130_fd_sc_hd__and3_1 _4498_ (.A(\current_src_addr[1][14] ),
    .B(\current_src_addr[1][15] ),
    .C(\current_src_addr[1][16] ),
    .X(_2305_));
 sky130_fd_sc_hd__and3_1 _4499_ (.A(\current_src_addr[1][17] ),
    .B(_2293_),
    .C(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__and3_1 _4500_ (.A(_2277_),
    .B(_2304_),
    .C(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__a311oi_1 _4501_ (.A1(\current_src_addr[1][16] ),
    .A2(_2287_),
    .A3(_2299_),
    .B1(\current_src_addr[1][17] ),
    .C1(net1247),
    .Y(_2308_));
 sky130_fd_sc_hd__nor2_1 _4502_ (.A(net340),
    .B(_1748_),
    .Y(_2309_));
 sky130_fd_sc_hd__nor3_1 _4503_ (.A(_2307_),
    .B(_2308_),
    .C(_2309_),
    .Y(_0169_));
 sky130_fd_sc_hd__a31oi_1 _4504_ (.A1(_2274_),
    .A2(_2280_),
    .A3(_2306_),
    .B1(_2250_),
    .Y(_2310_));
 sky130_fd_sc_hd__nor2_1 _4505_ (.A(_2249_),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__and3_1 _4506_ (.A(_2274_),
    .B(_2304_),
    .C(_2306_),
    .X(_2312_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(\current_src_addr[1][18] ),
    .B(_2312_),
    .Y(_2313_));
 sky130_fd_sc_hd__o221a_2 _4508_ (.A1(net342),
    .A2(net1245),
    .B1(_2311_),
    .B2(\current_src_addr[1][18] ),
    .C1(_2313_),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_1 _4509_ (.A(net343),
    .B(net1245),
    .Y(_2314_));
 sky130_fd_sc_hd__a211oi_1 _4510_ (.A1(\current_src_addr[1][18] ),
    .A2(_2307_),
    .B1(net1247),
    .C1(\current_src_addr[1][19] ),
    .Y(_2315_));
 sky130_fd_sc_hd__and3_1 _4511_ (.A(\current_src_addr[1][18] ),
    .B(\current_src_addr[1][19] ),
    .C(_2307_),
    .X(_2316_));
 sky130_fd_sc_hd__nor3_1 _4512_ (.A(_2314_),
    .B(_2315_),
    .C(_2316_),
    .Y(_0171_));
 sky130_fd_sc_hd__and3_1 _4513_ (.A(\current_src_addr[1][18] ),
    .B(\current_src_addr[1][19] ),
    .C(\current_src_addr[1][20] ),
    .X(_2317_));
 sky130_fd_sc_hd__a311oi_1 _4514_ (.A1(\current_src_addr[1][18] ),
    .A2(\current_src_addr[1][19] ),
    .A3(_2312_),
    .B1(net1247),
    .C1(\current_src_addr[1][20] ),
    .Y(_2318_));
 sky130_fd_sc_hd__nor2_1 _4515_ (.A(net344),
    .B(net1245),
    .Y(_2319_));
 sky130_fd_sc_hd__a211oi_1 _4516_ (.A1(_2312_),
    .A2(_2317_),
    .B1(_2318_),
    .C1(_2319_),
    .Y(_0172_));
 sky130_fd_sc_hd__nor2_1 _4517_ (.A(net345),
    .B(net1245),
    .Y(_2320_));
 sky130_fd_sc_hd__a211oi_1 _4518_ (.A1(_2307_),
    .A2(_2317_),
    .B1(\current_src_addr[1][21] ),
    .C1(net1247),
    .Y(_2321_));
 sky130_fd_sc_hd__a311oi_1 _4519_ (.A1(\current_src_addr[1][21] ),
    .A2(_2307_),
    .A3(_2317_),
    .B1(_2320_),
    .C1(_2321_),
    .Y(_0173_));
 sky130_fd_sc_hd__nor2_1 _4520_ (.A(net346),
    .B(net1245),
    .Y(_2322_));
 sky130_fd_sc_hd__a311oi_1 _4521_ (.A1(\current_src_addr[1][21] ),
    .A2(_2312_),
    .A3(_2317_),
    .B1(\current_src_addr[1][22] ),
    .C1(net1247),
    .Y(_2323_));
 sky130_fd_sc_hd__and4_1 _4522_ (.A(\current_src_addr[1][21] ),
    .B(\current_src_addr[1][22] ),
    .C(_2312_),
    .D(_2317_),
    .X(_2324_));
 sky130_fd_sc_hd__nor3_1 _4523_ (.A(_2322_),
    .B(_2323_),
    .C(_2324_),
    .Y(_0174_));
 sky130_fd_sc_hd__and3_1 _4524_ (.A(\current_src_addr[1][21] ),
    .B(\current_src_addr[1][22] ),
    .C(_2317_),
    .X(_2325_));
 sky130_fd_sc_hd__nand4_1 _4525_ (.A(_2277_),
    .B(_2280_),
    .C(_2306_),
    .D(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__nor2_1 _4526_ (.A(_2250_),
    .B(_2326_),
    .Y(_2327_));
 sky130_fd_sc_hd__a21oi_1 _4527_ (.A1(_2247_),
    .A2(_2326_),
    .B1(_2249_),
    .Y(_2328_));
 sky130_fd_sc_hd__nor2_1 _4528_ (.A(\current_src_addr[1][23] ),
    .B(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__nor2_1 _4529_ (.A(net347),
    .B(net1245),
    .Y(_2330_));
 sky130_fd_sc_hd__a211oi_1 _4530_ (.A1(\current_src_addr[1][23] ),
    .A2(_2327_),
    .B1(_2329_),
    .C1(_2330_),
    .Y(_0175_));
 sky130_fd_sc_hd__and4_1 _4531_ (.A(_2274_),
    .B(_2304_),
    .C(_2306_),
    .D(_2325_),
    .X(_2331_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input121 (.A(net1328),
    .X(net121));
 sky130_fd_sc_hd__a211oi_1 _4533_ (.A1(\current_src_addr[1][23] ),
    .A2(_2331_),
    .B1(net1247),
    .C1(\current_src_addr[1][24] ),
    .Y(_2333_));
 sky130_fd_sc_hd__nor2_1 _4534_ (.A(net348),
    .B(net1245),
    .Y(_2334_));
 sky130_fd_sc_hd__a311oi_1 _4535_ (.A1(\current_src_addr[1][23] ),
    .A2(\current_src_addr[1][24] ),
    .A3(_2331_),
    .B1(_2333_),
    .C1(_2334_),
    .Y(_0176_));
 sky130_fd_sc_hd__and3_1 _4536_ (.A(\current_src_addr[1][23] ),
    .B(\current_src_addr[1][24] ),
    .C(\current_src_addr[1][25] ),
    .X(_2335_));
 sky130_fd_sc_hd__nor2_1 _4537_ (.A(net349),
    .B(net1245),
    .Y(_2336_));
 sky130_fd_sc_hd__nand2_1 _4538_ (.A(\current_src_addr[1][23] ),
    .B(\current_src_addr[1][24] ),
    .Y(_2337_));
 sky130_fd_sc_hd__o21ai_0 _4539_ (.A1(_2326_),
    .A2(_2337_),
    .B1(_2247_),
    .Y(_2338_));
 sky130_fd_sc_hd__a21oi_1 _4540_ (.A1(_2257_),
    .A2(_2338_),
    .B1(\current_src_addr[1][25] ),
    .Y(_2339_));
 sky130_fd_sc_hd__a211oi_1 _4541_ (.A1(_2327_),
    .A2(_2335_),
    .B1(_2336_),
    .C1(_2339_),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_1 _4542_ (.A(net350),
    .B(net1245),
    .Y(_2340_));
 sky130_fd_sc_hd__a211oi_1 _4543_ (.A1(_2331_),
    .A2(_2335_),
    .B1(\current_src_addr[1][26] ),
    .C1(net1247),
    .Y(_2341_));
 sky130_fd_sc_hd__a311oi_1 _4544_ (.A1(\current_src_addr[1][26] ),
    .A2(_2331_),
    .A3(_2335_),
    .B1(_2340_),
    .C1(_2341_),
    .Y(_0178_));
 sky130_fd_sc_hd__and3_1 _4545_ (.A(\current_src_addr[1][26] ),
    .B(\current_src_addr[1][27] ),
    .C(_2335_),
    .X(_2342_));
 sky130_fd_sc_hd__a311oi_1 _4546_ (.A1(\current_src_addr[1][26] ),
    .A2(_2327_),
    .A3(_2335_),
    .B1(\current_src_addr[1][27] ),
    .C1(net1247),
    .Y(_2343_));
 sky130_fd_sc_hd__nor2_1 _4547_ (.A(net351),
    .B(net1245),
    .Y(_2344_));
 sky130_fd_sc_hd__a211oi_1 _4548_ (.A1(_2327_),
    .A2(_2342_),
    .B1(_2343_),
    .C1(_2344_),
    .Y(_0179_));
 sky130_fd_sc_hd__nor2_1 _4549_ (.A(net353),
    .B(net1245),
    .Y(_2345_));
 sky130_fd_sc_hd__a211oi_1 _4550_ (.A1(_2331_),
    .A2(_2342_),
    .B1(\current_src_addr[1][28] ),
    .C1(net1247),
    .Y(_2346_));
 sky130_fd_sc_hd__a311oi_1 _4551_ (.A1(\current_src_addr[1][28] ),
    .A2(_2331_),
    .A3(_2342_),
    .B1(_2345_),
    .C1(_2346_),
    .Y(_0180_));
 sky130_fd_sc_hd__and2_1 _4552_ (.A(\current_src_addr[1][28] ),
    .B(_2342_),
    .X(_2347_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(\current_src_addr[1][28] ),
    .B(_2342_),
    .Y(_2348_));
 sky130_fd_sc_hd__o21ai_0 _4554_ (.A1(_2326_),
    .A2(_2348_),
    .B1(_2247_),
    .Y(_2349_));
 sky130_fd_sc_hd__a21oi_1 _4555_ (.A1(_2257_),
    .A2(_2349_),
    .B1(\current_src_addr[1][29] ),
    .Y(_2350_));
 sky130_fd_sc_hd__nor2_1 _4556_ (.A(net354),
    .B(net1245),
    .Y(_2351_));
 sky130_fd_sc_hd__a311oi_1 _4557_ (.A1(\current_src_addr[1][29] ),
    .A2(_2327_),
    .A3(_2347_),
    .B1(_2350_),
    .C1(_2351_),
    .Y(_0181_));
 sky130_fd_sc_hd__and3_1 _4558_ (.A(\current_src_addr[1][29] ),
    .B(\current_src_addr[1][30] ),
    .C(_2347_),
    .X(_2352_));
 sky130_fd_sc_hd__a311oi_1 _4559_ (.A1(\current_src_addr[1][29] ),
    .A2(_2331_),
    .A3(_2347_),
    .B1(\current_src_addr[1][30] ),
    .C1(net1247),
    .Y(_2353_));
 sky130_fd_sc_hd__nor2_1 _4560_ (.A(net355),
    .B(net1245),
    .Y(_2354_));
 sky130_fd_sc_hd__a211oi_1 _4561_ (.A1(_2331_),
    .A2(_2352_),
    .B1(_2353_),
    .C1(_2354_),
    .Y(_0183_));
 sky130_fd_sc_hd__nor2_1 _4562_ (.A(net356),
    .B(net1245),
    .Y(_2355_));
 sky130_fd_sc_hd__a211oi_1 _4563_ (.A1(_2327_),
    .A2(_2352_),
    .B1(\current_src_addr[1][31] ),
    .C1(net1247),
    .Y(_2356_));
 sky130_fd_sc_hd__a311oi_1 _4564_ (.A1(\current_src_addr[1][31] ),
    .A2(_2327_),
    .A3(_2352_),
    .B1(_2355_),
    .C1(_2356_),
    .Y(_0184_));
 sky130_fd_sc_hd__nor2_1 _4565_ (.A(net262),
    .B(_1869_),
    .Y(_2357_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input120 (.A(net1312),
    .X(net120));
 sky130_fd_sc_hd__nor2_1 _4567_ (.A(_1866_),
    .B(_2357_),
    .Y(_2359_));
 sky130_fd_sc_hd__nand2b_1 _4568_ (.A_N(net262),
    .B(net1263),
    .Y(_2360_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(\current_src_addr[0][2] ),
    .B(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__a221o_1 _4570_ (.A1(net319),
    .A2(net1244),
    .B1(_2359_),
    .B2(\current_src_addr[0][2] ),
    .C1(_2361_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2i_1 _4571_ (.A0(\current_src_addr[0][3] ),
    .A1(net330),
    .S(net1244),
    .Y(_2362_));
 sky130_fd_sc_hd__nand2_1 _4572_ (.A(_0396_),
    .B(_2357_),
    .Y(_2363_));
 sky130_fd_sc_hd__o21ai_0 _4573_ (.A1(_2357_),
    .A2(_2362_),
    .B1(_2363_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(\current_src_addr[0][4] ),
    .B(_0395_),
    .Y(_2364_));
 sky130_fd_sc_hd__o22ai_1 _4575_ (.A1(net341),
    .A2(net1243),
    .B1(_2360_),
    .B2(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__nor2_1 _4576_ (.A(_0395_),
    .B(_2360_),
    .Y(_2366_));
 sky130_fd_sc_hd__nor2_1 _4577_ (.A(_2359_),
    .B(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__nor2_1 _4578_ (.A(\current_src_addr[0][4] ),
    .B(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__nor2_1 _4579_ (.A(_2365_),
    .B(_2368_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand3_1 _4580_ (.A(\current_src_addr[0][2] ),
    .B(\current_src_addr[0][3] ),
    .C(\current_src_addr[0][4] ),
    .Y(_2369_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(\current_src_addr[0][5] ),
    .B(_2357_),
    .Y(_2370_));
 sky130_fd_sc_hd__o22ai_1 _4582_ (.A1(net352),
    .A2(net1243),
    .B1(_2369_),
    .B2(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(net1243),
    .B(_2360_),
    .Y(_2372_));
 sky130_fd_sc_hd__nand2_1 _4584_ (.A(_2357_),
    .B(_2369_),
    .Y(_2373_));
 sky130_fd_sc_hd__a21oi_1 _4585_ (.A1(_2372_),
    .A2(_2373_),
    .B1(\current_src_addr[0][5] ),
    .Y(_2374_));
 sky130_fd_sc_hd__nor2_1 _4586_ (.A(_2371_),
    .B(_2374_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand3_1 _4587_ (.A(\current_src_addr[0][4] ),
    .B(_0395_),
    .C(\current_src_addr[0][5] ),
    .Y(_2375_));
 sky130_fd_sc_hd__nand2_1 _4588_ (.A(_2357_),
    .B(_2375_),
    .Y(_2376_));
 sky130_fd_sc_hd__a21oi_1 _4589_ (.A1(_2372_),
    .A2(_2376_),
    .B1(\current_src_addr[0][6] ),
    .Y(_2377_));
 sky130_fd_sc_hd__nand2_1 _4590_ (.A(\current_src_addr[0][5] ),
    .B(\current_src_addr[0][6] ),
    .Y(_2378_));
 sky130_fd_sc_hd__o32ai_1 _4591_ (.A1(_2360_),
    .A2(_2364_),
    .A3(_2378_),
    .B1(net1243),
    .B2(net363),
    .Y(_2379_));
 sky130_fd_sc_hd__nor2_1 _4592_ (.A(_2377_),
    .B(_2379_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand3_1 _4593_ (.A(\current_src_addr[0][5] ),
    .B(\current_src_addr[0][6] ),
    .C(\current_src_addr[0][7] ),
    .Y(_2380_));
 sky130_fd_sc_hd__nor4_1 _4594_ (.A(net262),
    .B(_1869_),
    .C(_2369_),
    .D(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__nor2_1 _4595_ (.A(net374),
    .B(_1880_),
    .Y(_2382_));
 sky130_fd_sc_hd__o21ai_0 _4596_ (.A1(_2369_),
    .A2(_2378_),
    .B1(_2357_),
    .Y(_2383_));
 sky130_fd_sc_hd__a21oi_1 _4597_ (.A1(_2372_),
    .A2(_2383_),
    .B1(\current_src_addr[0][7] ),
    .Y(_2384_));
 sky130_fd_sc_hd__nor3_1 _4598_ (.A(_2381_),
    .B(_2382_),
    .C(_2384_),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _4599_ (.A(_2364_),
    .B(_2380_),
    .Y(_2385_));
 sky130_fd_sc_hd__nor2_1 _4600_ (.A(_2360_),
    .B(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(_2359_),
    .B(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__nand3_1 _4602_ (.A(\current_src_addr[0][8] ),
    .B(_2357_),
    .C(_2385_),
    .Y(_2388_));
 sky130_fd_sc_hd__o221a_2 _4603_ (.A1(net385),
    .A2(net1243),
    .B1(_2387_),
    .B2(\current_src_addr[0][8] ),
    .C1(_2388_),
    .X(_0160_));
 sky130_fd_sc_hd__nor2_1 _4604_ (.A(net396),
    .B(net1243),
    .Y(_2389_));
 sky130_fd_sc_hd__a211oi_1 _4605_ (.A1(\current_src_addr[0][8] ),
    .A2(_2381_),
    .B1(net1244),
    .C1(\current_src_addr[0][9] ),
    .Y(_2390_));
 sky130_fd_sc_hd__and3_1 _4606_ (.A(\current_src_addr[0][8] ),
    .B(\current_src_addr[0][9] ),
    .C(_2381_),
    .X(_2391_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input119 (.A(net1548),
    .X(net119));
 sky130_fd_sc_hd__nor3_1 _4608_ (.A(_2389_),
    .B(_2390_),
    .C(_2391_),
    .Y(_0161_));
 sky130_fd_sc_hd__nor2_1 _4609_ (.A(net280),
    .B(net1243),
    .Y(_2393_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input118 (.A(net1521),
    .X(net118));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(\current_src_addr[0][8] ),
    .B(\current_src_addr[0][9] ),
    .Y(_2395_));
 sky130_fd_sc_hd__nor3_1 _4612_ (.A(_2364_),
    .B(_2380_),
    .C(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__nand2_1 _4613_ (.A(_2357_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__nor2_1 _4614_ (.A(_2360_),
    .B(_2396_),
    .Y(_2398_));
 sky130_fd_sc_hd__nor3_1 _4615_ (.A(\current_src_addr[0][10] ),
    .B(_2359_),
    .C(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__a21oi_1 _4616_ (.A1(\current_src_addr[0][10] ),
    .A2(_2397_),
    .B1(_2399_),
    .Y(_2400_));
 sky130_fd_sc_hd__nor2_1 _4617_ (.A(_2393_),
    .B(_2400_),
    .Y(_0132_));
 sky130_fd_sc_hd__nor2_1 _4618_ (.A(net291),
    .B(net1243),
    .Y(_2401_));
 sky130_fd_sc_hd__a211oi_1 _4619_ (.A1(\current_src_addr[0][10] ),
    .A2(_2391_),
    .B1(net1244),
    .C1(\current_src_addr[0][11] ),
    .Y(_2402_));
 sky130_fd_sc_hd__a311oi_1 _4620_ (.A1(\current_src_addr[0][10] ),
    .A2(\current_src_addr[0][11] ),
    .A3(_2391_),
    .B1(_2401_),
    .C1(_2402_),
    .Y(_0133_));
 sky130_fd_sc_hd__and2_1 _4621_ (.A(_2357_),
    .B(_2396_),
    .X(_2403_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input117 (.A(channel_dst_addr[8]),
    .X(net117));
 sky130_fd_sc_hd__a311oi_1 _4623_ (.A1(\current_src_addr[0][10] ),
    .A2(\current_src_addr[0][11] ),
    .A3(_2403_),
    .B1(net1244),
    .C1(\current_src_addr[0][12] ),
    .Y(_2405_));
 sky130_fd_sc_hd__a41oi_1 _4624_ (.A1(\current_src_addr[0][10] ),
    .A2(\current_src_addr[0][11] ),
    .A3(\current_src_addr[0][12] ),
    .A4(_2403_),
    .B1(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__o21a_1 _4625_ (.A1(net300),
    .A2(net1243),
    .B1(_2406_),
    .X(_0134_));
 sky130_fd_sc_hd__nor2_1 _4626_ (.A(\current_src_addr[0][13] ),
    .B(net1244),
    .Y(_2407_));
 sky130_fd_sc_hd__nand4_1 _4627_ (.A(\current_src_addr[0][10] ),
    .B(\current_src_addr[0][11] ),
    .C(\current_src_addr[0][12] ),
    .D(_2391_),
    .Y(_2408_));
 sky130_fd_sc_hd__and4_1 _4628_ (.A(\current_src_addr[0][10] ),
    .B(\current_src_addr[0][11] ),
    .C(\current_src_addr[0][12] ),
    .D(\current_src_addr[0][13] ),
    .X(_2409_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(_2391_),
    .B(_2409_),
    .Y(_2410_));
 sky130_fd_sc_hd__o21ai_0 _4630_ (.A1(net301),
    .A2(net1243),
    .B1(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__a21oi_1 _4631_ (.A1(_2407_),
    .A2(_2408_),
    .B1(_2411_),
    .Y(_0135_));
 sky130_fd_sc_hd__and2_1 _4632_ (.A(\current_src_addr[0][14] ),
    .B(_2409_),
    .X(_2412_));
 sky130_fd_sc_hd__a211oi_1 _4633_ (.A1(_2403_),
    .A2(_2409_),
    .B1(\current_src_addr[0][14] ),
    .C1(net1244),
    .Y(_2413_));
 sky130_fd_sc_hd__nor2_1 _4634_ (.A(net302),
    .B(net1243),
    .Y(_2414_));
 sky130_fd_sc_hd__a211oi_1 _4635_ (.A1(_2403_),
    .A2(_2412_),
    .B1(_2413_),
    .C1(_2414_),
    .Y(_0136_));
 sky130_fd_sc_hd__a211oi_1 _4636_ (.A1(_2391_),
    .A2(_2412_),
    .B1(\current_src_addr[0][15] ),
    .C1(net1244),
    .Y(_2415_));
 sky130_fd_sc_hd__a31oi_1 _4637_ (.A1(\current_src_addr[0][15] ),
    .A2(_2391_),
    .A3(_2412_),
    .B1(_2415_),
    .Y(_2416_));
 sky130_fd_sc_hd__o21a_1 _4638_ (.A1(net303),
    .A2(net1243),
    .B1(_2416_),
    .X(_0137_));
 sky130_fd_sc_hd__and3_1 _4639_ (.A(\current_src_addr[0][14] ),
    .B(\current_src_addr[0][15] ),
    .C(_2409_),
    .X(_2417_));
 sky130_fd_sc_hd__a211oi_1 _4640_ (.A1(_2403_),
    .A2(_2417_),
    .B1(\current_src_addr[0][16] ),
    .C1(net1244),
    .Y(_2418_));
 sky130_fd_sc_hd__nor2_1 _4641_ (.A(net304),
    .B(net1243),
    .Y(_2419_));
 sky130_fd_sc_hd__a311oi_1 _4642_ (.A1(\current_src_addr[0][16] ),
    .A2(_2403_),
    .A3(_2417_),
    .B1(_2418_),
    .C1(_2419_),
    .Y(_0138_));
 sky130_fd_sc_hd__nor2_1 _4643_ (.A(net305),
    .B(net1243),
    .Y(_2420_));
 sky130_fd_sc_hd__a311oi_1 _4644_ (.A1(\current_src_addr[0][16] ),
    .A2(_2391_),
    .A3(_2417_),
    .B1(\current_src_addr[0][17] ),
    .C1(net1244),
    .Y(_2421_));
 sky130_fd_sc_hd__and4_1 _4645_ (.A(\current_src_addr[0][16] ),
    .B(\current_src_addr[0][17] ),
    .C(_2391_),
    .D(_2417_),
    .X(_2422_));
 sky130_fd_sc_hd__nor3_1 _4646_ (.A(_2420_),
    .B(_2421_),
    .C(_2422_),
    .Y(_0139_));
 sky130_fd_sc_hd__and3_1 _4647_ (.A(\current_src_addr[0][15] ),
    .B(\current_src_addr[0][16] ),
    .C(\current_src_addr[0][17] ),
    .X(_2423_));
 sky130_fd_sc_hd__nand2_1 _4648_ (.A(_2412_),
    .B(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__nor2_1 _4649_ (.A(_2397_),
    .B(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__nand3_1 _4650_ (.A(_2396_),
    .B(_2412_),
    .C(_2423_),
    .Y(_2426_));
 sky130_fd_sc_hd__a21oi_1 _4651_ (.A1(_2357_),
    .A2(_2426_),
    .B1(_2359_),
    .Y(_2427_));
 sky130_fd_sc_hd__nor2_1 _4652_ (.A(\current_src_addr[0][18] ),
    .B(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__nor2_1 _4653_ (.A(net306),
    .B(net1243),
    .Y(_2429_));
 sky130_fd_sc_hd__a211oi_1 _4654_ (.A1(\current_src_addr[0][18] ),
    .A2(_2425_),
    .B1(_2428_),
    .C1(_2429_),
    .Y(_0140_));
 sky130_fd_sc_hd__nor2_1 _4655_ (.A(net307),
    .B(net1243),
    .Y(_2430_));
 sky130_fd_sc_hd__a211oi_1 _4656_ (.A1(\current_src_addr[0][18] ),
    .A2(_2422_),
    .B1(net1244),
    .C1(\current_src_addr[0][19] ),
    .Y(_2431_));
 sky130_fd_sc_hd__and3_1 _4657_ (.A(\current_src_addr[0][18] ),
    .B(\current_src_addr[0][19] ),
    .C(_2422_),
    .X(_2432_));
 sky130_fd_sc_hd__nor3_1 _4658_ (.A(_2430_),
    .B(_2431_),
    .C(_2432_),
    .Y(_0141_));
 sky130_fd_sc_hd__and3_1 _4659_ (.A(\current_src_addr[0][18] ),
    .B(\current_src_addr[0][19] ),
    .C(\current_src_addr[0][20] ),
    .X(_2433_));
 sky130_fd_sc_hd__a311oi_1 _4660_ (.A1(\current_src_addr[0][18] ),
    .A2(\current_src_addr[0][19] ),
    .A3(_2425_),
    .B1(net1244),
    .C1(\current_src_addr[0][20] ),
    .Y(_2434_));
 sky130_fd_sc_hd__nor2_1 _4661_ (.A(net309),
    .B(net1243),
    .Y(_2435_));
 sky130_fd_sc_hd__a211oi_1 _4662_ (.A1(_2425_),
    .A2(_2433_),
    .B1(_2434_),
    .C1(_2435_),
    .Y(_0142_));
 sky130_fd_sc_hd__nor2_1 _4663_ (.A(net310),
    .B(net1243),
    .Y(_2436_));
 sky130_fd_sc_hd__a211oi_1 _4664_ (.A1(_2422_),
    .A2(_2433_),
    .B1(\current_src_addr[0][21] ),
    .C1(net1244),
    .Y(_2437_));
 sky130_fd_sc_hd__a311oi_1 _4665_ (.A1(\current_src_addr[0][21] ),
    .A2(_2422_),
    .A3(_2433_),
    .B1(_2436_),
    .C1(_2437_),
    .Y(_0143_));
 sky130_fd_sc_hd__nor2_1 _4666_ (.A(net311),
    .B(net1243),
    .Y(_2438_));
 sky130_fd_sc_hd__a311oi_1 _4667_ (.A1(\current_src_addr[0][21] ),
    .A2(_2425_),
    .A3(_2433_),
    .B1(\current_src_addr[0][22] ),
    .C1(net1244),
    .Y(_2439_));
 sky130_fd_sc_hd__nand3_1 _4668_ (.A(\current_src_addr[0][21] ),
    .B(\current_src_addr[0][22] ),
    .C(_2433_),
    .Y(_2440_));
 sky130_fd_sc_hd__nor3_2 _4669_ (.A(_2397_),
    .B(_2424_),
    .C(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__nor3_1 _4670_ (.A(_2438_),
    .B(_2439_),
    .C(_2441_),
    .Y(_0144_));
 sky130_fd_sc_hd__nor2_1 _4671_ (.A(_2369_),
    .B(_2380_),
    .Y(_2442_));
 sky130_fd_sc_hd__nand4_1 _4672_ (.A(\current_src_addr[0][8] ),
    .B(\current_src_addr[0][9] ),
    .C(_2357_),
    .D(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__nor3_2 _4673_ (.A(_2443_),
    .B(_2424_),
    .C(_2440_),
    .Y(_2444_));
 sky130_fd_sc_hd__nor3_1 _4674_ (.A(\current_src_addr[0][23] ),
    .B(net1244),
    .C(net1229),
    .Y(_2445_));
 sky130_fd_sc_hd__nor2_1 _4675_ (.A(net312),
    .B(net1243),
    .Y(_2446_));
 sky130_fd_sc_hd__a211oi_1 _4676_ (.A1(\current_src_addr[0][23] ),
    .A2(net1229),
    .B1(_2445_),
    .C1(_2446_),
    .Y(_0145_));
 sky130_fd_sc_hd__nor2_1 _4677_ (.A(net313),
    .B(net1243),
    .Y(_2447_));
 sky130_fd_sc_hd__a211oi_1 _4678_ (.A1(\current_src_addr[0][23] ),
    .A2(net1228),
    .B1(net1244),
    .C1(\current_src_addr[0][24] ),
    .Y(_2448_));
 sky130_fd_sc_hd__a311oi_1 _4679_ (.A1(\current_src_addr[0][23] ),
    .A2(\current_src_addr[0][24] ),
    .A3(net1228),
    .B1(_2447_),
    .C1(_2448_),
    .Y(_0146_));
 sky130_fd_sc_hd__and3_1 _4680_ (.A(\current_src_addr[0][23] ),
    .B(\current_src_addr[0][24] ),
    .C(\current_src_addr[0][25] ),
    .X(_2449_));
 sky130_fd_sc_hd__a311oi_1 _4681_ (.A1(\current_src_addr[0][23] ),
    .A2(\current_src_addr[0][24] ),
    .A3(net1229),
    .B1(net1244),
    .C1(\current_src_addr[0][25] ),
    .Y(_2450_));
 sky130_fd_sc_hd__nor2_1 _4682_ (.A(net314),
    .B(net1243),
    .Y(_2451_));
 sky130_fd_sc_hd__a211oi_1 _4683_ (.A1(net1229),
    .A2(_2449_),
    .B1(_2450_),
    .C1(_2451_),
    .Y(_0147_));
 sky130_fd_sc_hd__nor2_1 _4684_ (.A(net315),
    .B(net1243),
    .Y(_2452_));
 sky130_fd_sc_hd__a211oi_1 _4685_ (.A1(net1228),
    .A2(_2449_),
    .B1(\current_src_addr[0][26] ),
    .C1(net1244),
    .Y(_2453_));
 sky130_fd_sc_hd__a311oi_1 _4686_ (.A1(\current_src_addr[0][26] ),
    .A2(net1228),
    .A3(_2449_),
    .B1(_2452_),
    .C1(_2453_),
    .Y(_0148_));
 sky130_fd_sc_hd__and3_1 _4687_ (.A(\current_src_addr[0][26] ),
    .B(\current_src_addr[0][27] ),
    .C(_2449_),
    .X(_2454_));
 sky130_fd_sc_hd__a311oi_1 _4688_ (.A1(\current_src_addr[0][26] ),
    .A2(net1229),
    .A3(_2449_),
    .B1(\current_src_addr[0][27] ),
    .C1(net1244),
    .Y(_2455_));
 sky130_fd_sc_hd__nor2_1 _4689_ (.A(net316),
    .B(net1243),
    .Y(_2456_));
 sky130_fd_sc_hd__a211oi_1 _4690_ (.A1(net1229),
    .A2(_2454_),
    .B1(_2455_),
    .C1(_2456_),
    .Y(_0149_));
 sky130_fd_sc_hd__nor2_1 _4691_ (.A(net317),
    .B(net1243),
    .Y(_2457_));
 sky130_fd_sc_hd__a211oi_1 _4692_ (.A1(net1228),
    .A2(_2454_),
    .B1(\current_src_addr[0][28] ),
    .C1(net1244),
    .Y(_2458_));
 sky130_fd_sc_hd__a311oi_1 _4693_ (.A1(\current_src_addr[0][28] ),
    .A2(net1228),
    .A3(_2454_),
    .B1(_2457_),
    .C1(_2458_),
    .Y(_0150_));
 sky130_fd_sc_hd__and3_1 _4694_ (.A(\current_src_addr[0][28] ),
    .B(\current_src_addr[0][29] ),
    .C(_2454_),
    .X(_2459_));
 sky130_fd_sc_hd__a311oi_1 _4695_ (.A1(\current_src_addr[0][28] ),
    .A2(net1229),
    .A3(_2454_),
    .B1(\current_src_addr[0][29] ),
    .C1(net1244),
    .Y(_2460_));
 sky130_fd_sc_hd__nor2_1 _4696_ (.A(net318),
    .B(net1243),
    .Y(_2461_));
 sky130_fd_sc_hd__a211oi_1 _4697_ (.A1(net1229),
    .A2(_2459_),
    .B1(_2460_),
    .C1(_2461_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor2_1 _4698_ (.A(net320),
    .B(net1243),
    .Y(_2462_));
 sky130_fd_sc_hd__a211oi_1 _4699_ (.A1(net1228),
    .A2(_2459_),
    .B1(\current_src_addr[0][30] ),
    .C1(net1244),
    .Y(_2463_));
 sky130_fd_sc_hd__a311oi_1 _4700_ (.A1(\current_src_addr[0][30] ),
    .A2(net1228),
    .A3(_2459_),
    .B1(_2462_),
    .C1(_2463_),
    .Y(_0153_));
 sky130_fd_sc_hd__nor2_1 _4701_ (.A(net321),
    .B(net1243),
    .Y(_2464_));
 sky130_fd_sc_hd__a311oi_1 _4702_ (.A1(\current_src_addr[0][30] ),
    .A2(net1229),
    .A3(_2459_),
    .B1(\current_src_addr[0][31] ),
    .C1(net1244),
    .Y(_2465_));
 sky130_fd_sc_hd__and4_1 _4703_ (.A(\current_src_addr[0][30] ),
    .B(\current_src_addr[0][31] ),
    .C(net1229),
    .D(_2459_),
    .X(_2466_));
 sky130_fd_sc_hd__nor3_1 _4704_ (.A(_2464_),
    .B(_2465_),
    .C(_2466_),
    .Y(_0154_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input116 (.A(net1404),
    .X(net116));
 sky130_fd_sc_hd__nor2_1 _4706_ (.A(_1465_),
    .B(net1267),
    .Y(_2468_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input115 (.A(net1314),
    .X(net115));
 sky130_fd_sc_hd__nand2_1 _4708_ (.A(net690),
    .B(net1234),
    .Y(_2470_));
 sky130_fd_sc_hd__o21ai_0 _4709_ (.A1(net690),
    .A2(net1268),
    .B1(_2470_),
    .Y(_0349_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input114 (.A(net1516),
    .X(net114));
 sky130_fd_sc_hd__nand2_1 _4711_ (.A(net691),
    .B(net1268),
    .Y(_2472_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input113 (.A(net1382),
    .X(net113));
 sky130_fd_sc_hd__nand2_1 _4713_ (.A(_0398_),
    .B(net1267),
    .Y(_2474_));
 sky130_fd_sc_hd__o21ai_0 _4714_ (.A1(_1465_),
    .A2(_2472_),
    .B1(_2474_),
    .Y(_0360_));
 sky130_fd_sc_hd__xor2_1 _4715_ (.A(net692),
    .B(_0397_),
    .X(_0670_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input112 (.A(net1431),
    .X(net112));
 sky130_fd_sc_hd__nand2_1 _4717_ (.A(_0397_),
    .B(net1267),
    .Y(_2476_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input111 (.A(net1313),
    .X(net111));
 sky130_fd_sc_hd__nor2_1 _4719_ (.A(_0397_),
    .B(net1268),
    .Y(_2478_));
 sky130_fd_sc_hd__o21ai_0 _4720_ (.A1(net1234),
    .A2(_2478_),
    .B1(net692),
    .Y(_2479_));
 sky130_fd_sc_hd__o21ai_0 _4721_ (.A1(net692),
    .A2(_2476_),
    .B1(_2479_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand3_1 _4722_ (.A(net690),
    .B(net691),
    .C(net692),
    .Y(_2480_));
 sky130_fd_sc_hd__xnor2_1 _4723_ (.A(net693),
    .B(_2480_),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(net1267),
    .B(_0666_),
    .Y(_2481_));
 sky130_fd_sc_hd__nand3_1 _4725_ (.A(net693),
    .B(_1473_),
    .C(net1268),
    .Y(_2482_));
 sky130_fd_sc_hd__nand2_1 _4726_ (.A(_2481_),
    .B(_2482_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand3_1 _4727_ (.A(net692),
    .B(_0397_),
    .C(net693),
    .Y(_2483_));
 sky130_fd_sc_hd__xnor2_1 _4728_ (.A(net568),
    .B(_2483_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(net1267),
    .B(_0686_),
    .Y(_2484_));
 sky130_fd_sc_hd__nand3_1 _4730_ (.A(net568),
    .B(_1473_),
    .C(net1268),
    .Y(_2485_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_2484_),
    .B(_2485_),
    .Y(_0375_));
 sky130_fd_sc_hd__and3_1 _4732_ (.A(net692),
    .B(net693),
    .C(net568),
    .X(_2486_));
 sky130_fd_sc_hd__nand3_1 _4733_ (.A(net690),
    .B(net691),
    .C(_2486_),
    .Y(_2487_));
 sky130_fd_sc_hd__xnor2_1 _4734_ (.A(net569),
    .B(_2487_),
    .Y(_0682_));
 sky130_fd_sc_hd__a31oi_1 _4735_ (.A1(net690),
    .A2(net691),
    .A3(_2486_),
    .B1(net1268),
    .Y(_2488_));
 sky130_fd_sc_hd__o21ai_0 _4736_ (.A1(net1234),
    .A2(_2488_),
    .B1(net569),
    .Y(_2489_));
 sky130_fd_sc_hd__o31ai_1 _4737_ (.A1(net569),
    .A2(net1268),
    .A3(_2487_),
    .B1(_2489_),
    .Y(_0376_));
 sky130_fd_sc_hd__and4_1 _4738_ (.A(net692),
    .B(_0397_),
    .C(net693),
    .D(net568),
    .X(_2490_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(net569),
    .B(_2490_),
    .Y(_2491_));
 sky130_fd_sc_hd__xnor2_1 _4740_ (.A(net570),
    .B(_2491_),
    .Y(_0678_));
 sky130_fd_sc_hd__a21oi_1 _4741_ (.A1(net569),
    .A2(_2490_),
    .B1(net1268),
    .Y(_2492_));
 sky130_fd_sc_hd__o21ai_0 _4742_ (.A1(net1234),
    .A2(_2492_),
    .B1(net570),
    .Y(_2493_));
 sky130_fd_sc_hd__o31ai_1 _4743_ (.A1(net570),
    .A2(net1268),
    .A3(_2491_),
    .B1(_2493_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_1 _4744_ (.A(net693),
    .B(net568),
    .Y(_2494_));
 sky130_fd_sc_hd__nand2_1 _4745_ (.A(net569),
    .B(net570),
    .Y(_2495_));
 sky130_fd_sc_hd__or3_1 _4746_ (.A(_2480_),
    .B(_2494_),
    .C(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input110 (.A(net1325),
    .X(net110));
 sky130_fd_sc_hd__xnor2_1 _4748_ (.A(net571),
    .B(_2496_),
    .Y(_0674_));
 sky130_fd_sc_hd__and2_1 _4749_ (.A(net1267),
    .B(_2496_),
    .X(_2498_));
 sky130_fd_sc_hd__o21ai_0 _4750_ (.A1(net1234),
    .A2(_2498_),
    .B1(net571),
    .Y(_2499_));
 sky130_fd_sc_hd__o31ai_1 _4751_ (.A1(net571),
    .A2(net1268),
    .A3(_2496_),
    .B1(_2499_),
    .Y(_0378_));
 sky130_fd_sc_hd__and2_1 _4752_ (.A(net569),
    .B(net570),
    .X(_2500_));
 sky130_fd_sc_hd__and3_1 _4753_ (.A(net571),
    .B(_2490_),
    .C(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__xor2_1 _4754_ (.A(net572),
    .B(_2501_),
    .X(_0718_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(net1267),
    .B(_2501_),
    .Y(_2502_));
 sky130_fd_sc_hd__nor2_1 _4756_ (.A(net1268),
    .B(_2501_),
    .Y(_2503_));
 sky130_fd_sc_hd__o21ai_0 _4757_ (.A1(net1234),
    .A2(_2503_),
    .B1(net572),
    .Y(_2504_));
 sky130_fd_sc_hd__o21ai_0 _4758_ (.A1(net572),
    .A2(_2502_),
    .B1(_2504_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(net571),
    .B(net572),
    .Y(_2505_));
 sky130_fd_sc_hd__nor4_1 _4760_ (.A(_2480_),
    .B(_2494_),
    .C(_2495_),
    .D(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__xor2_1 _4761_ (.A(net573),
    .B(_2506_),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(net1267),
    .B(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__nor2_1 _4763_ (.A(net1268),
    .B(_2506_),
    .Y(_2508_));
 sky130_fd_sc_hd__o21ai_0 _4764_ (.A1(net1234),
    .A2(_2508_),
    .B1(net573),
    .Y(_2509_));
 sky130_fd_sc_hd__o21ai_0 _4765_ (.A1(net573),
    .A2(_2507_),
    .B1(_2509_),
    .Y(_0380_));
 sky130_fd_sc_hd__and3_1 _4766_ (.A(net572),
    .B(net573),
    .C(_2501_),
    .X(_2510_));
 sky130_fd_sc_hd__xor2_1 _4767_ (.A(net574),
    .B(_2510_),
    .X(_0710_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(net1267),
    .B(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input109 (.A(net1309),
    .X(net109));
 sky130_fd_sc_hd__nand2_1 _4770_ (.A(_1473_),
    .B(net1268),
    .Y(_2513_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input108 (.A(net1300),
    .X(net108));
 sky130_fd_sc_hd__o21ai_0 _4772_ (.A1(net1268),
    .A2(_2510_),
    .B1(_2513_),
    .Y(_2515_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(net574),
    .B(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__o21ai_0 _4774_ (.A1(net574),
    .A2(_2511_),
    .B1(_2516_),
    .Y(_0350_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input107 (.A(net1409),
    .X(net107));
 sky130_fd_sc_hd__and3_1 _4776_ (.A(net573),
    .B(net574),
    .C(_2506_),
    .X(_2518_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input106 (.A(net1524),
    .X(net106));
 sky130_fd_sc_hd__xor2_1 _4778_ (.A(net575),
    .B(_2518_),
    .X(_0706_));
 sky130_fd_sc_hd__o21ai_0 _4779_ (.A1(net1268),
    .A2(_2518_),
    .B1(_2513_),
    .Y(_2520_));
 sky130_fd_sc_hd__nor2_1 _4780_ (.A(net575),
    .B(net1268),
    .Y(_2521_));
 sky130_fd_sc_hd__a22o_1 _4781_ (.A1(net575),
    .A2(_2520_),
    .B1(_2521_),
    .B2(_2518_),
    .X(_0351_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input105 (.A(net1381),
    .X(net105));
 sky130_fd_sc_hd__and4_1 _4783_ (.A(net571),
    .B(net572),
    .C(net573),
    .D(net574),
    .X(_2523_));
 sky130_fd_sc_hd__nand4_1 _4784_ (.A(net575),
    .B(_2490_),
    .C(_2500_),
    .D(_2523_),
    .Y(_2524_));
 sky130_fd_sc_hd__xnor2_1 _4785_ (.A(net576),
    .B(_2524_),
    .Y(_0702_));
 sky130_fd_sc_hd__and2_1 _4786_ (.A(net1267),
    .B(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__o21ai_0 _4787_ (.A1(net1234),
    .A2(_2525_),
    .B1(net576),
    .Y(_2526_));
 sky130_fd_sc_hd__o31ai_1 _4788_ (.A1(net576),
    .A2(net1268),
    .A3(_2524_),
    .B1(_2526_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand3_1 _4789_ (.A(net575),
    .B(net576),
    .C(_2518_),
    .Y(_2527_));
 sky130_fd_sc_hd__xnor2_1 _4790_ (.A(net577),
    .B(_2527_),
    .Y(_0698_));
 sky130_fd_sc_hd__a31oi_1 _4791_ (.A1(net575),
    .A2(net576),
    .A3(_2518_),
    .B1(net1268),
    .Y(_2528_));
 sky130_fd_sc_hd__o21ai_0 _4792_ (.A1(net1234),
    .A2(_2528_),
    .B1(net577),
    .Y(_2529_));
 sky130_fd_sc_hd__o31ai_1 _4793_ (.A1(net577),
    .A2(net1268),
    .A3(_2527_),
    .B1(_2529_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(net576),
    .B(net577),
    .Y(_2530_));
 sky130_fd_sc_hd__nor2_1 _4795_ (.A(_2524_),
    .B(_2530_),
    .Y(_2531_));
 sky130_fd_sc_hd__xor2_1 _4796_ (.A(net579),
    .B(_2531_),
    .X(_0694_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(net1267),
    .B(_2531_),
    .Y(_2532_));
 sky130_fd_sc_hd__o21ai_0 _4798_ (.A1(net1268),
    .A2(_2531_),
    .B1(_2513_),
    .Y(_2533_));
 sky130_fd_sc_hd__nand2_1 _4799_ (.A(net579),
    .B(_2533_),
    .Y(_2534_));
 sky130_fd_sc_hd__o21ai_0 _4800_ (.A1(net579),
    .A2(_2532_),
    .B1(_2534_),
    .Y(_0354_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input104 (.A(net1396),
    .X(net104));
 sky130_fd_sc_hd__and3_1 _4802_ (.A(net576),
    .B(net577),
    .C(net579),
    .X(_2536_));
 sky130_fd_sc_hd__nand3_1 _4803_ (.A(net575),
    .B(_2523_),
    .C(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__nor2_2 _4804_ (.A(_2496_),
    .B(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__xor2_1 _4805_ (.A(net580),
    .B(_2538_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(net1267),
    .B(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__o21ai_0 _4807_ (.A1(net1268),
    .A2(_2538_),
    .B1(_2513_),
    .Y(_2540_));
 sky130_fd_sc_hd__nand2_1 _4808_ (.A(net580),
    .B(_2540_),
    .Y(_2541_));
 sky130_fd_sc_hd__o21ai_0 _4809_ (.A1(net580),
    .A2(_2539_),
    .B1(_2541_),
    .Y(_0355_));
 sky130_fd_sc_hd__nand3_1 _4810_ (.A(net579),
    .B(net580),
    .C(_2531_),
    .Y(_2542_));
 sky130_fd_sc_hd__xnor2_1 _4811_ (.A(net581),
    .B(_2542_),
    .Y(_0782_));
 sky130_fd_sc_hd__a31oi_1 _4812_ (.A1(net579),
    .A2(net580),
    .A3(_2531_),
    .B1(net1268),
    .Y(_2543_));
 sky130_fd_sc_hd__o21ai_0 _4813_ (.A1(net1234),
    .A2(_2543_),
    .B1(net581),
    .Y(_2544_));
 sky130_fd_sc_hd__o31ai_1 _4814_ (.A1(net581),
    .A2(net1268),
    .A3(_2542_),
    .B1(_2544_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand3_1 _4815_ (.A(net580),
    .B(net581),
    .C(_2538_),
    .Y(_2545_));
 sky130_fd_sc_hd__xnor2_1 _4816_ (.A(net582),
    .B(_2545_),
    .Y(_0778_));
 sky130_fd_sc_hd__a31oi_1 _4817_ (.A1(net580),
    .A2(net581),
    .A3(_2538_),
    .B1(net1268),
    .Y(_2546_));
 sky130_fd_sc_hd__o21ai_0 _4818_ (.A1(net1234),
    .A2(_2546_),
    .B1(net582),
    .Y(_2547_));
 sky130_fd_sc_hd__o31ai_1 _4819_ (.A1(net582),
    .A2(net1268),
    .A3(_2545_),
    .B1(_2547_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand3_1 _4820_ (.A(net576),
    .B(net577),
    .C(net579),
    .Y(_2548_));
 sky130_fd_sc_hd__nand3_1 _4821_ (.A(net580),
    .B(net581),
    .C(net582),
    .Y(_2549_));
 sky130_fd_sc_hd__nor3_1 _4822_ (.A(_2524_),
    .B(_2548_),
    .C(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__xor2_1 _4823_ (.A(net583),
    .B(_2550_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _4824_ (.A(net1267),
    .B(_2550_),
    .Y(_2551_));
 sky130_fd_sc_hd__o21ai_0 _4825_ (.A1(net1268),
    .A2(_2550_),
    .B1(_2513_),
    .Y(_2552_));
 sky130_fd_sc_hd__nand2_1 _4826_ (.A(net583),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__o21ai_0 _4827_ (.A1(net583),
    .A2(_2551_),
    .B1(_2553_),
    .Y(_0358_));
 sky130_fd_sc_hd__and4_1 _4828_ (.A(net580),
    .B(net581),
    .C(net582),
    .D(net583),
    .X(_2554_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input103 (.A(net1344),
    .X(net103));
 sky130_fd_sc_hd__nand2_1 _4830_ (.A(_2538_),
    .B(_2554_),
    .Y(_2556_));
 sky130_fd_sc_hd__xnor2_1 _4831_ (.A(net584),
    .B(_2556_),
    .Y(_0770_));
 sky130_fd_sc_hd__a21oi_1 _4832_ (.A1(_2538_),
    .A2(_2554_),
    .B1(net1268),
    .Y(_2557_));
 sky130_fd_sc_hd__o21ai_0 _4833_ (.A1(net1234),
    .A2(_2557_),
    .B1(net584),
    .Y(_2558_));
 sky130_fd_sc_hd__o31ai_1 _4834_ (.A1(net584),
    .A2(net1268),
    .A3(_2556_),
    .B1(_2558_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _4835_ (.A(net584),
    .B(_2554_),
    .Y(_2559_));
 sky130_fd_sc_hd__nor3_1 _4836_ (.A(_2524_),
    .B(_2548_),
    .C(_2559_),
    .Y(_2560_));
 sky130_fd_sc_hd__xor2_1 _4837_ (.A(net585),
    .B(_2560_),
    .X(_0766_));
 sky130_fd_sc_hd__nand2_1 _4838_ (.A(net1267),
    .B(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__o21ai_0 _4839_ (.A1(net1268),
    .A2(_2560_),
    .B1(_2513_),
    .Y(_2562_));
 sky130_fd_sc_hd__nand2_1 _4840_ (.A(net585),
    .B(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__o21ai_0 _4841_ (.A1(net585),
    .A2(_2561_),
    .B1(_2563_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand4_1 _4842_ (.A(net584),
    .B(net585),
    .C(_2538_),
    .D(_2554_),
    .Y(_2564_));
 sky130_fd_sc_hd__xnor2_1 _4843_ (.A(net586),
    .B(_2564_),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_1 _4844_ (.A(net586),
    .Y(_2565_));
 sky130_fd_sc_hd__a21oi_1 _4845_ (.A1(net1267),
    .A2(_2564_),
    .B1(net1234),
    .Y(_2566_));
 sky130_fd_sc_hd__nor3_1 _4846_ (.A(net586),
    .B(net1268),
    .C(_2564_),
    .Y(_2567_));
 sky130_fd_sc_hd__o21bai_1 _4847_ (.A1(_2565_),
    .A2(_2566_),
    .B1_N(_2567_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand4_1 _4848_ (.A(net584),
    .B(net585),
    .C(net586),
    .D(_2554_),
    .Y(_2568_));
 sky130_fd_sc_hd__nor3_1 _4849_ (.A(_2524_),
    .B(_2548_),
    .C(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__xor2_1 _4850_ (.A(net587),
    .B(_2569_),
    .X(_0758_));
 sky130_fd_sc_hd__nand2_1 _4851_ (.A(net1267),
    .B(_2569_),
    .Y(_2570_));
 sky130_fd_sc_hd__o21ai_0 _4852_ (.A1(net1268),
    .A2(_2569_),
    .B1(_2513_),
    .Y(_2571_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(net587),
    .B(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__o21ai_0 _4854_ (.A1(net587),
    .A2(_2570_),
    .B1(_2572_),
    .Y(_0363_));
 sky130_fd_sc_hd__and4_1 _4855_ (.A(net584),
    .B(net585),
    .C(net586),
    .D(net587),
    .X(_2573_));
 sky130_fd_sc_hd__nand3_1 _4856_ (.A(_2538_),
    .B(_2554_),
    .C(_2573_),
    .Y(_2574_));
 sky130_fd_sc_hd__xnor2_1 _4857_ (.A(net588),
    .B(_2574_),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_1 _4858_ (.A(net588),
    .Y(_2575_));
 sky130_fd_sc_hd__a21oi_1 _4859_ (.A1(net1267),
    .A2(_2574_),
    .B1(net1234),
    .Y(_2576_));
 sky130_fd_sc_hd__nand2_1 _4860_ (.A(_2575_),
    .B(net1267),
    .Y(_2577_));
 sky130_fd_sc_hd__o22ai_1 _4861_ (.A1(_2575_),
    .A2(_2576_),
    .B1(_2577_),
    .B2(_2574_),
    .Y(_0364_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input102 (.A(net1399),
    .X(net102));
 sky130_fd_sc_hd__nand3_1 _4863_ (.A(net588),
    .B(_2554_),
    .C(_2573_),
    .Y(_2579_));
 sky130_fd_sc_hd__nor3_2 _4864_ (.A(_2524_),
    .B(_2548_),
    .C(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__xor2_1 _4865_ (.A(net590),
    .B(_2580_),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(net1267),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__o21ai_0 _4867_ (.A1(net1268),
    .A2(_2580_),
    .B1(_2513_),
    .Y(_2582_));
 sky130_fd_sc_hd__nand2_1 _4868_ (.A(net590),
    .B(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__o21ai_0 _4869_ (.A1(net590),
    .A2(_2581_),
    .B1(_2583_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor3_1 _4870_ (.A(_2496_),
    .B(_2537_),
    .C(_2579_),
    .Y(_2584_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(net590),
    .B(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__xnor2_1 _4872_ (.A(net591),
    .B(_2585_),
    .Y(_0746_));
 sky130_fd_sc_hd__a21oi_1 _4873_ (.A1(net590),
    .A2(_2584_),
    .B1(net1268),
    .Y(_2586_));
 sky130_fd_sc_hd__o21ai_0 _4874_ (.A1(net1234),
    .A2(_2586_),
    .B1(net591),
    .Y(_2587_));
 sky130_fd_sc_hd__o31ai_1 _4875_ (.A1(net591),
    .A2(net1268),
    .A3(_2585_),
    .B1(_2587_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand3_1 _4876_ (.A(net590),
    .B(net591),
    .C(_2580_),
    .Y(_2588_));
 sky130_fd_sc_hd__xnor2_1 _4877_ (.A(net592),
    .B(_2588_),
    .Y(_0742_));
 sky130_fd_sc_hd__a31oi_1 _4878_ (.A1(net590),
    .A2(net591),
    .A3(_2580_),
    .B1(net1268),
    .Y(_2589_));
 sky130_fd_sc_hd__o21ai_0 _4879_ (.A1(net1234),
    .A2(_2589_),
    .B1(net592),
    .Y(_2590_));
 sky130_fd_sc_hd__o31ai_1 _4880_ (.A1(net592),
    .A2(net1268),
    .A3(_2588_),
    .B1(_2590_),
    .Y(_0367_));
 sky130_fd_sc_hd__and4_1 _4881_ (.A(net590),
    .B(net591),
    .C(net592),
    .D(_2584_),
    .X(_2591_));
 sky130_fd_sc_hd__xor2_1 _4882_ (.A(net593),
    .B(_2591_),
    .X(_0738_));
 sky130_fd_sc_hd__nand2b_1 _4883_ (.A_N(_2591_),
    .B(net1267),
    .Y(_2592_));
 sky130_fd_sc_hd__a21oi_1 _4884_ (.A1(net1267),
    .A2(_2591_),
    .B1(net593),
    .Y(_2593_));
 sky130_fd_sc_hd__a31oi_1 _4885_ (.A1(net593),
    .A2(_2513_),
    .A3(_2592_),
    .B1(_2593_),
    .Y(_0368_));
 sky130_fd_sc_hd__and4_1 _4886_ (.A(net590),
    .B(net591),
    .C(net592),
    .D(net593),
    .X(_2594_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(_2580_),
    .B(_2594_),
    .Y(_2595_));
 sky130_fd_sc_hd__xnor2_1 _4888_ (.A(net594),
    .B(_2595_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_1 _4889_ (.A1(_2580_),
    .A2(_2594_),
    .B1(net1268),
    .Y(_2596_));
 sky130_fd_sc_hd__o21ai_0 _4890_ (.A1(net1234),
    .A2(_2596_),
    .B1(net594),
    .Y(_2597_));
 sky130_fd_sc_hd__o31ai_1 _4891_ (.A1(net594),
    .A2(net1268),
    .A3(_2595_),
    .B1(_2597_),
    .Y(_0369_));
 sky130_fd_sc_hd__and3_1 _4892_ (.A(net594),
    .B(_2584_),
    .C(_2594_),
    .X(_2598_));
 sky130_fd_sc_hd__xor2_1 _4893_ (.A(net595),
    .B(_2598_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2b_1 _4894_ (.A_N(_2598_),
    .B(net1267),
    .Y(_2599_));
 sky130_fd_sc_hd__a21oi_1 _4895_ (.A1(net1267),
    .A2(_2598_),
    .B1(net595),
    .Y(_2600_));
 sky130_fd_sc_hd__a31oi_1 _4896_ (.A1(net595),
    .A2(_2513_),
    .A3(_2599_),
    .B1(_2600_),
    .Y(_0370_));
 sky130_fd_sc_hd__and3_1 _4897_ (.A(net594),
    .B(net595),
    .C(_2594_),
    .X(_2601_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_2580_),
    .B(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__xnor2_1 _4899_ (.A(net596),
    .B(_2602_),
    .Y(_0726_));
 sky130_fd_sc_hd__a21oi_1 _4900_ (.A1(_2580_),
    .A2(_2601_),
    .B1(net1268),
    .Y(_2603_));
 sky130_fd_sc_hd__o21ai_0 _4901_ (.A1(net1234),
    .A2(_2603_),
    .B1(net596),
    .Y(_2604_));
 sky130_fd_sc_hd__o31ai_1 _4902_ (.A1(net596),
    .A2(net1268),
    .A3(_2602_),
    .B1(_2604_),
    .Y(_0372_));
 sky130_fd_sc_hd__and3_1 _4903_ (.A(net596),
    .B(_2584_),
    .C(_2601_),
    .X(_2605_));
 sky130_fd_sc_hd__xor2_1 _4904_ (.A(net597),
    .B(_2605_),
    .X(_0722_));
 sky130_fd_sc_hd__nand2b_1 _4905_ (.A_N(_2605_),
    .B(net1267),
    .Y(_2606_));
 sky130_fd_sc_hd__a21oi_1 _4906_ (.A1(net1267),
    .A2(_2605_),
    .B1(net597),
    .Y(_2607_));
 sky130_fd_sc_hd__a31oi_1 _4907_ (.A1(net597),
    .A2(_2513_),
    .A3(_2606_),
    .B1(_2607_),
    .Y(_0373_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input101 (.A(net1377),
    .X(net101));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input100 (.A(net1484),
    .X(net100));
 sky130_fd_sc_hd__nor2_2 _4910_ (.A(_1604_),
    .B(_1611_),
    .Y(_2610_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input99 (.A(net1503),
    .X(net99));
 sky130_fd_sc_hd__nand2_1 _4912_ (.A(net655),
    .B(net1233),
    .Y(_2612_));
 sky130_fd_sc_hd__o21ai_0 _4913_ (.A1(net655),
    .A2(net1266),
    .B1(_2612_),
    .Y(_0317_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input98 (.A(net1310),
    .X(net98));
 sky130_fd_sc_hd__nand2_1 _4915_ (.A(net656),
    .B(net1266),
    .Y(_2614_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input97 (.A(net1376),
    .X(net97));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_0400_),
    .B(_1611_),
    .Y(_2616_));
 sky130_fd_sc_hd__o21ai_0 _4918_ (.A1(_1604_),
    .A2(_2614_),
    .B1(_2616_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_1 _4919_ (.A(net657),
    .B(_0399_),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(_0399_),
    .B(_1611_),
    .Y(_2617_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input96 (.A(net1427),
    .X(net96));
 sky130_fd_sc_hd__nor2_1 _4922_ (.A(_0399_),
    .B(net1266),
    .Y(_2619_));
 sky130_fd_sc_hd__o21ai_0 _4923_ (.A1(_2610_),
    .A2(_2619_),
    .B1(net657),
    .Y(_2620_));
 sky130_fd_sc_hd__o21ai_0 _4924_ (.A1(net657),
    .A2(_2617_),
    .B1(_2620_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand3_1 _4925_ (.A(net655),
    .B(net656),
    .C(net657),
    .Y(_2621_));
 sky130_fd_sc_hd__xnor2_1 _4926_ (.A(net658),
    .B(_2621_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _4927_ (.A(_1611_),
    .B(_0791_),
    .Y(_2622_));
 sky130_fd_sc_hd__nand3_1 _4928_ (.A(net658),
    .B(_1618_),
    .C(net1266),
    .Y(_2623_));
 sky130_fd_sc_hd__nand2_1 _4929_ (.A(_2622_),
    .B(_2623_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand3_1 _4930_ (.A(net657),
    .B(_0399_),
    .C(net658),
    .Y(_2624_));
 sky130_fd_sc_hd__xnor2_1 _4931_ (.A(net659),
    .B(_2624_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_1611_),
    .B(_0811_),
    .Y(_2625_));
 sky130_fd_sc_hd__nand3_1 _4933_ (.A(net659),
    .B(_1618_),
    .C(net1266),
    .Y(_2626_));
 sky130_fd_sc_hd__nand2_1 _4934_ (.A(_2625_),
    .B(_2626_),
    .Y(_0343_));
 sky130_fd_sc_hd__and3_1 _4935_ (.A(net657),
    .B(net658),
    .C(net659),
    .X(_2627_));
 sky130_fd_sc_hd__nand3_1 _4936_ (.A(net655),
    .B(net656),
    .C(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__xnor2_1 _4937_ (.A(net660),
    .B(_2628_),
    .Y(_0807_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input95 (.A(net1625),
    .X(net95));
 sky130_fd_sc_hd__a31oi_1 _4939_ (.A1(net655),
    .A2(net656),
    .A3(_2627_),
    .B1(net1266),
    .Y(_2630_));
 sky130_fd_sc_hd__o21ai_0 _4940_ (.A1(net1233),
    .A2(_2630_),
    .B1(net660),
    .Y(_2631_));
 sky130_fd_sc_hd__o31ai_1 _4941_ (.A1(net660),
    .A2(net1266),
    .A3(_2628_),
    .B1(_2631_),
    .Y(_0344_));
 sky130_fd_sc_hd__and4_1 _4942_ (.A(net657),
    .B(_0399_),
    .C(net658),
    .D(net659),
    .X(_2632_));
 sky130_fd_sc_hd__and2_1 _4943_ (.A(net660),
    .B(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__xor2_1 _4944_ (.A(net662),
    .B(_2633_),
    .X(_0803_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(_1611_),
    .B(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__nor2_1 _4946_ (.A(net1266),
    .B(_2633_),
    .Y(_2635_));
 sky130_fd_sc_hd__o21ai_0 _4947_ (.A1(net1233),
    .A2(_2635_),
    .B1(net662),
    .Y(_2636_));
 sky130_fd_sc_hd__o21ai_0 _4948_ (.A1(net662),
    .A2(_2634_),
    .B1(_2636_),
    .Y(_0345_));
 sky130_fd_sc_hd__and2_1 _4949_ (.A(net660),
    .B(net662),
    .X(_2637_));
 sky130_fd_sc_hd__nand4_1 _4950_ (.A(net655),
    .B(net656),
    .C(_2627_),
    .D(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__xnor2_1 _4951_ (.A(net1270),
    .B(net1241),
    .Y(_0799_));
 sky130_fd_sc_hd__and4_1 _4952_ (.A(net655),
    .B(net656),
    .C(_2627_),
    .D(_2637_),
    .X(_2639_));
 sky130_fd_sc_hd__nor2_1 _4953_ (.A(net1266),
    .B(_2639_),
    .Y(_2640_));
 sky130_fd_sc_hd__o21ai_0 _4954_ (.A1(net1233),
    .A2(_2640_),
    .B1(net1270),
    .Y(_2641_));
 sky130_fd_sc_hd__o31ai_1 _4955_ (.A1(net1270),
    .A2(net1266),
    .A3(net1241),
    .B1(_2641_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand3_1 _4956_ (.A(net1270),
    .B(_2632_),
    .C(_2637_),
    .Y(_2642_));
 sky130_fd_sc_hd__xnor2_1 _4957_ (.A(net664),
    .B(_2642_),
    .Y(_0843_));
 sky130_fd_sc_hd__and3_1 _4958_ (.A(net1270),
    .B(_2632_),
    .C(_2637_),
    .X(_2643_));
 sky130_fd_sc_hd__nor2_1 _4959_ (.A(net1266),
    .B(_2643_),
    .Y(_2644_));
 sky130_fd_sc_hd__o21ai_0 _4960_ (.A1(net1233),
    .A2(_2644_),
    .B1(net664),
    .Y(_2645_));
 sky130_fd_sc_hd__o31ai_1 _4961_ (.A1(net664),
    .A2(net1266),
    .A3(_2642_),
    .B1(_2645_),
    .Y(_0347_));
 sky130_fd_sc_hd__and3_1 _4962_ (.A(net1270),
    .B(net664),
    .C(_2639_),
    .X(_2646_));
 sky130_fd_sc_hd__xor2_1 _4963_ (.A(net665),
    .B(_2646_),
    .X(_0839_));
 sky130_fd_sc_hd__nand2_1 _4964_ (.A(_1611_),
    .B(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__nand2_1 _4965_ (.A(_1618_),
    .B(net1266),
    .Y(_2648_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input94 (.A(net1494),
    .X(net94));
 sky130_fd_sc_hd__o21ai_0 _4967_ (.A1(net1266),
    .A2(_2646_),
    .B1(_2648_),
    .Y(_2650_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(net665),
    .B(_2650_),
    .Y(_2651_));
 sky130_fd_sc_hd__o21ai_0 _4969_ (.A1(net665),
    .A2(_2647_),
    .B1(_2651_),
    .Y(_0348_));
 sky130_fd_sc_hd__and3_1 _4970_ (.A(net664),
    .B(net665),
    .C(_2643_),
    .X(_2652_));
 sky130_fd_sc_hd__xor2_1 _4971_ (.A(net666),
    .B(_2652_),
    .X(_0835_));
 sky130_fd_sc_hd__o21ai_0 _4972_ (.A1(net1266),
    .A2(_2652_),
    .B1(_2648_),
    .Y(_2653_));
 sky130_fd_sc_hd__nor2_1 _4973_ (.A(net666),
    .B(net1266),
    .Y(_2654_));
 sky130_fd_sc_hd__a22o_1 _4974_ (.A1(net666),
    .A2(_2653_),
    .B1(_2654_),
    .B2(_2652_),
    .X(_0318_));
 sky130_fd_sc_hd__and4_1 _4975_ (.A(net1270),
    .B(net664),
    .C(net665),
    .D(net666),
    .X(_2655_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input93 (.A(net1301),
    .X(net93));
 sky130_fd_sc_hd__nand2_1 _4977_ (.A(_2639_),
    .B(_2655_),
    .Y(_2657_));
 sky130_fd_sc_hd__xnor2_1 _4978_ (.A(net667),
    .B(_2657_),
    .Y(_0831_));
 sky130_fd_sc_hd__a21oi_1 _4979_ (.A1(_2639_),
    .A2(_2655_),
    .B1(net1266),
    .Y(_2658_));
 sky130_fd_sc_hd__o21ai_0 _4980_ (.A1(net1233),
    .A2(_2658_),
    .B1(net667),
    .Y(_2659_));
 sky130_fd_sc_hd__o31ai_1 _4981_ (.A1(net667),
    .A2(net1266),
    .A3(_2657_),
    .B1(_2659_),
    .Y(_0319_));
 sky130_fd_sc_hd__nand4_1 _4982_ (.A(net667),
    .B(_2632_),
    .C(_2637_),
    .D(_2655_),
    .Y(_2660_));
 sky130_fd_sc_hd__xnor2_1 _4983_ (.A(net668),
    .B(_2660_),
    .Y(_0827_));
 sky130_fd_sc_hd__and2_0 _4984_ (.A(_1611_),
    .B(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__o21ai_0 _4985_ (.A1(net1233),
    .A2(_2661_),
    .B1(net668),
    .Y(_2662_));
 sky130_fd_sc_hd__o31ai_1 _4986_ (.A1(net668),
    .A2(net1266),
    .A3(_2660_),
    .B1(_2662_),
    .Y(_0320_));
 sky130_fd_sc_hd__nand4_1 _4987_ (.A(net667),
    .B(net668),
    .C(_2639_),
    .D(_2655_),
    .Y(_2663_));
 sky130_fd_sc_hd__xnor2_1 _4988_ (.A(net669),
    .B(_2663_),
    .Y(_0823_));
 sky130_fd_sc_hd__a21o_1 _4989_ (.A1(_1611_),
    .A2(_2663_),
    .B1(net1233),
    .X(_2664_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(net669),
    .B(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__o31ai_1 _4991_ (.A1(net669),
    .A2(net1266),
    .A3(_2663_),
    .B1(_2665_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _4992_ (.A(net668),
    .B(net669),
    .Y(_2666_));
 sky130_fd_sc_hd__nor2_1 _4993_ (.A(_2660_),
    .B(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__xor2_1 _4994_ (.A(net670),
    .B(_2667_),
    .X(_0819_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_1611_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__o21ai_0 _4996_ (.A1(net1266),
    .A2(_2667_),
    .B1(_2648_),
    .Y(_2669_));
 sky130_fd_sc_hd__nand2_1 _4997_ (.A(net670),
    .B(_2669_),
    .Y(_2670_));
 sky130_fd_sc_hd__o21ai_0 _4998_ (.A1(net670),
    .A2(_2668_),
    .B1(_2670_),
    .Y(_0322_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input92 (.A(net1345),
    .X(net92));
 sky130_fd_sc_hd__nand2_1 _5000_ (.A(net667),
    .B(_2655_),
    .Y(_2672_));
 sky130_fd_sc_hd__nand3_1 _5001_ (.A(net668),
    .B(net669),
    .C(net670),
    .Y(_2673_));
 sky130_fd_sc_hd__nor3_2 _5002_ (.A(net1241),
    .B(_2672_),
    .C(_2673_),
    .Y(_2674_));
 sky130_fd_sc_hd__xor2_1 _5003_ (.A(net671),
    .B(_2674_),
    .X(_0815_));
 sky130_fd_sc_hd__nand2_1 _5004_ (.A(_1611_),
    .B(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__o21ai_0 _5005_ (.A1(net1266),
    .A2(_2674_),
    .B1(_2648_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_1 _5006_ (.A(net671),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__o21ai_0 _5007_ (.A1(net671),
    .A2(_2675_),
    .B1(_2677_),
    .Y(_0323_));
 sky130_fd_sc_hd__nand3_1 _5008_ (.A(net670),
    .B(net671),
    .C(_2667_),
    .Y(_2678_));
 sky130_fd_sc_hd__xnor2_1 _5009_ (.A(net673),
    .B(_2678_),
    .Y(_0907_));
 sky130_fd_sc_hd__a31oi_1 _5010_ (.A1(net670),
    .A2(net671),
    .A3(_2667_),
    .B1(net1266),
    .Y(_2679_));
 sky130_fd_sc_hd__o21ai_0 _5011_ (.A1(net1233),
    .A2(_2679_),
    .B1(net673),
    .Y(_2680_));
 sky130_fd_sc_hd__o31ai_1 _5012_ (.A1(net673),
    .A2(net1266),
    .A3(_2678_),
    .B1(_2680_),
    .Y(_0324_));
 sky130_fd_sc_hd__nand3_1 _5013_ (.A(net671),
    .B(net673),
    .C(_2674_),
    .Y(_2681_));
 sky130_fd_sc_hd__xnor2_1 _5014_ (.A(net674),
    .B(_2681_),
    .Y(_0903_));
 sky130_fd_sc_hd__a31oi_1 _5015_ (.A1(net671),
    .A2(net673),
    .A3(_2674_),
    .B1(net1266),
    .Y(_2682_));
 sky130_fd_sc_hd__o21ai_0 _5016_ (.A1(net1233),
    .A2(_2682_),
    .B1(net674),
    .Y(_2683_));
 sky130_fd_sc_hd__o31ai_1 _5017_ (.A1(net674),
    .A2(net1266),
    .A3(_2681_),
    .B1(_2683_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand3_1 _5018_ (.A(net671),
    .B(net673),
    .C(net674),
    .Y(_2684_));
 sky130_fd_sc_hd__nor3_1 _5019_ (.A(_2660_),
    .B(_2673_),
    .C(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__xor2_1 _5020_ (.A(net675),
    .B(_2685_),
    .X(_0899_));
 sky130_fd_sc_hd__nand2_1 _5021_ (.A(_1611_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__o21ai_0 _5022_ (.A1(net1266),
    .A2(_2685_),
    .B1(_2648_),
    .Y(_2687_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(net675),
    .B(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__o21ai_0 _5024_ (.A1(net675),
    .A2(_2686_),
    .B1(_2688_),
    .Y(_0326_));
 sky130_fd_sc_hd__and4_1 _5025_ (.A(net671),
    .B(net673),
    .C(net674),
    .D(net675),
    .X(_2689_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input91 (.A(net1336),
    .X(net91));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_2674_),
    .B(_2689_),
    .Y(_2691_));
 sky130_fd_sc_hd__xnor2_1 _5028_ (.A(net676),
    .B(_2691_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_1 _5029_ (.A(_1611_),
    .B(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__a31oi_1 _5030_ (.A1(_1611_),
    .A2(_2674_),
    .A3(_2689_),
    .B1(net676),
    .Y(_2693_));
 sky130_fd_sc_hd__a31oi_1 _5031_ (.A1(net676),
    .A2(_2648_),
    .A3(_2692_),
    .B1(_2693_),
    .Y(_0327_));
 sky130_fd_sc_hd__and2_1 _5032_ (.A(net676),
    .B(_2689_),
    .X(_2694_));
 sky130_fd_sc_hd__nor3b_1 _5033_ (.A(_2660_),
    .B(_2673_),
    .C_N(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__xor2_1 _5034_ (.A(net677),
    .B(_2695_),
    .X(_0891_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_1611_),
    .B(_2695_),
    .Y(_2696_));
 sky130_fd_sc_hd__o21ai_0 _5036_ (.A1(net1266),
    .A2(_2695_),
    .B1(_2648_),
    .Y(_2697_));
 sky130_fd_sc_hd__nand2_1 _5037_ (.A(net677),
    .B(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__o21ai_0 _5038_ (.A1(net677),
    .A2(_2696_),
    .B1(_2698_),
    .Y(_0329_));
 sky130_fd_sc_hd__and3_1 _5039_ (.A(net677),
    .B(_2674_),
    .C(_2694_),
    .X(_2699_));
 sky130_fd_sc_hd__xor2_1 _5040_ (.A(net678),
    .B(_2699_),
    .X(_0887_));
 sky130_fd_sc_hd__o21ai_0 _5041_ (.A1(net1266),
    .A2(_2699_),
    .B1(_2648_),
    .Y(_2700_));
 sky130_fd_sc_hd__nor2_1 _5042_ (.A(net678),
    .B(net1266),
    .Y(_2701_));
 sky130_fd_sc_hd__a22o_1 _5043_ (.A1(net678),
    .A2(_2700_),
    .B1(_2701_),
    .B2(_2699_),
    .X(_0330_));
 sky130_fd_sc_hd__nor2_1 _5044_ (.A(_2660_),
    .B(_2673_),
    .Y(_2702_));
 sky130_fd_sc_hd__and3_1 _5045_ (.A(net676),
    .B(net677),
    .C(net678),
    .X(_2703_));
 sky130_fd_sc_hd__nand3_1 _5046_ (.A(_2702_),
    .B(_2689_),
    .C(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__xnor2_1 _5047_ (.A(net679),
    .B(_2704_),
    .Y(_0883_));
 sky130_fd_sc_hd__a31oi_1 _5048_ (.A1(_2702_),
    .A2(_2689_),
    .A3(_2703_),
    .B1(net1266),
    .Y(_2705_));
 sky130_fd_sc_hd__o21ai_0 _5049_ (.A1(net1233),
    .A2(_2705_),
    .B1(net679),
    .Y(_2706_));
 sky130_fd_sc_hd__o31ai_1 _5050_ (.A1(net679),
    .A2(net1266),
    .A3(_2704_),
    .B1(_2706_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_1 _5051_ (.A(net680),
    .Y(_2707_));
 sky130_fd_sc_hd__and3_1 _5052_ (.A(net668),
    .B(net669),
    .C(net670),
    .X(_2708_));
 sky130_fd_sc_hd__nand4_1 _5053_ (.A(net679),
    .B(_2708_),
    .C(_2689_),
    .D(_2703_),
    .Y(_2709_));
 sky130_fd_sc_hd__nor3_1 _5054_ (.A(net1241),
    .B(_2672_),
    .C(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__xnor2_1 _5055_ (.A(_2707_),
    .B(_2710_),
    .Y(_0879_));
 sky130_fd_sc_hd__nand2_1 _5056_ (.A(_1611_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__o21ai_0 _5057_ (.A1(net1266),
    .A2(_2710_),
    .B1(_2648_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand2_1 _5058_ (.A(net680),
    .B(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__o21ai_0 _5059_ (.A1(net680),
    .A2(_2711_),
    .B1(_2713_),
    .Y(_0332_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input90 (.A(net1298),
    .X(net90));
 sky130_fd_sc_hd__nor3_2 _5061_ (.A(_2707_),
    .B(_2660_),
    .C(_2709_),
    .Y(_2715_));
 sky130_fd_sc_hd__xor2_1 _5062_ (.A(net681),
    .B(_2715_),
    .X(_0875_));
 sky130_fd_sc_hd__nand2_1 _5063_ (.A(_1611_),
    .B(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__o21ai_0 _5064_ (.A1(net1266),
    .A2(_2715_),
    .B1(_2648_),
    .Y(_2717_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(net681),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__o21ai_0 _5066_ (.A1(net681),
    .A2(_2716_),
    .B1(_2718_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand3_1 _5067_ (.A(net680),
    .B(net681),
    .C(_2710_),
    .Y(_2719_));
 sky130_fd_sc_hd__xnor2_1 _5068_ (.A(net682),
    .B(_2719_),
    .Y(_0871_));
 sky130_fd_sc_hd__a31oi_1 _5069_ (.A1(net680),
    .A2(net681),
    .A3(_2710_),
    .B1(net1266),
    .Y(_2720_));
 sky130_fd_sc_hd__o21ai_0 _5070_ (.A1(net1233),
    .A2(_2720_),
    .B1(net682),
    .Y(_2721_));
 sky130_fd_sc_hd__o31ai_1 _5071_ (.A1(net682),
    .A2(net1266),
    .A3(_2719_),
    .B1(_2721_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand3_1 _5072_ (.A(net681),
    .B(net682),
    .C(_2715_),
    .Y(_2722_));
 sky130_fd_sc_hd__xnor2_1 _5073_ (.A(net684),
    .B(_2722_),
    .Y(_0867_));
 sky130_fd_sc_hd__a31oi_1 _5074_ (.A1(net681),
    .A2(net682),
    .A3(_2715_),
    .B1(net1266),
    .Y(_2723_));
 sky130_fd_sc_hd__o21ai_0 _5075_ (.A1(net1233),
    .A2(_2723_),
    .B1(net684),
    .Y(_2724_));
 sky130_fd_sc_hd__o31ai_1 _5076_ (.A1(net684),
    .A2(net1266),
    .A3(_2722_),
    .B1(_2724_),
    .Y(_0335_));
 sky130_fd_sc_hd__and3_1 _5077_ (.A(net681),
    .B(net682),
    .C(net684),
    .X(_2725_));
 sky130_fd_sc_hd__nand2_1 _5078_ (.A(net680),
    .B(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__or4_4 _5079_ (.A(net1241),
    .B(_2672_),
    .C(_2709_),
    .D(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__xnor2_1 _5080_ (.A(net685),
    .B(_2727_),
    .Y(_0863_));
 sky130_fd_sc_hd__nand2_1 _5081_ (.A(_1611_),
    .B(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__nor2_1 _5082_ (.A(net1266),
    .B(_2727_),
    .Y(_2729_));
 sky130_fd_sc_hd__nor2_1 _5083_ (.A(net685),
    .B(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__a31oi_1 _5084_ (.A1(net685),
    .A2(_2648_),
    .A3(_2728_),
    .B1(_2730_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand3_1 _5085_ (.A(net685),
    .B(_2715_),
    .C(_2725_),
    .Y(_2731_));
 sky130_fd_sc_hd__xnor2_1 _5086_ (.A(net686),
    .B(_2731_),
    .Y(_0859_));
 sky130_fd_sc_hd__o211ai_1 _5087_ (.A1(net1266),
    .A2(_2731_),
    .B1(net686),
    .C1(_1618_),
    .Y(_2732_));
 sky130_fd_sc_hd__o31ai_1 _5088_ (.A1(net686),
    .A2(net1266),
    .A3(_2731_),
    .B1(_2732_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _5089_ (.A(net685),
    .B(net686),
    .Y(_2733_));
 sky130_fd_sc_hd__nor2_2 _5090_ (.A(_2727_),
    .B(_2733_),
    .Y(_2734_));
 sky130_fd_sc_hd__xor2_1 _5091_ (.A(net687),
    .B(_2734_),
    .X(_0855_));
 sky130_fd_sc_hd__o21ai_0 _5092_ (.A1(net1266),
    .A2(_2734_),
    .B1(_2648_),
    .Y(_2735_));
 sky130_fd_sc_hd__nor2_1 _5093_ (.A(net687),
    .B(net1266),
    .Y(_2736_));
 sky130_fd_sc_hd__a22o_1 _5094_ (.A1(net687),
    .A2(_2735_),
    .B1(_2736_),
    .B2(_2734_),
    .X(_0338_));
 sky130_fd_sc_hd__and4_1 _5095_ (.A(net685),
    .B(net686),
    .C(net687),
    .D(_2725_),
    .X(_2737_));
 sky130_fd_sc_hd__nand2_1 _5096_ (.A(_2715_),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__xnor2_1 _5097_ (.A(net688),
    .B(_2738_),
    .Y(_0851_));
 sky130_fd_sc_hd__a21oi_1 _5098_ (.A1(_2715_),
    .A2(_2737_),
    .B1(net1266),
    .Y(_2739_));
 sky130_fd_sc_hd__o21ai_0 _5099_ (.A1(net1233),
    .A2(_2739_),
    .B1(net688),
    .Y(_2740_));
 sky130_fd_sc_hd__o31ai_1 _5100_ (.A1(net688),
    .A2(net1266),
    .A3(_2738_),
    .B1(_2740_),
    .Y(_0340_));
 sky130_fd_sc_hd__nand4_1 _5101_ (.A(net680),
    .B(net688),
    .C(_2710_),
    .D(_2737_),
    .Y(_2741_));
 sky130_fd_sc_hd__xnor2_1 _5102_ (.A(net689),
    .B(_2741_),
    .Y(_0847_));
 sky130_fd_sc_hd__o211ai_1 _5103_ (.A1(net1266),
    .A2(_2741_),
    .B1(net689),
    .C1(_1618_),
    .Y(_2742_));
 sky130_fd_sc_hd__o31ai_1 _5104_ (.A1(net689),
    .A2(net1266),
    .A3(_2741_),
    .B1(_2742_),
    .Y(_0341_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input89 (.A(net1297),
    .X(net89));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input88 (.A(net1458),
    .X(net88));
 sky130_fd_sc_hd__nor2_2 _5107_ (.A(_1733_),
    .B(net1264),
    .Y(_2745_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input87 (.A(net1609),
    .X(net87));
 sky130_fd_sc_hd__nand2_1 _5109_ (.A(net620),
    .B(net1232),
    .Y(_2747_));
 sky130_fd_sc_hd__o21ai_0 _5110_ (.A1(net620),
    .A2(net1265),
    .B1(_2747_),
    .Y(_0285_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input86 (.A(net1549),
    .X(net86));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(net621),
    .B(net1265),
    .Y(_2749_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input85 (.A(net1500),
    .X(net85));
 sky130_fd_sc_hd__nand2_1 _5114_ (.A(_0402_),
    .B(net1264),
    .Y(_2751_));
 sky130_fd_sc_hd__o21ai_0 _5115_ (.A1(_1733_),
    .A2(_2749_),
    .B1(_2751_),
    .Y(_0296_));
 sky130_fd_sc_hd__xor2_1 _5116_ (.A(net622),
    .B(_0401_),
    .X(_0545_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input84 (.A(net1616),
    .X(net84));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_0401_),
    .B(net1264),
    .Y(_2753_));
 sky130_fd_sc_hd__nor2_1 _5119_ (.A(_0401_),
    .B(net1265),
    .Y(_2754_));
 sky130_fd_sc_hd__o21ai_0 _5120_ (.A1(net1232),
    .A2(_2754_),
    .B1(net622),
    .Y(_2755_));
 sky130_fd_sc_hd__o21ai_0 _5121_ (.A1(net622),
    .A2(_2753_),
    .B1(_2755_),
    .Y(_0307_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input83 (.A(net1479),
    .X(net83));
 sky130_fd_sc_hd__nand3_1 _5123_ (.A(net620),
    .B(net621),
    .C(net622),
    .Y(_2757_));
 sky130_fd_sc_hd__xnor2_1 _5124_ (.A(net623),
    .B(_2757_),
    .Y(_0541_));
 sky130_fd_sc_hd__and3_1 _5125_ (.A(net620),
    .B(net621),
    .C(net622),
    .X(_2758_));
 sky130_fd_sc_hd__nor2_1 _5126_ (.A(net1265),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__o21ai_0 _5127_ (.A1(net1232),
    .A2(_2759_),
    .B1(net623),
    .Y(_2760_));
 sky130_fd_sc_hd__o31ai_1 _5128_ (.A1(net623),
    .A2(net1265),
    .A3(_2757_),
    .B1(_2760_),
    .Y(_0310_));
 sky130_fd_sc_hd__nand3_1 _5129_ (.A(net622),
    .B(_0401_),
    .C(net623),
    .Y(_2761_));
 sky130_fd_sc_hd__xnor2_1 _5130_ (.A(net624),
    .B(_2761_),
    .Y(_0561_));
 sky130_fd_sc_hd__a22o_1 _5131_ (.A1(net624),
    .A2(net1232),
    .B1(_0561_),
    .B2(net1264),
    .X(_0311_));
 sky130_fd_sc_hd__nand3_1 _5132_ (.A(net623),
    .B(net624),
    .C(_2758_),
    .Y(_2762_));
 sky130_fd_sc_hd__xnor2_1 _5133_ (.A(net625),
    .B(_2762_),
    .Y(_0557_));
 sky130_fd_sc_hd__a22o_1 _5134_ (.A1(net625),
    .A2(net1232),
    .B1(_0557_),
    .B2(net1264),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _5135_ (.A(net622),
    .B(_0401_),
    .Y(_2763_));
 sky130_fd_sc_hd__nand3_1 _5136_ (.A(net623),
    .B(net624),
    .C(net625),
    .Y(_2764_));
 sky130_fd_sc_hd__nor2_1 _5137_ (.A(_2763_),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__xor2_1 _5138_ (.A(net626),
    .B(_2765_),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _5139_ (.A1(net626),
    .A2(net1232),
    .B1(_0553_),
    .B2(net1264),
    .X(_0313_));
 sky130_fd_sc_hd__inv_1 _5140_ (.A(net627),
    .Y(_2766_));
 sky130_fd_sc_hd__nand4_1 _5141_ (.A(net623),
    .B(net624),
    .C(net625),
    .D(net626),
    .Y(_2767_));
 sky130_fd_sc_hd__nor2_1 _5142_ (.A(_2757_),
    .B(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__xnor2_1 _5143_ (.A(_2766_),
    .B(_2768_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(net1264),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__nor2_1 _5145_ (.A(net1265),
    .B(_2768_),
    .Y(_2770_));
 sky130_fd_sc_hd__o21ai_0 _5146_ (.A1(net1232),
    .A2(_2770_),
    .B1(net627),
    .Y(_2771_));
 sky130_fd_sc_hd__o21ai_0 _5147_ (.A1(net627),
    .A2(_2769_),
    .B1(_2771_),
    .Y(_0314_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input82 (.A(net1402),
    .X(net82));
 sky130_fd_sc_hd__or3_1 _5149_ (.A(_2766_),
    .B(_2763_),
    .C(_2767_),
    .X(_2773_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input81 (.A(net1620),
    .X(net81));
 sky130_fd_sc_hd__xnor2_1 _5151_ (.A(net629),
    .B(_2773_),
    .Y(_0593_));
 sky130_fd_sc_hd__and2_1 _5152_ (.A(net1264),
    .B(_2773_),
    .X(_2775_));
 sky130_fd_sc_hd__o21ai_0 _5153_ (.A1(net1232),
    .A2(_2775_),
    .B1(net629),
    .Y(_2776_));
 sky130_fd_sc_hd__o31ai_1 _5154_ (.A1(net629),
    .A2(net1265),
    .A3(_2773_),
    .B1(_2776_),
    .Y(_0315_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input80 (.A(net1433),
    .X(net80));
 sky130_fd_sc_hd__and4_1 _5156_ (.A(net623),
    .B(net624),
    .C(net625),
    .D(net626),
    .X(_2778_));
 sky130_fd_sc_hd__nand4_1 _5157_ (.A(net627),
    .B(net629),
    .C(_2758_),
    .D(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__xnor2_1 _5158_ (.A(net630),
    .B(_2779_),
    .Y(_0589_));
 sky130_fd_sc_hd__and2_1 _5159_ (.A(net1264),
    .B(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__o21ai_0 _5160_ (.A1(net1232),
    .A2(_2780_),
    .B1(net630),
    .Y(_2781_));
 sky130_fd_sc_hd__o31ai_1 _5161_ (.A1(net630),
    .A2(net1265),
    .A3(_2779_),
    .B1(_2781_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _5162_ (.A(net629),
    .B(net630),
    .Y(_2782_));
 sky130_fd_sc_hd__nor4_1 _5163_ (.A(_2766_),
    .B(_2763_),
    .C(_2767_),
    .D(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__xor2_1 _5164_ (.A(net631),
    .B(net1231),
    .X(_0585_));
 sky130_fd_sc_hd__nand2_1 _5165_ (.A(net1264),
    .B(net1231),
    .Y(_2784_));
 sky130_fd_sc_hd__nor2_1 _5166_ (.A(net1265),
    .B(net1231),
    .Y(_2785_));
 sky130_fd_sc_hd__o21ai_0 _5167_ (.A1(net1232),
    .A2(_2785_),
    .B1(net631),
    .Y(_2786_));
 sky130_fd_sc_hd__o21ai_0 _5168_ (.A1(net631),
    .A2(_2784_),
    .B1(_2786_),
    .Y(_0286_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input79 (.A(net1614),
    .X(net79));
 sky130_fd_sc_hd__nand2_1 _5170_ (.A(net630),
    .B(net631),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2_1 _5171_ (.A(_2779_),
    .B(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__xor2_1 _5172_ (.A(net632),
    .B(_2789_),
    .X(_0581_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(net1264),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input78 (.A(net1490),
    .X(net78));
 sky130_fd_sc_hd__nand2_1 _5175_ (.A(_1748_),
    .B(net1265),
    .Y(_2792_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input77 (.A(net1587),
    .X(net77));
 sky130_fd_sc_hd__o21ai_0 _5177_ (.A1(net1265),
    .A2(_2789_),
    .B1(_2792_),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(net632),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__o21ai_0 _5179_ (.A1(net632),
    .A2(_2790_),
    .B1(_2795_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand3_1 _5180_ (.A(net631),
    .B(net632),
    .C(net1231),
    .Y(_2796_));
 sky130_fd_sc_hd__xnor2_1 _5181_ (.A(net633),
    .B(_2796_),
    .Y(_0577_));
 sky130_fd_sc_hd__a31oi_1 _5182_ (.A1(net631),
    .A2(net632),
    .A3(net1231),
    .B1(net1265),
    .Y(_2797_));
 sky130_fd_sc_hd__o21ai_0 _5183_ (.A1(net1232),
    .A2(_2797_),
    .B1(net633),
    .Y(_2798_));
 sky130_fd_sc_hd__o31ai_1 _5184_ (.A1(net633),
    .A2(net1265),
    .A3(_2796_),
    .B1(_2798_),
    .Y(_0288_));
 sky130_fd_sc_hd__and3_1 _5185_ (.A(net632),
    .B(net633),
    .C(_2789_),
    .X(_2799_));
 sky130_fd_sc_hd__xor2_1 _5186_ (.A(net634),
    .B(_2799_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _5187_ (.A(net1264),
    .B(_2799_),
    .Y(_2800_));
 sky130_fd_sc_hd__a31oi_1 _5188_ (.A1(net632),
    .A2(net633),
    .A3(_2789_),
    .B1(net1265),
    .Y(_2801_));
 sky130_fd_sc_hd__o21ai_0 _5189_ (.A1(net1232),
    .A2(_2801_),
    .B1(net634),
    .Y(_2802_));
 sky130_fd_sc_hd__o21ai_0 _5190_ (.A1(net634),
    .A2(_2800_),
    .B1(_2802_),
    .Y(_0289_));
 sky130_fd_sc_hd__and4_1 _5191_ (.A(net631),
    .B(net632),
    .C(net633),
    .D(net634),
    .X(_2803_));
 sky130_fd_sc_hd__and2_1 _5192_ (.A(net1231),
    .B(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__xor2_1 _5193_ (.A(net635),
    .B(_2804_),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_1 _5194_ (.A(net1264),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__o21ai_0 _5195_ (.A1(net1265),
    .A2(_2804_),
    .B1(_2792_),
    .Y(_2806_));
 sky130_fd_sc_hd__nand2_1 _5196_ (.A(net635),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__o21ai_0 _5197_ (.A1(net635),
    .A2(_2805_),
    .B1(_2807_),
    .Y(_0290_));
 sky130_fd_sc_hd__nand3_1 _5198_ (.A(net627),
    .B(_2758_),
    .C(_2778_),
    .Y(_2808_));
 sky130_fd_sc_hd__nand4_2 _5199_ (.A(net629),
    .B(net630),
    .C(net635),
    .D(_2803_),
    .Y(_2809_));
 sky130_fd_sc_hd__nor2_1 _5200_ (.A(_2808_),
    .B(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__xor2_1 _5201_ (.A(net636),
    .B(_2810_),
    .X(_0565_));
 sky130_fd_sc_hd__nand2_1 _5202_ (.A(net1264),
    .B(_2810_),
    .Y(_2811_));
 sky130_fd_sc_hd__o21ai_0 _5203_ (.A1(net1265),
    .A2(_2810_),
    .B1(_2792_),
    .Y(_2812_));
 sky130_fd_sc_hd__nand2_1 _5204_ (.A(net636),
    .B(_2812_),
    .Y(_2813_));
 sky130_fd_sc_hd__o21ai_0 _5205_ (.A1(net636),
    .A2(_2811_),
    .B1(_2813_),
    .Y(_0291_));
 sky130_fd_sc_hd__nand4_1 _5206_ (.A(net635),
    .B(net636),
    .C(net1231),
    .D(_2803_),
    .Y(_2814_));
 sky130_fd_sc_hd__xnor2_1 _5207_ (.A(net637),
    .B(_2814_),
    .Y(_0657_));
 sky130_fd_sc_hd__a21o_1 _5208_ (.A1(net1264),
    .A2(_2814_),
    .B1(net1232),
    .X(_2815_));
 sky130_fd_sc_hd__nand2_1 _5209_ (.A(net637),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__o31ai_1 _5210_ (.A1(net637),
    .A2(net1265),
    .A3(_2814_),
    .B1(_2816_),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _5211_ (.A(net636),
    .B(net637),
    .Y(_2817_));
 sky130_fd_sc_hd__nor3_1 _5212_ (.A(_2808_),
    .B(_2809_),
    .C(_2817_),
    .Y(_2818_));
 sky130_fd_sc_hd__xor2_1 _5213_ (.A(net638),
    .B(_2818_),
    .X(_0653_));
 sky130_fd_sc_hd__o21ai_0 _5214_ (.A1(net1265),
    .A2(_2818_),
    .B1(_2792_),
    .Y(_2819_));
 sky130_fd_sc_hd__nand2_1 _5215_ (.A(net638),
    .B(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__nand3b_1 _5216_ (.A_N(net638),
    .B(net1264),
    .C(_2818_),
    .Y(_2821_));
 sky130_fd_sc_hd__nand2_1 _5217_ (.A(_2820_),
    .B(_2821_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand3_1 _5218_ (.A(net636),
    .B(net637),
    .C(net638),
    .Y(_2822_));
 sky130_fd_sc_hd__nor3_1 _5219_ (.A(_2773_),
    .B(_2809_),
    .C(_2822_),
    .Y(_2823_));
 sky130_fd_sc_hd__xor2_1 _5220_ (.A(net640),
    .B(_2823_),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_1 _5221_ (.A(net1264),
    .B(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__o21ai_0 _5222_ (.A1(net1265),
    .A2(_2823_),
    .B1(_2792_),
    .Y(_2825_));
 sky130_fd_sc_hd__nand2_1 _5223_ (.A(net640),
    .B(_2825_),
    .Y(_2826_));
 sky130_fd_sc_hd__o21ai_0 _5224_ (.A1(net640),
    .A2(_2824_),
    .B1(_2826_),
    .Y(_0294_));
 sky130_fd_sc_hd__and4_1 _5225_ (.A(net636),
    .B(net637),
    .C(net638),
    .D(net640),
    .X(_2827_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input76 (.A(net1393),
    .X(net76));
 sky130_fd_sc_hd__nand2_1 _5227_ (.A(_2810_),
    .B(_2827_),
    .Y(_2829_));
 sky130_fd_sc_hd__xnor2_1 _5228_ (.A(net641),
    .B(_2829_),
    .Y(_0645_));
 sky130_fd_sc_hd__a21oi_1 _5229_ (.A1(_2810_),
    .A2(_2827_),
    .B1(net1265),
    .Y(_2830_));
 sky130_fd_sc_hd__o21ai_0 _5230_ (.A1(net1232),
    .A2(_2830_),
    .B1(net641),
    .Y(_2831_));
 sky130_fd_sc_hd__o31ai_1 _5231_ (.A1(net641),
    .A2(net1265),
    .A3(_2829_),
    .B1(_2831_),
    .Y(_0295_));
 sky130_fd_sc_hd__nor2_1 _5232_ (.A(_2773_),
    .B(_2809_),
    .Y(_2832_));
 sky130_fd_sc_hd__nand3_1 _5233_ (.A(net641),
    .B(_2832_),
    .C(_2827_),
    .Y(_2833_));
 sky130_fd_sc_hd__xnor2_1 _5234_ (.A(net642),
    .B(_2833_),
    .Y(_0641_));
 sky130_fd_sc_hd__a31oi_1 _5235_ (.A1(net641),
    .A2(_2832_),
    .A3(_2827_),
    .B1(net1265),
    .Y(_2834_));
 sky130_fd_sc_hd__o21ai_0 _5236_ (.A1(net1232),
    .A2(_2834_),
    .B1(net642),
    .Y(_2835_));
 sky130_fd_sc_hd__o31ai_1 _5237_ (.A1(net642),
    .A2(net1265),
    .A3(_2833_),
    .B1(_2835_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_1 _5238_ (.A(net643),
    .Y(_2836_));
 sky130_fd_sc_hd__nand3_1 _5239_ (.A(net641),
    .B(net642),
    .C(_2827_),
    .Y(_2837_));
 sky130_fd_sc_hd__nor3_1 _5240_ (.A(_2808_),
    .B(_2809_),
    .C(_2837_),
    .Y(_2838_));
 sky130_fd_sc_hd__xnor2_1 _5241_ (.A(_2836_),
    .B(_2838_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(net1264),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__o21ai_0 _5243_ (.A1(net1265),
    .A2(_2838_),
    .B1(_2792_),
    .Y(_2840_));
 sky130_fd_sc_hd__nand2_1 _5244_ (.A(net643),
    .B(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__o21ai_0 _5245_ (.A1(net643),
    .A2(_2839_),
    .B1(_2841_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor4_1 _5246_ (.A(_2836_),
    .B(_2773_),
    .C(_2809_),
    .D(_2837_),
    .Y(_2842_));
 sky130_fd_sc_hd__xor2_1 _5247_ (.A(net644),
    .B(_2842_),
    .X(_0633_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(net1264),
    .B(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__o21ai_0 _5249_ (.A1(net1265),
    .A2(_2842_),
    .B1(_2792_),
    .Y(_2844_));
 sky130_fd_sc_hd__nand2_1 _5250_ (.A(net644),
    .B(_2844_),
    .Y(_2845_));
 sky130_fd_sc_hd__o21ai_0 _5251_ (.A1(net644),
    .A2(_2843_),
    .B1(_2845_),
    .Y(_0299_));
 sky130_fd_sc_hd__and4_1 _5252_ (.A(net641),
    .B(net642),
    .C(net643),
    .D(net644),
    .X(_2846_));
 sky130_fd_sc_hd__nand2_1 _5253_ (.A(_2827_),
    .B(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nor3_1 _5254_ (.A(_2808_),
    .B(_2809_),
    .C(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__xor2_1 _5255_ (.A(net645),
    .B(_2848_),
    .X(_0628_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(net1264),
    .B(_2848_),
    .Y(_2849_));
 sky130_fd_sc_hd__o21ai_0 _5257_ (.A1(net1265),
    .A2(_2848_),
    .B1(_2792_),
    .Y(_2850_));
 sky130_fd_sc_hd__nand2_1 _5258_ (.A(net645),
    .B(_2850_),
    .Y(_2851_));
 sky130_fd_sc_hd__o21ai_0 _5259_ (.A1(net645),
    .A2(_2849_),
    .B1(_2851_),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_1 _5260_ (.A(net646),
    .Y(_2852_));
 sky130_fd_sc_hd__nand3_1 _5261_ (.A(net645),
    .B(_2827_),
    .C(_2846_),
    .Y(_2853_));
 sky130_fd_sc_hd__nor3_1 _5262_ (.A(_2773_),
    .B(_2809_),
    .C(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__xnor2_1 _5263_ (.A(_2852_),
    .B(_2854_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _5264_ (.A(net1264),
    .B(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__o21ai_0 _5265_ (.A1(net1265),
    .A2(_2854_),
    .B1(_2792_),
    .Y(_2856_));
 sky130_fd_sc_hd__nand2_1 _5266_ (.A(net646),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__o21ai_0 _5267_ (.A1(net646),
    .A2(_2855_),
    .B1(_2857_),
    .Y(_0301_));
 sky130_fd_sc_hd__nor4_1 _5268_ (.A(_2852_),
    .B(_2808_),
    .C(_2809_),
    .D(_2853_),
    .Y(_2858_));
 sky130_fd_sc_hd__xor2_1 _5269_ (.A(net647),
    .B(_2858_),
    .X(_0621_));
 sky130_fd_sc_hd__nand2_1 _5270_ (.A(net1264),
    .B(_2858_),
    .Y(_2859_));
 sky130_fd_sc_hd__o21ai_0 _5271_ (.A1(net1265),
    .A2(_2858_),
    .B1(_2792_),
    .Y(_2860_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(net647),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__o21ai_0 _5273_ (.A1(net647),
    .A2(_2859_),
    .B1(_2861_),
    .Y(_0302_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input75 (.A(net1450),
    .X(net75));
 sky130_fd_sc_hd__and2_1 _5275_ (.A(net646),
    .B(net647),
    .X(_2863_));
 sky130_fd_sc_hd__nand4_1 _5276_ (.A(net645),
    .B(_2827_),
    .C(_2846_),
    .D(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__nor3_2 _5277_ (.A(_2773_),
    .B(_2809_),
    .C(_2864_),
    .Y(_2865_));
 sky130_fd_sc_hd__xor2_1 _5278_ (.A(net648),
    .B(_2865_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(net1264),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__o21ai_0 _5280_ (.A1(net1265),
    .A2(_2865_),
    .B1(_2792_),
    .Y(_2867_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(net648),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__o21ai_0 _5282_ (.A1(net648),
    .A2(_2866_),
    .B1(_2868_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(net635),
    .B(_2803_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand3_1 _5284_ (.A(net629),
    .B(net630),
    .C(net648),
    .Y(_2870_));
 sky130_fd_sc_hd__or3_1 _5285_ (.A(_2808_),
    .B(_2869_),
    .C(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__nor2_1 _5286_ (.A(_2864_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__xor2_1 _5287_ (.A(net649),
    .B(_2872_),
    .X(_0613_));
 sky130_fd_sc_hd__nor2b_1 _5288_ (.A(_2853_),
    .B_N(_2863_),
    .Y(_2873_));
 sky130_fd_sc_hd__nand3_1 _5289_ (.A(net648),
    .B(_2810_),
    .C(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__nand2_1 _5290_ (.A(net1264),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__a21oi_1 _5291_ (.A1(net1264),
    .A2(_2872_),
    .B1(net649),
    .Y(_2876_));
 sky130_fd_sc_hd__a31oi_1 _5292_ (.A1(net649),
    .A2(_2792_),
    .A3(_2875_),
    .B1(_2876_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand3_1 _5293_ (.A(net648),
    .B(net649),
    .C(_2865_),
    .Y(_2877_));
 sky130_fd_sc_hd__xnor2_1 _5294_ (.A(net651),
    .B(_2877_),
    .Y(_0609_));
 sky130_fd_sc_hd__o211ai_1 _5295_ (.A1(net1265),
    .A2(_2877_),
    .B1(net651),
    .C1(_1748_),
    .Y(_2878_));
 sky130_fd_sc_hd__o31ai_1 _5296_ (.A1(net651),
    .A2(net1265),
    .A3(_2877_),
    .B1(_2878_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _5297_ (.A(net649),
    .B(net651),
    .Y(_2879_));
 sky130_fd_sc_hd__nor2_1 _5298_ (.A(_2874_),
    .B(_2879_),
    .Y(_2880_));
 sky130_fd_sc_hd__xor2_1 _5299_ (.A(net652),
    .B(_2880_),
    .X(_0605_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(net652),
    .B(net1264),
    .Y(_2881_));
 sky130_fd_sc_hd__or4_1 _5301_ (.A(net652),
    .B(net1265),
    .C(_2874_),
    .D(_2879_),
    .X(_2882_));
 sky130_fd_sc_hd__nand2_1 _5302_ (.A(net652),
    .B(net1232),
    .Y(_2883_));
 sky130_fd_sc_hd__o211ai_1 _5303_ (.A1(_2880_),
    .A2(_2881_),
    .B1(_2882_),
    .C1(_2883_),
    .Y(_0306_));
 sky130_fd_sc_hd__and3_1 _5304_ (.A(net649),
    .B(net651),
    .C(net652),
    .X(_2884_));
 sky130_fd_sc_hd__nand3_1 _5305_ (.A(net648),
    .B(_2865_),
    .C(_2884_),
    .Y(_2885_));
 sky130_fd_sc_hd__xnor2_1 _5306_ (.A(net653),
    .B(_2885_),
    .Y(_0600_));
 sky130_fd_sc_hd__a31oi_1 _5307_ (.A1(net648),
    .A2(_2865_),
    .A3(_2884_),
    .B1(net1265),
    .Y(_2886_));
 sky130_fd_sc_hd__o21ai_0 _5308_ (.A1(net1232),
    .A2(_2886_),
    .B1(net653),
    .Y(_2887_));
 sky130_fd_sc_hd__o31ai_1 _5309_ (.A1(net653),
    .A2(net1265),
    .A3(_2885_),
    .B1(_2887_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand3_1 _5310_ (.A(net653),
    .B(_2863_),
    .C(_2884_),
    .Y(_2888_));
 sky130_fd_sc_hd__nor3_1 _5311_ (.A(_2853_),
    .B(_2871_),
    .C(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__xor2_1 _5312_ (.A(net654),
    .B(_2889_),
    .X(_0597_));
 sky130_fd_sc_hd__nand2_1 _5313_ (.A(net654),
    .B(net1264),
    .Y(_2890_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(net654),
    .B(net1232),
    .Y(_2891_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(net654),
    .B(net1265),
    .Y(_2892_));
 sky130_fd_sc_hd__nand2_1 _5316_ (.A(_2889_),
    .B(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__o211ai_1 _5317_ (.A1(_2889_),
    .A2(_2890_),
    .B1(_2891_),
    .C1(_2893_),
    .Y(_0309_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input74 (.A(net1401),
    .X(net74));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input73 (.A(channel_dst_addr[4]),
    .X(net73));
 sky130_fd_sc_hd__nor2_2 _5320_ (.A(_1866_),
    .B(net1263),
    .Y(_2896_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input72 (.A(net1461),
    .X(net72));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(net567),
    .B(net1230),
    .Y(_2898_));
 sky130_fd_sc_hd__o21ai_0 _5323_ (.A1(net567),
    .A2(_1869_),
    .B1(_2898_),
    .Y(_0253_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input71 (.A(net1607),
    .X(net71));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(net606),
    .B(_1869_),
    .Y(_2900_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input70 (.A(net1635),
    .X(net70));
 sky130_fd_sc_hd__nand2_1 _5327_ (.A(_0404_),
    .B(net1263),
    .Y(_2902_));
 sky130_fd_sc_hd__o21ai_0 _5328_ (.A1(_1866_),
    .A2(_2900_),
    .B1(_2902_),
    .Y(_0264_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input69 (.A(net1470),
    .X(net69));
 sky130_fd_sc_hd__xor2_1 _5330_ (.A(net617),
    .B(_0403_),
    .X(_0527_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input68 (.A(net1570),
    .X(net68));
 sky130_fd_sc_hd__nand2_1 _5332_ (.A(_0403_),
    .B(net1263),
    .Y(_2905_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input67 (.A(net1436),
    .X(net67));
 sky130_fd_sc_hd__nor2_1 _5334_ (.A(_0403_),
    .B(_1869_),
    .Y(_2907_));
 sky130_fd_sc_hd__o21ai_0 _5335_ (.A1(net1230),
    .A2(_2907_),
    .B1(net617),
    .Y(_2908_));
 sky130_fd_sc_hd__o21ai_0 _5336_ (.A1(net617),
    .A2(_2905_),
    .B1(_2908_),
    .Y(_0275_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input66 (.A(channel_dst_addr[43]),
    .X(net66));
 sky130_fd_sc_hd__nand3_2 _5338_ (.A(net567),
    .B(net606),
    .C(net617),
    .Y(_2910_));
 sky130_fd_sc_hd__xnor2_1 _5339_ (.A(net628),
    .B(_2910_),
    .Y(_0523_));
 sky130_fd_sc_hd__and3_1 _5340_ (.A(net567),
    .B(net606),
    .C(net617),
    .X(_2911_));
 sky130_fd_sc_hd__nor2_1 _5341_ (.A(_1869_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__o21ai_0 _5342_ (.A1(net1230),
    .A2(_2912_),
    .B1(net628),
    .Y(_2913_));
 sky130_fd_sc_hd__o31ai_1 _5343_ (.A1(net628),
    .A2(_1869_),
    .A3(_2910_),
    .B1(_2913_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand3_1 _5344_ (.A(net617),
    .B(_0403_),
    .C(net628),
    .Y(_2914_));
 sky130_fd_sc_hd__xnor2_1 _5345_ (.A(net639),
    .B(_2914_),
    .Y(_0519_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input65 (.A(net1366),
    .X(net65));
 sky130_fd_sc_hd__a22o_1 _5347_ (.A1(net639),
    .A2(net1230),
    .B1(_0519_),
    .B2(net1263),
    .X(_0279_));
 sky130_fd_sc_hd__nand3_1 _5348_ (.A(net628),
    .B(net639),
    .C(_2911_),
    .Y(_2916_));
 sky130_fd_sc_hd__xnor2_1 _5349_ (.A(net650),
    .B(_2916_),
    .Y(_0515_));
 sky130_fd_sc_hd__a22o_1 _5350_ (.A1(net650),
    .A2(net1230),
    .B1(_0515_),
    .B2(net1263),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(net617),
    .B(_0403_),
    .Y(_2917_));
 sky130_fd_sc_hd__nand3_1 _5352_ (.A(net628),
    .B(net639),
    .C(net650),
    .Y(_2918_));
 sky130_fd_sc_hd__nor2_1 _5353_ (.A(_2917_),
    .B(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__xor2_1 _5354_ (.A(net661),
    .B(_2919_),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _5355_ (.A1(net661),
    .A2(net1230),
    .B1(_0511_),
    .B2(net1263),
    .X(_0281_));
 sky130_fd_sc_hd__inv_1 _5356_ (.A(net672),
    .Y(_2920_));
 sky130_fd_sc_hd__nand4_2 _5357_ (.A(net628),
    .B(net639),
    .C(net650),
    .D(net661),
    .Y(_2921_));
 sky130_fd_sc_hd__nor2_1 _5358_ (.A(_2910_),
    .B(_2921_),
    .Y(_2922_));
 sky130_fd_sc_hd__xnor2_1 _5359_ (.A(_2920_),
    .B(_2922_),
    .Y(_0506_));
 sky130_fd_sc_hd__nand2_1 _5360_ (.A(net1263),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input64 (.A(net1636),
    .X(net64));
 sky130_fd_sc_hd__nor2_1 _5362_ (.A(_1869_),
    .B(_2922_),
    .Y(_2925_));
 sky130_fd_sc_hd__o21ai_0 _5363_ (.A1(net1230),
    .A2(_2925_),
    .B1(net672),
    .Y(_2926_));
 sky130_fd_sc_hd__o21ai_0 _5364_ (.A1(net672),
    .A2(_2923_),
    .B1(_2926_),
    .Y(_0282_));
 sky130_fd_sc_hd__or3_1 _5365_ (.A(_2920_),
    .B(_2917_),
    .C(_2921_),
    .X(_2927_));
 sky130_fd_sc_hd__xnor2_1 _5366_ (.A(net683),
    .B(_2927_),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_1 _5367_ (.A(net683),
    .Y(_2928_));
 sky130_fd_sc_hd__a21oi_1 _5368_ (.A1(net1263),
    .A2(_2927_),
    .B1(net1230),
    .Y(_2929_));
 sky130_fd_sc_hd__or3_1 _5369_ (.A(net683),
    .B(_1869_),
    .C(_2927_),
    .X(_2930_));
 sky130_fd_sc_hd__o21ai_0 _5370_ (.A1(_2928_),
    .A2(_2929_),
    .B1(_2930_),
    .Y(_0283_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input63 (.A(net1473),
    .X(net63));
 sky130_fd_sc_hd__or4_1 _5372_ (.A(_2920_),
    .B(_2928_),
    .C(_2910_),
    .D(_2921_),
    .X(_2932_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input62 (.A(net1519),
    .X(net62));
 sky130_fd_sc_hd__xnor2_1 _5374_ (.A(net694),
    .B(_2932_),
    .Y(_0499_));
 sky130_fd_sc_hd__and2_0 _5375_ (.A(net1263),
    .B(_2932_),
    .X(_2934_));
 sky130_fd_sc_hd__o21ai_0 _5376_ (.A1(net1230),
    .A2(_2934_),
    .B1(net694),
    .Y(_2935_));
 sky130_fd_sc_hd__o31ai_1 _5377_ (.A1(net694),
    .A2(_1869_),
    .A3(_2932_),
    .B1(_2935_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand4_1 _5378_ (.A(net617),
    .B(_0403_),
    .C(net672),
    .D(net683),
    .Y(_2936_));
 sky130_fd_sc_hd__nor2_1 _5379_ (.A(_2921_),
    .B(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(net694),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__xnor2_1 _5381_ (.A(net578),
    .B(_2938_),
    .Y(_0495_));
 sky130_fd_sc_hd__a21oi_1 _5382_ (.A1(net694),
    .A2(_2937_),
    .B1(_1869_),
    .Y(_2939_));
 sky130_fd_sc_hd__o21ai_0 _5383_ (.A1(net1230),
    .A2(_2939_),
    .B1(net578),
    .Y(_2940_));
 sky130_fd_sc_hd__o31ai_1 _5384_ (.A1(net578),
    .A2(_1869_),
    .A3(_2938_),
    .B1(_2940_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _5385_ (.A(net694),
    .B(net578),
    .Y(_2941_));
 sky130_fd_sc_hd__nor2_1 _5386_ (.A(_2932_),
    .B(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__xor2_1 _5387_ (.A(net589),
    .B(_2942_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_1 _5388_ (.A(net1263),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__nor2_1 _5389_ (.A(_1869_),
    .B(_2942_),
    .Y(_2944_));
 sky130_fd_sc_hd__o21ai_0 _5390_ (.A1(net1230),
    .A2(_2944_),
    .B1(net589),
    .Y(_2945_));
 sky130_fd_sc_hd__o21ai_0 _5391_ (.A1(net589),
    .A2(_2943_),
    .B1(_2945_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand3_1 _5392_ (.A(net683),
    .B(net694),
    .C(net578),
    .Y(_2946_));
 sky130_fd_sc_hd__nor4_1 _5393_ (.A(_2920_),
    .B(_2917_),
    .C(_2921_),
    .D(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__nand2_1 _5394_ (.A(net589),
    .B(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__xnor2_1 _5395_ (.A(net598),
    .B(_2948_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21oi_1 _5396_ (.A1(net589),
    .A2(_2947_),
    .B1(_1869_),
    .Y(_2949_));
 sky130_fd_sc_hd__o21ai_0 _5397_ (.A1(net1230),
    .A2(_2949_),
    .B1(net598),
    .Y(_2950_));
 sky130_fd_sc_hd__o31ai_1 _5398_ (.A1(net598),
    .A2(_1869_),
    .A3(_2948_),
    .B1(_2950_),
    .Y(_0256_));
 sky130_fd_sc_hd__and3_1 _5399_ (.A(net589),
    .B(net598),
    .C(_2942_),
    .X(_2951_));
 sky130_fd_sc_hd__xor2_1 _5400_ (.A(net599),
    .B(_2951_),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _5401_ (.A1(net599),
    .A2(net1230),
    .B1(_0483_),
    .B2(net1263),
    .X(_0257_));
 sky130_fd_sc_hd__and4_1 _5402_ (.A(net589),
    .B(net598),
    .C(net599),
    .D(_2947_),
    .X(_2952_));
 sky130_fd_sc_hd__xor2_1 _5403_ (.A(net600),
    .B(_2952_),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(net1263),
    .B(_2952_),
    .Y(_2953_));
 sky130_fd_sc_hd__nor2_1 _5405_ (.A(_1869_),
    .B(_2952_),
    .Y(_2954_));
 sky130_fd_sc_hd__o21ai_0 _5406_ (.A1(net1230),
    .A2(_2954_),
    .B1(net600),
    .Y(_2955_));
 sky130_fd_sc_hd__o21ai_0 _5407_ (.A1(net600),
    .A2(_2953_),
    .B1(_2955_),
    .Y(_0258_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input61 (.A(net1459),
    .X(net61));
 sky130_fd_sc_hd__and4_1 _5409_ (.A(net589),
    .B(net598),
    .C(net599),
    .D(net600),
    .X(_2957_));
 sky130_fd_sc_hd__nand3_1 _5410_ (.A(net694),
    .B(net578),
    .C(_2957_),
    .Y(_2958_));
 sky130_fd_sc_hd__nor2_4 _5411_ (.A(_2932_),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__xor2_1 _5412_ (.A(net601),
    .B(_2959_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(net1263),
    .B(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__nor2_1 _5414_ (.A(_1869_),
    .B(_2959_),
    .Y(_2961_));
 sky130_fd_sc_hd__o21ai_0 _5415_ (.A1(net1230),
    .A2(_2961_),
    .B1(net601),
    .Y(_2962_));
 sky130_fd_sc_hd__o21ai_0 _5416_ (.A1(net601),
    .A2(_2960_),
    .B1(_2962_),
    .Y(_0259_));
 sky130_fd_sc_hd__and3_1 _5417_ (.A(net601),
    .B(_2947_),
    .C(_2957_),
    .X(_2963_));
 sky130_fd_sc_hd__xor2_1 _5418_ (.A(net602),
    .B(_2963_),
    .X(_0471_));
 sky130_fd_sc_hd__nand2_1 _5419_ (.A(net1263),
    .B(_2963_),
    .Y(_2964_));
 sky130_fd_sc_hd__nor2_1 _5420_ (.A(_1869_),
    .B(_2963_),
    .Y(_2965_));
 sky130_fd_sc_hd__o21ai_0 _5421_ (.A1(net1230),
    .A2(_2965_),
    .B1(net602),
    .Y(_2966_));
 sky130_fd_sc_hd__o21ai_0 _5422_ (.A1(net602),
    .A2(_2964_),
    .B1(_2966_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand3_1 _5423_ (.A(net601),
    .B(net602),
    .C(_2959_),
    .Y(_2967_));
 sky130_fd_sc_hd__xnor2_1 _5424_ (.A(net603),
    .B(_2967_),
    .Y(_0467_));
 sky130_fd_sc_hd__a31oi_1 _5425_ (.A1(net601),
    .A2(net602),
    .A3(_2959_),
    .B1(_1869_),
    .Y(_2968_));
 sky130_fd_sc_hd__o21ai_0 _5426_ (.A1(net1230),
    .A2(_2968_),
    .B1(net603),
    .Y(_2969_));
 sky130_fd_sc_hd__o31ai_1 _5427_ (.A1(net603),
    .A2(_1869_),
    .A3(_2967_),
    .B1(_2969_),
    .Y(_0261_));
 sky130_fd_sc_hd__or4b_1 _5428_ (.A(_2921_),
    .B(_2936_),
    .C(_2941_),
    .D_N(_2957_),
    .X(_2970_));
 sky130_fd_sc_hd__nand3_1 _5429_ (.A(net601),
    .B(net602),
    .C(net603),
    .Y(_2971_));
 sky130_fd_sc_hd__nor2_1 _5430_ (.A(_2970_),
    .B(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__xor2_1 _5431_ (.A(net604),
    .B(_2972_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _5432_ (.A(net1263),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__nor2_1 _5433_ (.A(_1869_),
    .B(_2972_),
    .Y(_2974_));
 sky130_fd_sc_hd__o21ai_0 _5434_ (.A1(net1230),
    .A2(_2974_),
    .B1(net604),
    .Y(_2975_));
 sky130_fd_sc_hd__o21ai_0 _5435_ (.A1(net604),
    .A2(_2973_),
    .B1(_2975_),
    .Y(_0262_));
 sky130_fd_sc_hd__and4_1 _5436_ (.A(net601),
    .B(net602),
    .C(net603),
    .D(net604),
    .X(_2976_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input60 (.A(net1581),
    .X(net60));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_2959_),
    .B(_2976_),
    .Y(_2978_));
 sky130_fd_sc_hd__xnor2_1 _5439_ (.A(net605),
    .B(_2978_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21oi_1 _5440_ (.A1(_2959_),
    .A2(_2976_),
    .B1(_1869_),
    .Y(_2979_));
 sky130_fd_sc_hd__o21ai_0 _5441_ (.A1(_2896_),
    .A2(_2979_),
    .B1(net605),
    .Y(_2980_));
 sky130_fd_sc_hd__o31ai_1 _5442_ (.A1(net605),
    .A2(_1869_),
    .A3(_2978_),
    .B1(_2980_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _5443_ (.A(net605),
    .B(_2976_),
    .Y(_2981_));
 sky130_fd_sc_hd__nor2_1 _5444_ (.A(_2970_),
    .B(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__xor2_1 _5445_ (.A(net607),
    .B(_2982_),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _5446_ (.A(net1263),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__nor2_1 _5447_ (.A(_1869_),
    .B(_2982_),
    .Y(_2984_));
 sky130_fd_sc_hd__o21ai_0 _5448_ (.A1(_2896_),
    .A2(_2984_),
    .B1(net607),
    .Y(_2985_));
 sky130_fd_sc_hd__o21ai_0 _5449_ (.A1(net607),
    .A2(_2983_),
    .B1(_2985_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand4_1 _5450_ (.A(net605),
    .B(net607),
    .C(_2959_),
    .D(_2976_),
    .Y(_2986_));
 sky130_fd_sc_hd__xnor2_1 _5451_ (.A(net608),
    .B(_2986_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_1 _5452_ (.A(net608),
    .Y(_2987_));
 sky130_fd_sc_hd__a21oi_1 _5453_ (.A1(net1263),
    .A2(_2986_),
    .B1(_2896_),
    .Y(_2988_));
 sky130_fd_sc_hd__or3_1 _5454_ (.A(net608),
    .B(_1869_),
    .C(_2986_),
    .X(_2989_));
 sky130_fd_sc_hd__o21ai_0 _5455_ (.A1(_2987_),
    .A2(_2988_),
    .B1(_2989_),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_1 _5456_ (.A(net609),
    .Y(_2990_));
 sky130_fd_sc_hd__and3_1 _5457_ (.A(net605),
    .B(net607),
    .C(net608),
    .X(_2991_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_2976_),
    .B(_2991_),
    .Y(_2992_));
 sky130_fd_sc_hd__nor2_1 _5459_ (.A(_2970_),
    .B(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__xnor2_1 _5460_ (.A(_2990_),
    .B(_2993_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_1 _5461_ (.A(net1263),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__nor2_1 _5462_ (.A(_1869_),
    .B(_2993_),
    .Y(_2995_));
 sky130_fd_sc_hd__o21ai_0 _5463_ (.A1(_2896_),
    .A2(_2995_),
    .B1(net609),
    .Y(_2996_));
 sky130_fd_sc_hd__o21ai_0 _5464_ (.A1(net609),
    .A2(_2994_),
    .B1(_2996_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor4_1 _5465_ (.A(_2990_),
    .B(_2932_),
    .C(_2958_),
    .D(_2992_),
    .Y(_2997_));
 sky130_fd_sc_hd__xor2_1 _5466_ (.A(net610),
    .B(_2997_),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(net1263),
    .B(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__nor2_1 _5468_ (.A(_1869_),
    .B(_2997_),
    .Y(_2999_));
 sky130_fd_sc_hd__o21ai_0 _5469_ (.A1(_2896_),
    .A2(_2999_),
    .B1(net610),
    .Y(_3000_));
 sky130_fd_sc_hd__o21ai_0 _5470_ (.A1(net610),
    .A2(_2998_),
    .B1(_3000_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand3_1 _5471_ (.A(net609),
    .B(net610),
    .C(_2993_),
    .Y(_3001_));
 sky130_fd_sc_hd__xnor2_1 _5472_ (.A(net611),
    .B(_3001_),
    .Y(_0439_));
 sky130_fd_sc_hd__a31oi_1 _5473_ (.A1(net609),
    .A2(net610),
    .A3(_2993_),
    .B1(_1869_),
    .Y(_3002_));
 sky130_fd_sc_hd__o21ai_0 _5474_ (.A1(_2896_),
    .A2(_3002_),
    .B1(net611),
    .Y(_3003_));
 sky130_fd_sc_hd__o31ai_1 _5475_ (.A1(net611),
    .A2(_1869_),
    .A3(_3001_),
    .B1(_3003_),
    .Y(_0269_));
 sky130_fd_sc_hd__and3_1 _5476_ (.A(net609),
    .B(net610),
    .C(net611),
    .X(_3004_));
 sky130_fd_sc_hd__or4b_4 _5477_ (.A(_2932_),
    .B(_2958_),
    .C(_2992_),
    .D_N(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__xnor2_1 _5478_ (.A(net612),
    .B(_3005_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21o_1 _5479_ (.A1(net1263),
    .A2(_3005_),
    .B1(_2896_),
    .X(_3006_));
 sky130_fd_sc_hd__nand2_1 _5480_ (.A(net612),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__o31ai_1 _5481_ (.A1(net612),
    .A2(_1869_),
    .A3(_3005_),
    .B1(_3007_),
    .Y(_0270_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input59 (.A(net1643),
    .X(net59));
 sky130_fd_sc_hd__nand4_1 _5483_ (.A(net612),
    .B(_2976_),
    .C(_2991_),
    .D(_3004_),
    .Y(_3009_));
 sky130_fd_sc_hd__nor2_1 _5484_ (.A(_2970_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__xor2_1 _5485_ (.A(net613),
    .B(_3010_),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(net1263),
    .B(_3010_),
    .Y(_3011_));
 sky130_fd_sc_hd__nor2_1 _5487_ (.A(_1869_),
    .B(_3010_),
    .Y(_3012_));
 sky130_fd_sc_hd__o21ai_0 _5488_ (.A1(_2896_),
    .A2(_3012_),
    .B1(net613),
    .Y(_3013_));
 sky130_fd_sc_hd__o21ai_0 _5489_ (.A1(net613),
    .A2(_3011_),
    .B1(_3013_),
    .Y(_0271_));
 sky130_fd_sc_hd__nor3_4 _5490_ (.A(_2932_),
    .B(_2958_),
    .C(_3009_),
    .Y(_3014_));
 sky130_fd_sc_hd__nand2_1 _5491_ (.A(net613),
    .B(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__xnor2_1 _5492_ (.A(net614),
    .B(_3015_),
    .Y(_0427_));
 sky130_fd_sc_hd__a21oi_1 _5493_ (.A1(net613),
    .A2(_3014_),
    .B1(_1869_),
    .Y(_3016_));
 sky130_fd_sc_hd__o21ai_0 _5494_ (.A1(_2896_),
    .A2(_3016_),
    .B1(net614),
    .Y(_3017_));
 sky130_fd_sc_hd__o31ai_1 _5495_ (.A1(net614),
    .A2(_1869_),
    .A3(_3015_),
    .B1(_3017_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand3_1 _5496_ (.A(net613),
    .B(net614),
    .C(_3010_),
    .Y(_3018_));
 sky130_fd_sc_hd__xnor2_1 _5497_ (.A(net615),
    .B(_3018_),
    .Y(_0423_));
 sky130_fd_sc_hd__a31oi_1 _5498_ (.A1(net613),
    .A2(net614),
    .A3(_3010_),
    .B1(_1869_),
    .Y(_3019_));
 sky130_fd_sc_hd__o21ai_0 _5499_ (.A1(_2896_),
    .A2(_3019_),
    .B1(net615),
    .Y(_3020_));
 sky130_fd_sc_hd__o31ai_1 _5500_ (.A1(net615),
    .A2(_1869_),
    .A3(_3018_),
    .B1(_3020_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand4_1 _5501_ (.A(net613),
    .B(net614),
    .C(net615),
    .D(_3014_),
    .Y(_3021_));
 sky130_fd_sc_hd__xnor2_1 _5502_ (.A(net616),
    .B(_3021_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_1 _5503_ (.A(net616),
    .Y(_3022_));
 sky130_fd_sc_hd__a21oi_1 _5504_ (.A1(net1263),
    .A2(_3021_),
    .B1(_2896_),
    .Y(_3023_));
 sky130_fd_sc_hd__or3_1 _5505_ (.A(net616),
    .B(_1869_),
    .C(_3021_),
    .X(_3024_));
 sky130_fd_sc_hd__o21ai_0 _5506_ (.A1(_3022_),
    .A2(_3023_),
    .B1(_3024_),
    .Y(_0274_));
 sky130_fd_sc_hd__and4_1 _5507_ (.A(net613),
    .B(net614),
    .C(net615),
    .D(net616),
    .X(_3025_));
 sky130_fd_sc_hd__nand2_1 _5508_ (.A(_3010_),
    .B(_3025_),
    .Y(_3026_));
 sky130_fd_sc_hd__xnor2_1 _5509_ (.A(net618),
    .B(_3026_),
    .Y(_0415_));
 sky130_fd_sc_hd__a21oi_1 _5510_ (.A1(_3010_),
    .A2(_3025_),
    .B1(_1869_),
    .Y(_3027_));
 sky130_fd_sc_hd__o21ai_0 _5511_ (.A1(_2896_),
    .A2(_3027_),
    .B1(net618),
    .Y(_3028_));
 sky130_fd_sc_hd__o31ai_1 _5512_ (.A1(net618),
    .A2(_1869_),
    .A3(_3026_),
    .B1(_3028_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand3_1 _5513_ (.A(net618),
    .B(_3014_),
    .C(_3025_),
    .Y(_3029_));
 sky130_fd_sc_hd__xnor2_1 _5514_ (.A(net619),
    .B(_3029_),
    .Y(_0411_));
 sky130_fd_sc_hd__a31oi_1 _5515_ (.A1(net618),
    .A2(_3014_),
    .A3(_3025_),
    .B1(_1869_),
    .Y(_3030_));
 sky130_fd_sc_hd__o21ai_0 _5516_ (.A1(_2896_),
    .A2(_3030_),
    .B1(net619),
    .Y(_3031_));
 sky130_fd_sc_hd__o31ai_1 _5517_ (.A1(net619),
    .A2(_1869_),
    .A3(_3029_),
    .B1(_3031_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_1 _5518_ (.A(\active_channel_count[0] ),
    .Y(_0405_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input58 (.A(net1628),
    .X(net58));
 sky130_fd_sc_hd__xor2_1 _5520_ (.A(net554),
    .B(net557),
    .X(_3033_));
 sky130_fd_sc_hd__nand2_1 _5521_ (.A(net129),
    .B(net538),
    .Y(_3034_));
 sky130_fd_sc_hd__a21oi_2 _5522_ (.A1(net558),
    .A2(_3033_),
    .B1(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input57 (.A(net1342),
    .X(net57));
 sky130_fd_sc_hd__xor2_1 _5524_ (.A(net1273),
    .B(net1272),
    .X(_3037_));
 sky130_fd_sc_hd__nand2_1 _5525_ (.A(net130),
    .B(net539),
    .Y(_3038_));
 sky130_fd_sc_hd__a21oi_1 _5526_ (.A1(net1271),
    .A2(_3037_),
    .B1(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input56 (.A(net1582),
    .X(net56));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input55 (.A(net1299),
    .X(net55));
 sky130_fd_sc_hd__xor2_1 _5529_ (.A(net555),
    .B(net565),
    .X(_3042_));
 sky130_fd_sc_hd__nand2_1 _5530_ (.A(net132),
    .B(net541),
    .Y(_3043_));
 sky130_fd_sc_hd__a21oi_1 _5531_ (.A1(net556),
    .A2(_3042_),
    .B1(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input54 (.A(net1302),
    .X(net54));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input53 (.A(channel_dst_addr[31]),
    .X(net53));
 sky130_fd_sc_hd__xor2_1 _5534_ (.A(net563),
    .B(net562),
    .X(_3047_));
 sky130_fd_sc_hd__nand2_1 _5535_ (.A(net131),
    .B(net540),
    .Y(_3048_));
 sky130_fd_sc_hd__a21oi_2 _5536_ (.A1(net564),
    .A2(_3047_),
    .B1(_3048_),
    .Y(_3049_));
 sky130_fd_sc_hd__nor4_1 _5537_ (.A(net1240),
    .B(_3039_),
    .C(_3044_),
    .D(net1239),
    .Y(_3050_));
 sky130_fd_sc_hd__nor2_1 _5538_ (.A(\active_channel_count[0] ),
    .B(_3050_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2b_1 _5539_ (.A(_3050_),
    .B_N(_0408_),
    .Y(_0001_));
 sky130_fd_sc_hd__xnor2_1 _5540_ (.A(_0409_),
    .B(\active_channel_count[2] ),
    .Y(_3051_));
 sky130_fd_sc_hd__nor2_1 _5541_ (.A(_3050_),
    .B(_3051_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand3_1 _5542_ (.A(\active_channel_count[0] ),
    .B(\active_channel_count[2] ),
    .C(\active_channel_count[1] ),
    .Y(_3052_));
 sky130_fd_sc_hd__xor2_1 _5543_ (.A(\active_channel_count[3] ),
    .B(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__nor2_1 _5544_ (.A(_3050_),
    .B(_3053_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand3_1 _5545_ (.A(_0477_),
    .B(_0485_),
    .C(_0481_),
    .Y(_3054_));
 sky130_fd_sc_hd__a211oi_1 _5546_ (.A1(_0501_),
    .A2(_0504_),
    .B1(_0500_),
    .C1(_0496_),
    .Y(_3055_));
 sky130_fd_sc_hd__o21ai_0 _5547_ (.A1(_0497_),
    .A2(_0496_),
    .B1(_0493_),
    .Y(_3056_));
 sky130_fd_sc_hd__o21bai_1 _5548_ (.A1(_3055_),
    .A2(_3056_),
    .B1_N(_0492_),
    .Y(_3057_));
 sky130_fd_sc_hd__a21oi_1 _5549_ (.A1(_0489_),
    .A2(_3057_),
    .B1(_0488_),
    .Y(_3058_));
 sky130_fd_sc_hd__nor2_1 _5550_ (.A(_3054_),
    .B(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__a21oi_1 _5551_ (.A1(_0521_),
    .A2(_0524_),
    .B1(_0520_),
    .Y(_3060_));
 sky130_fd_sc_hd__nor2b_1 _5552_ (.A(_0534_),
    .B_N(_0533_),
    .Y(_3061_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_0532_),
    .B(_0529_),
    .Y(_3062_));
 sky130_fd_sc_hd__a21oi_1 _5554_ (.A1(_0529_),
    .A2(_0531_),
    .B1(_0528_),
    .Y(_3063_));
 sky130_fd_sc_hd__o21ai_0 _5555_ (.A1(_3061_),
    .A2(_3062_),
    .B1(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__nand3_1 _5556_ (.A(_0521_),
    .B(_0525_),
    .C(_3064_),
    .Y(_3065_));
 sky130_fd_sc_hd__nand4_1 _5557_ (.A(_0493_),
    .B(_0505_),
    .C(_0501_),
    .D(_0497_),
    .Y(_3066_));
 sky130_fd_sc_hd__nor2_1 _5558_ (.A(_3054_),
    .B(_3066_),
    .Y(_3067_));
 sky130_fd_sc_hd__nand2_1 _5559_ (.A(_0489_),
    .B(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__nand3_1 _5560_ (.A(_0509_),
    .B(_0517_),
    .C(_0513_),
    .Y(_3069_));
 sky130_fd_sc_hd__a211oi_1 _5561_ (.A1(_3060_),
    .A2(_3065_),
    .B1(_3068_),
    .C1(_3069_),
    .Y(_3070_));
 sky130_fd_sc_hd__a21o_1 _5562_ (.A1(_0513_),
    .A2(_0516_),
    .B1(_0512_),
    .X(_3071_));
 sky130_fd_sc_hd__a21oi_1 _5563_ (.A1(_0509_),
    .A2(_3071_),
    .B1(_0508_),
    .Y(_3072_));
 sky130_fd_sc_hd__a21o_1 _5564_ (.A1(_0481_),
    .A2(_0484_),
    .B1(_0480_),
    .X(_3073_));
 sky130_fd_sc_hd__a21oi_1 _5565_ (.A1(_0477_),
    .A2(_3073_),
    .B1(_0476_),
    .Y(_3074_));
 sky130_fd_sc_hd__o21ai_0 _5566_ (.A1(_3068_),
    .A2(_3072_),
    .B1(_3074_),
    .Y(_3075_));
 sky130_fd_sc_hd__nand4_1 _5567_ (.A(_0429_),
    .B(_0441_),
    .C(_0437_),
    .D(_0433_),
    .Y(_3076_));
 sky130_fd_sc_hd__nand4_1 _5568_ (.A(_0461_),
    .B(_0473_),
    .C(_0469_),
    .D(_0465_),
    .Y(_3077_));
 sky130_fd_sc_hd__nand4_1 _5569_ (.A(_0445_),
    .B(_0457_),
    .C(_0453_),
    .D(_0449_),
    .Y(_3078_));
 sky130_fd_sc_hd__nand4_1 _5570_ (.A(_0413_),
    .B(_0425_),
    .C(_0421_),
    .D(_0417_),
    .Y(_3079_));
 sky130_fd_sc_hd__nor4_1 _5571_ (.A(_3076_),
    .B(_3077_),
    .C(_3078_),
    .D(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__o31ai_1 _5572_ (.A1(_3059_),
    .A2(_3070_),
    .A3(_3075_),
    .B1(_3080_),
    .Y(_3081_));
 sky130_fd_sc_hd__inv_1 _5573_ (.A(net397),
    .Y(_3082_));
 sky130_fd_sc_hd__and3_1 _5574_ (.A(net397),
    .B(net129),
    .C(_1865_),
    .X(_3083_));
 sky130_fd_sc_hd__a31oi_1 _5575_ (.A1(net558),
    .A2(net554),
    .A3(_3082_),
    .B1(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__o21a_1 _5576_ (.A1(net557),
    .A2(_3084_),
    .B1(net542),
    .X(_3085_));
 sky130_fd_sc_hd__nand2_1 _5577_ (.A(_0445_),
    .B(_0449_),
    .Y(_3086_));
 sky130_fd_sc_hd__nand2_1 _5578_ (.A(_0457_),
    .B(_0453_),
    .Y(_3087_));
 sky130_fd_sc_hd__nor2_1 _5579_ (.A(_3086_),
    .B(_3087_),
    .Y(_3088_));
 sky130_fd_sc_hd__nand2_1 _5580_ (.A(_0461_),
    .B(_0465_),
    .Y(_3089_));
 sky130_fd_sc_hd__a21oi_1 _5581_ (.A1(_0469_),
    .A2(_0472_),
    .B1(_0468_),
    .Y(_3090_));
 sky130_fd_sc_hd__a21oi_1 _5582_ (.A1(_0461_),
    .A2(_0464_),
    .B1(_0460_),
    .Y(_3091_));
 sky130_fd_sc_hd__o21ai_0 _5583_ (.A1(_3089_),
    .A2(_3090_),
    .B1(_3091_),
    .Y(_3092_));
 sky130_fd_sc_hd__a21oi_1 _5584_ (.A1(_0453_),
    .A2(_0456_),
    .B1(_0452_),
    .Y(_3093_));
 sky130_fd_sc_hd__a21oi_1 _5585_ (.A1(_0445_),
    .A2(_0448_),
    .B1(_0444_),
    .Y(_3094_));
 sky130_fd_sc_hd__o21ai_0 _5586_ (.A1(_3086_),
    .A2(_3093_),
    .B1(_3094_),
    .Y(_3095_));
 sky130_fd_sc_hd__nand2_1 _5587_ (.A(_0429_),
    .B(_0433_),
    .Y(_3096_));
 sky130_fd_sc_hd__a21oi_1 _5588_ (.A1(_0437_),
    .A2(_0440_),
    .B1(_0436_),
    .Y(_3097_));
 sky130_fd_sc_hd__a21oi_1 _5589_ (.A1(_0429_),
    .A2(_0432_),
    .B1(_0428_),
    .Y(_3098_));
 sky130_fd_sc_hd__o21ai_0 _5590_ (.A1(_3096_),
    .A2(_3097_),
    .B1(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__a211oi_1 _5591_ (.A1(_3088_),
    .A2(_3092_),
    .B1(_3095_),
    .C1(_3099_),
    .Y(_3100_));
 sky130_fd_sc_hd__nor2b_1 _5592_ (.A(_3099_),
    .B_N(_3076_),
    .Y(_3101_));
 sky130_fd_sc_hd__nor3_1 _5593_ (.A(_3079_),
    .B(_3100_),
    .C(_3101_),
    .Y(_3102_));
 sky130_fd_sc_hd__a21oi_1 _5594_ (.A1(_0421_),
    .A2(_0424_),
    .B1(_0420_),
    .Y(_3103_));
 sky130_fd_sc_hd__nor2b_1 _5595_ (.A(_3103_),
    .B_N(_0417_),
    .Y(_3104_));
 sky130_fd_sc_hd__o21ai_0 _5596_ (.A1(_0416_),
    .A2(_3104_),
    .B1(_0413_),
    .Y(_3105_));
 sky130_fd_sc_hd__nand2b_1 _5597_ (.A_N(_0412_),
    .B(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__nor3_1 _5598_ (.A(_3085_),
    .B(_3102_),
    .C(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__nor2_1 _5599_ (.A(net1263),
    .B(_3085_),
    .Y(_3108_));
 sky130_fd_sc_hd__a21oi_1 _5600_ (.A1(_3081_),
    .A2(_3107_),
    .B1(_3108_),
    .Y(_3428_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(net1271),
    .B(net1273),
    .Y(_3109_));
 sky130_fd_sc_hd__nor2_1 _5602_ (.A(net398),
    .B(_3109_),
    .Y(_3110_));
 sky130_fd_sc_hd__a31oi_1 _5603_ (.A1(net398),
    .A2(net130),
    .A3(_1732_),
    .B1(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__o21ai_0 _5604_ (.A1(net1272),
    .A2(_3111_),
    .B1(net543),
    .Y(_3112_));
 sky130_fd_sc_hd__a21oi_1 _5605_ (.A1(_0607_),
    .A2(_0610_),
    .B1(_0606_),
    .Y(_3113_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_0599_),
    .B(_0603_),
    .Y(_3114_));
 sky130_fd_sc_hd__a21oi_1 _5607_ (.A1(_0599_),
    .A2(_0602_),
    .B1(_0598_),
    .Y(_3115_));
 sky130_fd_sc_hd__o21a_1 _5608_ (.A1(_0635_),
    .A2(_0634_),
    .B1(_0631_),
    .X(_3116_));
 sky130_fd_sc_hd__nand4_1 _5609_ (.A(_0643_),
    .B(_0639_),
    .C(_0647_),
    .D(_0651_),
    .Y(_3117_));
 sky130_fd_sc_hd__a21oi_1 _5610_ (.A1(_0655_),
    .A2(_0658_),
    .B1(_0654_),
    .Y(_3118_));
 sky130_fd_sc_hd__nand2_1 _5611_ (.A(_0631_),
    .B(_0634_),
    .Y(_3119_));
 sky130_fd_sc_hd__a211oi_1 _5612_ (.A1(_0639_),
    .A2(_0642_),
    .B1(_0638_),
    .C1(_0630_),
    .Y(_3120_));
 sky130_fd_sc_hd__o211ai_1 _5613_ (.A1(_3117_),
    .A2(_3118_),
    .B1(_3119_),
    .C1(_3120_),
    .Y(_3121_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(_0643_),
    .B(_0639_),
    .Y(_3122_));
 sky130_fd_sc_hd__a21oi_1 _5615_ (.A1(_0647_),
    .A2(_0650_),
    .B1(_0646_),
    .Y(_3123_));
 sky130_fd_sc_hd__nor2_1 _5616_ (.A(_3122_),
    .B(_3123_),
    .Y(_3124_));
 sky130_fd_sc_hd__nand4_1 _5617_ (.A(_0599_),
    .B(_0611_),
    .C(_0607_),
    .D(_0603_),
    .Y(_3125_));
 sky130_fd_sc_hd__nand2_1 _5618_ (.A(_0615_),
    .B(_0619_),
    .Y(_3126_));
 sky130_fd_sc_hd__nand2_1 _5619_ (.A(_0627_),
    .B(_0623_),
    .Y(_3127_));
 sky130_fd_sc_hd__nor3_1 _5620_ (.A(_3125_),
    .B(_3126_),
    .C(_3127_),
    .Y(_3128_));
 sky130_fd_sc_hd__o221ai_1 _5621_ (.A1(_0630_),
    .A2(_3116_),
    .B1(_3121_),
    .B2(_3124_),
    .C1(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__a21oi_1 _5622_ (.A1(_0623_),
    .A2(_0626_),
    .B1(_0622_),
    .Y(_3130_));
 sky130_fd_sc_hd__a21oi_1 _5623_ (.A1(_0615_),
    .A2(_0618_),
    .B1(_0614_),
    .Y(_3131_));
 sky130_fd_sc_hd__o21ai_0 _5624_ (.A1(_3130_),
    .A2(_3126_),
    .B1(_3131_),
    .Y(_3132_));
 sky130_fd_sc_hd__nand2b_1 _5625_ (.A_N(_3125_),
    .B(_3132_),
    .Y(_3133_));
 sky130_fd_sc_hd__o2111ai_1 _5626_ (.A1(_3113_),
    .A2(_3114_),
    .B1(_3115_),
    .C1(_3129_),
    .D1(_3133_),
    .Y(_3134_));
 sky130_fd_sc_hd__and4_1 _5627_ (.A(_0583_),
    .B(_0595_),
    .C(_0591_),
    .D(_0587_),
    .X(_3135_));
 sky130_fd_sc_hd__a21oi_1 _5628_ (.A1(_0559_),
    .A2(_0562_),
    .B1(_0558_),
    .Y(_3136_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(_0551_),
    .B(_0555_),
    .Y(_3137_));
 sky130_fd_sc_hd__a21oi_1 _5630_ (.A1(_0551_),
    .A2(_0554_),
    .B1(_0550_),
    .Y(_3138_));
 sky130_fd_sc_hd__o21ai_0 _5631_ (.A1(_3136_),
    .A2(_3137_),
    .B1(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__nand2_1 _5632_ (.A(_3135_),
    .B(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hd__inv_1 _5633_ (.A(_0542_),
    .Y(_3141_));
 sky130_fd_sc_hd__o21ai_0 _5634_ (.A1(_0547_),
    .A2(_0546_),
    .B1(_0543_),
    .Y(_3142_));
 sky130_fd_sc_hd__inv_1 _5635_ (.A(_0535_),
    .Y(_3143_));
 sky130_fd_sc_hd__o21ai_0 _5636_ (.A1(_0536_),
    .A2(_3143_),
    .B1(_0539_),
    .Y(_3144_));
 sky130_fd_sc_hd__nor3_1 _5637_ (.A(_0538_),
    .B(_0542_),
    .C(_0546_),
    .Y(_3145_));
 sky130_fd_sc_hd__and4_1 _5638_ (.A(_0551_),
    .B(_0563_),
    .C(_0559_),
    .D(_0555_),
    .X(_3146_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_3135_),
    .B(_3146_),
    .Y(_3147_));
 sky130_fd_sc_hd__a221o_1 _5640_ (.A1(_3141_),
    .A2(_3142_),
    .B1(_3144_),
    .B2(_3145_),
    .C1(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__a21oi_1 _5641_ (.A1(_0575_),
    .A2(_0578_),
    .B1(_0574_),
    .Y(_3149_));
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(_0567_),
    .B(_0571_),
    .Y(_3150_));
 sky130_fd_sc_hd__a21oi_1 _5643_ (.A1(_0567_),
    .A2(_0570_),
    .B1(_0566_),
    .Y(_3151_));
 sky130_fd_sc_hd__o21ai_0 _5644_ (.A1(_3149_),
    .A2(_3150_),
    .B1(_3151_),
    .Y(_3152_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(_0583_),
    .B(_0587_),
    .Y(_3153_));
 sky130_fd_sc_hd__a21oi_1 _5646_ (.A1(_0591_),
    .A2(_0594_),
    .B1(_0590_),
    .Y(_3154_));
 sky130_fd_sc_hd__nor2_1 _5647_ (.A(_3153_),
    .B(_3154_),
    .Y(_3155_));
 sky130_fd_sc_hd__a2111oi_0 _5648_ (.A1(_0583_),
    .A2(_0586_),
    .B1(_3152_),
    .C1(_3155_),
    .D1(_0582_),
    .Y(_3156_));
 sky130_fd_sc_hd__a41oi_1 _5649_ (.A1(_0567_),
    .A2(_0579_),
    .A3(_0575_),
    .A4(_0571_),
    .B1(_3152_),
    .Y(_3157_));
 sky130_fd_sc_hd__nand4_1 _5650_ (.A(_0631_),
    .B(_0659_),
    .C(_0655_),
    .D(_0635_),
    .Y(_3158_));
 sky130_fd_sc_hd__nor2_1 _5651_ (.A(_3117_),
    .B(_3158_),
    .Y(_3159_));
 sky130_fd_sc_hd__nand2_1 _5652_ (.A(_3128_),
    .B(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__a311oi_1 _5653_ (.A1(_3140_),
    .A2(_3148_),
    .A3(_3156_),
    .B1(_3157_),
    .C1(_3160_),
    .Y(_3161_));
 sky130_fd_sc_hd__o21ai_0 _5654_ (.A1(_3134_),
    .A2(_3161_),
    .B1(net1264),
    .Y(_3162_));
 sky130_fd_sc_hd__nand2_1 _5655_ (.A(_3112_),
    .B(_3162_),
    .Y(_3426_));
 sky130_fd_sc_hd__nand4_1 _5656_ (.A(_0724_),
    .B(_0736_),
    .C(_0732_),
    .D(_0728_),
    .Y(_3163_));
 sky130_fd_sc_hd__nand4_1 _5657_ (.A(_0740_),
    .B(_0752_),
    .C(_0748_),
    .D(_0744_),
    .Y(_3164_));
 sky130_fd_sc_hd__nand2_1 _5658_ (.A(_0756_),
    .B(_0760_),
    .Y(_3165_));
 sky130_fd_sc_hd__nor3_1 _5659_ (.A(_3163_),
    .B(_3164_),
    .C(_3165_),
    .Y(_3166_));
 sky130_fd_sc_hd__o21ai_0 _5660_ (.A1(_0704_),
    .A2(_0703_),
    .B1(_0700_),
    .Y(_3167_));
 sky130_fd_sc_hd__nor2_1 _5661_ (.A(_0695_),
    .B(_0699_),
    .Y(_3168_));
 sky130_fd_sc_hd__o21ai_0 _5662_ (.A1(_0696_),
    .A2(_0695_),
    .B1(_0692_),
    .Y(_3169_));
 sky130_fd_sc_hd__a21oi_1 _5663_ (.A1(_3167_),
    .A2(_3168_),
    .B1(_3169_),
    .Y(_3170_));
 sky130_fd_sc_hd__or2_2 _5664_ (.A(_0691_),
    .B(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__nand4_1 _5665_ (.A(_0708_),
    .B(_0720_),
    .C(_0716_),
    .D(_0712_),
    .Y(_3172_));
 sky130_fd_sc_hd__nor2b_1 _5666_ (.A(_0661_),
    .B_N(_0660_),
    .Y(_3173_));
 sky130_fd_sc_hd__nand2_1 _5667_ (.A(_0664_),
    .B(_0672_),
    .Y(_3174_));
 sky130_fd_sc_hd__a211oi_1 _5668_ (.A1(_0672_),
    .A2(_0663_),
    .B1(_0667_),
    .C1(_0671_),
    .Y(_3175_));
 sky130_fd_sc_hd__o21ai_0 _5669_ (.A1(_3173_),
    .A2(_3174_),
    .B1(_3175_),
    .Y(_3176_));
 sky130_fd_sc_hd__nand2_1 _5670_ (.A(_0676_),
    .B(_0680_),
    .Y(_3177_));
 sky130_fd_sc_hd__nand2_1 _5671_ (.A(_0688_),
    .B(_0684_),
    .Y(_3178_));
 sky130_fd_sc_hd__nor2_1 _5672_ (.A(_0668_),
    .B(_0667_),
    .Y(_3179_));
 sky130_fd_sc_hd__nor3_1 _5673_ (.A(_3177_),
    .B(_3178_),
    .C(_3179_),
    .Y(_3180_));
 sky130_fd_sc_hd__a21oi_1 _5674_ (.A1(_0684_),
    .A2(_0687_),
    .B1(_0683_),
    .Y(_3181_));
 sky130_fd_sc_hd__a21oi_1 _5675_ (.A1(_0676_),
    .A2(_0679_),
    .B1(_0675_),
    .Y(_3182_));
 sky130_fd_sc_hd__o21ai_0 _5676_ (.A1(_3181_),
    .A2(_3177_),
    .B1(_3182_),
    .Y(_3183_));
 sky130_fd_sc_hd__a21oi_1 _5677_ (.A1(_3176_),
    .A2(_3180_),
    .B1(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__a21o_1 _5678_ (.A1(_0716_),
    .A2(_0719_),
    .B1(_0715_),
    .X(_3185_));
 sky130_fd_sc_hd__a21o_1 _5679_ (.A1(_0712_),
    .A2(_3185_),
    .B1(_0711_),
    .X(_3186_));
 sky130_fd_sc_hd__a21oi_1 _5680_ (.A1(_0700_),
    .A2(_0703_),
    .B1(_0699_),
    .Y(_3187_));
 sky130_fd_sc_hd__nand2_1 _5681_ (.A(_0692_),
    .B(_0696_),
    .Y(_3188_));
 sky130_fd_sc_hd__a211oi_1 _5682_ (.A1(_0692_),
    .A2(_0695_),
    .B1(_0707_),
    .C1(_0691_),
    .Y(_3189_));
 sky130_fd_sc_hd__o21ai_0 _5683_ (.A1(_3187_),
    .A2(_3188_),
    .B1(_3189_),
    .Y(_3190_));
 sky130_fd_sc_hd__a21oi_1 _5684_ (.A1(_0708_),
    .A2(_3186_),
    .B1(_3190_),
    .Y(_3191_));
 sky130_fd_sc_hd__o21ai_0 _5685_ (.A1(_3172_),
    .A2(_3184_),
    .B1(_3191_),
    .Y(_3192_));
 sky130_fd_sc_hd__nand3_1 _5686_ (.A(_0768_),
    .B(_0772_),
    .C(_0776_),
    .Y(_3193_));
 sky130_fd_sc_hd__nand3_1 _5687_ (.A(_0764_),
    .B(_0784_),
    .C(_0780_),
    .Y(_3194_));
 sky130_fd_sc_hd__nor2_1 _5688_ (.A(_3193_),
    .B(_3194_),
    .Y(_3195_));
 sky130_fd_sc_hd__a21oi_1 _5689_ (.A1(_0748_),
    .A2(_0751_),
    .B1(_0747_),
    .Y(_3196_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_0740_),
    .B(_0744_),
    .Y(_3197_));
 sky130_fd_sc_hd__nor2_1 _5691_ (.A(_3196_),
    .B(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hd__a211oi_1 _5692_ (.A1(_0740_),
    .A2(_0743_),
    .B1(_3198_),
    .C1(_0739_),
    .Y(_3199_));
 sky130_fd_sc_hd__a21oi_1 _5693_ (.A1(_0772_),
    .A2(_0775_),
    .B1(_0771_),
    .Y(_3200_));
 sky130_fd_sc_hd__nor2b_1 _5694_ (.A(_3200_),
    .B_N(_0768_),
    .Y(_3201_));
 sky130_fd_sc_hd__a21oi_1 _5695_ (.A1(_0780_),
    .A2(_0783_),
    .B1(_0779_),
    .Y(_3202_));
 sky130_fd_sc_hd__nor2_1 _5696_ (.A(_0763_),
    .B(_0767_),
    .Y(_3203_));
 sky130_fd_sc_hd__o21ai_0 _5697_ (.A1(_3193_),
    .A2(_3202_),
    .B1(_3203_),
    .Y(_3204_));
 sky130_fd_sc_hd__o221ai_1 _5698_ (.A1(_0764_),
    .A2(_0763_),
    .B1(_3201_),
    .B2(_3204_),
    .C1(_3166_),
    .Y(_3205_));
 sky130_fd_sc_hd__a211oi_1 _5699_ (.A1(_0732_),
    .A2(_0735_),
    .B1(_0731_),
    .C1(_0727_),
    .Y(_3206_));
 sky130_fd_sc_hd__o21ai_0 _5700_ (.A1(_0728_),
    .A2(_0727_),
    .B1(_0724_),
    .Y(_3207_));
 sky130_fd_sc_hd__nor2_1 _5701_ (.A(_3206_),
    .B(_3207_),
    .Y(_3208_));
 sky130_fd_sc_hd__a21oi_1 _5702_ (.A1(_0756_),
    .A2(_0759_),
    .B1(_0755_),
    .Y(_3209_));
 sky130_fd_sc_hd__nor3_1 _5703_ (.A(_3163_),
    .B(_3164_),
    .C(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__nor3_1 _5704_ (.A(_0723_),
    .B(_3208_),
    .C(_3210_),
    .Y(_3211_));
 sky130_fd_sc_hd__o211ai_1 _5705_ (.A1(_3163_),
    .A2(_3199_),
    .B1(_3205_),
    .C1(_3211_),
    .Y(_3212_));
 sky130_fd_sc_hd__a41oi_1 _5706_ (.A1(_3166_),
    .A2(_3171_),
    .A3(_3192_),
    .A4(_3195_),
    .B1(_3212_),
    .Y(_3213_));
 sky130_fd_sc_hd__inv_1 _5707_ (.A(net556),
    .Y(_3214_));
 sky130_fd_sc_hd__nor2_1 _5708_ (.A(_3214_),
    .B(net400),
    .Y(_3215_));
 sky130_fd_sc_hd__a32oi_1 _5709_ (.A1(_3214_),
    .A2(net132),
    .A3(_1464_),
    .B1(_3215_),
    .B2(net565),
    .Y(_3216_));
 sky130_fd_sc_hd__o21ai_0 _5710_ (.A1(net555),
    .A2(_3216_),
    .B1(net545),
    .Y(_3217_));
 sky130_fd_sc_hd__o21ai_0 _5711_ (.A1(net1268),
    .A2(_3213_),
    .B1(_3217_),
    .Y(_3425_));
 sky130_fd_sc_hd__nand4_1 _5712_ (.A(_0849_),
    .B(_0861_),
    .C(_0857_),
    .D(_0853_),
    .Y(_3218_));
 sky130_fd_sc_hd__nand4_1 _5713_ (.A(_0865_),
    .B(_0877_),
    .C(_0873_),
    .D(_0869_),
    .Y(_3219_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(_0881_),
    .B(_0885_),
    .Y(_3220_));
 sky130_fd_sc_hd__nor3_1 _5715_ (.A(_3218_),
    .B(_3219_),
    .C(_3220_),
    .Y(_3221_));
 sky130_fd_sc_hd__o21ai_0 _5716_ (.A1(_0829_),
    .A2(_0828_),
    .B1(_0825_),
    .Y(_3222_));
 sky130_fd_sc_hd__nor2_1 _5717_ (.A(_0820_),
    .B(_0824_),
    .Y(_3223_));
 sky130_fd_sc_hd__o21ai_0 _5718_ (.A1(_0821_),
    .A2(_0820_),
    .B1(_0817_),
    .Y(_3224_));
 sky130_fd_sc_hd__a21oi_1 _5719_ (.A1(_3222_),
    .A2(_3223_),
    .B1(_3224_),
    .Y(_3225_));
 sky130_fd_sc_hd__or2_2 _5720_ (.A(_0816_),
    .B(_3225_),
    .X(_3226_));
 sky130_fd_sc_hd__nand4_1 _5721_ (.A(_0833_),
    .B(_0845_),
    .C(_0841_),
    .D(_0837_),
    .Y(_3227_));
 sky130_fd_sc_hd__nor2b_1 _5722_ (.A(_0786_),
    .B_N(_0785_),
    .Y(_3228_));
 sky130_fd_sc_hd__nand2_1 _5723_ (.A(_0789_),
    .B(_0797_),
    .Y(_3229_));
 sky130_fd_sc_hd__a211oi_1 _5724_ (.A1(_0797_),
    .A2(_0788_),
    .B1(_0792_),
    .C1(_0796_),
    .Y(_3230_));
 sky130_fd_sc_hd__o21ai_0 _5725_ (.A1(_3228_),
    .A2(_3229_),
    .B1(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__nand2_1 _5726_ (.A(_0801_),
    .B(_0805_),
    .Y(_3232_));
 sky130_fd_sc_hd__nand2_1 _5727_ (.A(_0813_),
    .B(_0809_),
    .Y(_3233_));
 sky130_fd_sc_hd__nor2_1 _5728_ (.A(_0793_),
    .B(_0792_),
    .Y(_3234_));
 sky130_fd_sc_hd__nor3_1 _5729_ (.A(_3232_),
    .B(_3233_),
    .C(_3234_),
    .Y(_3235_));
 sky130_fd_sc_hd__a21oi_1 _5730_ (.A1(_0809_),
    .A2(_0812_),
    .B1(_0808_),
    .Y(_3236_));
 sky130_fd_sc_hd__a21oi_1 _5731_ (.A1(_0801_),
    .A2(_0804_),
    .B1(_0800_),
    .Y(_3237_));
 sky130_fd_sc_hd__o21ai_0 _5732_ (.A1(_3236_),
    .A2(_3232_),
    .B1(_3237_),
    .Y(_3238_));
 sky130_fd_sc_hd__a21oi_1 _5733_ (.A1(_3231_),
    .A2(_3235_),
    .B1(_3238_),
    .Y(_3239_));
 sky130_fd_sc_hd__a21o_1 _5734_ (.A1(_0841_),
    .A2(_0844_),
    .B1(_0840_),
    .X(_3240_));
 sky130_fd_sc_hd__a21o_1 _5735_ (.A1(_0837_),
    .A2(_3240_),
    .B1(_0836_),
    .X(_3241_));
 sky130_fd_sc_hd__a21oi_1 _5736_ (.A1(_0825_),
    .A2(_0828_),
    .B1(_0824_),
    .Y(_3242_));
 sky130_fd_sc_hd__nand2_1 _5737_ (.A(_0817_),
    .B(_0821_),
    .Y(_3243_));
 sky130_fd_sc_hd__a211oi_1 _5738_ (.A1(_0817_),
    .A2(_0820_),
    .B1(_0832_),
    .C1(_0816_),
    .Y(_3244_));
 sky130_fd_sc_hd__o21ai_0 _5739_ (.A1(_3242_),
    .A2(_3243_),
    .B1(_3244_),
    .Y(_3245_));
 sky130_fd_sc_hd__a21oi_1 _5740_ (.A1(_0833_),
    .A2(_3241_),
    .B1(_3245_),
    .Y(_3246_));
 sky130_fd_sc_hd__o21ai_0 _5741_ (.A1(_3227_),
    .A2(_3239_),
    .B1(_3246_),
    .Y(_3247_));
 sky130_fd_sc_hd__nand3_1 _5742_ (.A(_0893_),
    .B(_0897_),
    .C(_0901_),
    .Y(_3248_));
 sky130_fd_sc_hd__nand3_1 _5743_ (.A(_0889_),
    .B(_0909_),
    .C(_0905_),
    .Y(_3249_));
 sky130_fd_sc_hd__nor2_1 _5744_ (.A(_3248_),
    .B(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__a21oi_1 _5745_ (.A1(_0873_),
    .A2(_0876_),
    .B1(_0872_),
    .Y(_3251_));
 sky130_fd_sc_hd__nand2_1 _5746_ (.A(_0865_),
    .B(_0869_),
    .Y(_3252_));
 sky130_fd_sc_hd__nor2_1 _5747_ (.A(_3251_),
    .B(_3252_),
    .Y(_3253_));
 sky130_fd_sc_hd__a211oi_1 _5748_ (.A1(_0865_),
    .A2(_0868_),
    .B1(_3253_),
    .C1(_0864_),
    .Y(_3254_));
 sky130_fd_sc_hd__a211oi_1 _5749_ (.A1(_0857_),
    .A2(_0860_),
    .B1(_0856_),
    .C1(_0852_),
    .Y(_3255_));
 sky130_fd_sc_hd__o21ai_0 _5750_ (.A1(_0853_),
    .A2(_0852_),
    .B1(_0849_),
    .Y(_3256_));
 sky130_fd_sc_hd__nor2_1 _5751_ (.A(_3255_),
    .B(_3256_),
    .Y(_3257_));
 sky130_fd_sc_hd__a21oi_1 _5752_ (.A1(_0881_),
    .A2(_0884_),
    .B1(_0880_),
    .Y(_3258_));
 sky130_fd_sc_hd__nor3_1 _5753_ (.A(_3218_),
    .B(_3219_),
    .C(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__nor3_1 _5754_ (.A(_0848_),
    .B(_3257_),
    .C(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__a21oi_1 _5755_ (.A1(_0897_),
    .A2(_0900_),
    .B1(_0896_),
    .Y(_3261_));
 sky130_fd_sc_hd__nor2b_1 _5756_ (.A(_3261_),
    .B_N(_0893_),
    .Y(_3262_));
 sky130_fd_sc_hd__a21oi_1 _5757_ (.A1(_0905_),
    .A2(_0908_),
    .B1(_0904_),
    .Y(_3263_));
 sky130_fd_sc_hd__nor2_1 _5758_ (.A(_0888_),
    .B(_0892_),
    .Y(_3264_));
 sky130_fd_sc_hd__o21ai_0 _5759_ (.A1(_3248_),
    .A2(_3263_),
    .B1(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__o221ai_1 _5760_ (.A1(_0889_),
    .A2(_0888_),
    .B1(_3262_),
    .B2(_3265_),
    .C1(_3221_),
    .Y(_3266_));
 sky130_fd_sc_hd__o211ai_1 _5761_ (.A1(_3218_),
    .A2(_3254_),
    .B1(_3260_),
    .C1(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__a41oi_1 _5762_ (.A1(_3221_),
    .A2(_3226_),
    .A3(_3247_),
    .A4(_3250_),
    .B1(_3267_),
    .Y(_3268_));
 sky130_fd_sc_hd__inv_1 _5763_ (.A(net564),
    .Y(_3269_));
 sky130_fd_sc_hd__nor2_1 _5764_ (.A(_3269_),
    .B(net399),
    .Y(_3270_));
 sky130_fd_sc_hd__a32oi_1 _5765_ (.A1(_3269_),
    .A2(net131),
    .A3(_1603_),
    .B1(_3270_),
    .B2(net562),
    .Y(_3271_));
 sky130_fd_sc_hd__o21ai_0 _5766_ (.A1(net563),
    .A2(_3271_),
    .B1(net544),
    .Y(_3272_));
 sky130_fd_sc_hd__o21ai_0 _5767_ (.A1(net1266),
    .A2(net1227),
    .B1(_3272_),
    .Y(_3423_));
 sky130_fd_sc_hd__nor2_1 _5768_ (.A(_3214_),
    .B(net555),
    .Y(_3273_));
 sky130_fd_sc_hd__nor4bb_4 _5769_ (.A(net556),
    .B(net565),
    .C_N(net537),
    .D_N(net555),
    .Y(_3274_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input52 (.A(net1615),
    .X(net52));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input51 (.A(net1606),
    .X(net51));
 sky130_fd_sc_hd__a311o_1 _5772_ (.A1(net565),
    .A2(net400),
    .A3(_3273_),
    .B1(_2513_),
    .C1(net1262),
    .X(_3431_));
 sky130_fd_sc_hd__a22o_1 _5773_ (.A1(net555),
    .A2(_1464_),
    .B1(_3042_),
    .B2(_3214_),
    .X(_3432_));
 sky130_fd_sc_hd__or3_1 _5774_ (.A(_3214_),
    .B(net555),
    .C(net565),
    .X(_3277_));
 sky130_fd_sc_hd__nand2_1 _5775_ (.A(net565),
    .B(net400),
    .Y(_3278_));
 sky130_fd_sc_hd__o21ai_0 _5776_ (.A1(net565),
    .A2(net404),
    .B1(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__mux2_2 _5777_ (.A0(net565),
    .A1(_1464_),
    .S(net556),
    .X(_3280_));
 sky130_fd_sc_hd__a22oi_1 _5778_ (.A1(_3273_),
    .A2(_3279_),
    .B1(_3280_),
    .B2(net555),
    .Y(_3281_));
 sky130_fd_sc_hd__o21ai_0 _5779_ (.A1(_3213_),
    .A2(_3277_),
    .B1(_3281_),
    .Y(_3433_));
 sky130_fd_sc_hd__nor2_1 _5780_ (.A(_3269_),
    .B(net563),
    .Y(_3282_));
 sky130_fd_sc_hd__nor4bb_4 _5781_ (.A(net564),
    .B(net562),
    .C_N(net536),
    .D_N(net563),
    .Y(_3283_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input50 (.A(net1585),
    .X(net50));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input49 (.A(net1621),
    .X(net49));
 sky130_fd_sc_hd__a31oi_1 _5784_ (.A1(net562),
    .A2(net399),
    .A3(_3282_),
    .B1(_3283_),
    .Y(_3286_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(_2610_),
    .B(_3286_),
    .Y(_3434_));
 sky130_fd_sc_hd__a22o_1 _5786_ (.A1(net563),
    .A2(_1603_),
    .B1(_3047_),
    .B2(_3269_),
    .X(_3435_));
 sky130_fd_sc_hd__or3_1 _5787_ (.A(_3269_),
    .B(net563),
    .C(net562),
    .X(_3287_));
 sky130_fd_sc_hd__nand2_1 _5788_ (.A(net562),
    .B(net399),
    .Y(_3288_));
 sky130_fd_sc_hd__o21ai_0 _5789_ (.A1(net562),
    .A2(net403),
    .B1(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__mux2_2 _5790_ (.A0(net562),
    .A1(_1603_),
    .S(net564),
    .X(_3290_));
 sky130_fd_sc_hd__a22oi_1 _5791_ (.A1(_3282_),
    .A2(_3289_),
    .B1(_3290_),
    .B2(net563),
    .Y(_3291_));
 sky130_fd_sc_hd__o21ai_0 _5792_ (.A1(net1227),
    .A2(_3287_),
    .B1(_3291_),
    .Y(_3436_));
 sky130_fd_sc_hd__and3_2 _5793_ (.A(net1272),
    .B(net535),
    .C(_1732_),
    .X(_3292_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input48 (.A(net1577),
    .X(net48));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input47 (.A(net1578),
    .X(net47));
 sky130_fd_sc_hd__a31oi_1 _5796_ (.A1(net1271),
    .A2(net1273),
    .A3(_1731_),
    .B1(net1238),
    .Y(_3295_));
 sky130_fd_sc_hd__nand2_1 _5797_ (.A(net1232),
    .B(_3295_),
    .Y(_3437_));
 sky130_fd_sc_hd__nand2b_1 _5798_ (.A_N(net1271),
    .B(_3037_),
    .Y(_3296_));
 sky130_fd_sc_hd__nand3b_1 _5799_ (.A_N(net1273),
    .B(net1272),
    .C(net398),
    .Y(_3297_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(_3296_),
    .B(_3297_),
    .Y(_3438_));
 sky130_fd_sc_hd__nand3b_1 _5801_ (.A_N(net1271),
    .B(net1273),
    .C(net1272),
    .Y(_3298_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input46 (.A(net1569),
    .X(net46));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input45 (.A(net1623),
    .X(net45));
 sky130_fd_sc_hd__inv_1 _5804_ (.A(net1272),
    .Y(_3301_));
 sky130_fd_sc_hd__nor2_1 _5805_ (.A(_3301_),
    .B(net398),
    .Y(_3302_));
 sky130_fd_sc_hd__nor2_1 _5806_ (.A(net1273),
    .B(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__o21ai_0 _5807_ (.A1(_1731_),
    .A2(_3303_),
    .B1(net1271),
    .Y(_3304_));
 sky130_fd_sc_hd__a21oi_1 _5808_ (.A1(_3301_),
    .A2(net1293),
    .B1(_3302_),
    .Y(_3305_));
 sky130_fd_sc_hd__a2111oi_0 _5809_ (.A1(net1271),
    .A2(_3305_),
    .B1(_3161_),
    .C1(_3134_),
    .D1(net1273),
    .Y(_3306_));
 sky130_fd_sc_hd__a21oi_1 _5810_ (.A1(net1258),
    .A2(_3304_),
    .B1(_3306_),
    .Y(_3439_));
 sky130_fd_sc_hd__and3_1 _5811_ (.A(net557),
    .B(net534),
    .C(_1865_),
    .X(_3307_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input44 (.A(net1553),
    .X(net44));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input43 (.A(channel_dst_addr[22]),
    .X(net43));
 sky130_fd_sc_hd__a31oi_1 _5814_ (.A1(net558),
    .A2(net554),
    .A3(_1864_),
    .B1(_3307_),
    .Y(_3310_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(_2896_),
    .B(_3310_),
    .Y(_3440_));
 sky130_fd_sc_hd__nand2b_1 _5816_ (.A_N(net558),
    .B(_3033_),
    .Y(_3311_));
 sky130_fd_sc_hd__inv_1 _5817_ (.A(net554),
    .Y(_3312_));
 sky130_fd_sc_hd__nand3_1 _5818_ (.A(_3312_),
    .B(net557),
    .C(net397),
    .Y(_3313_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_3311_),
    .B(_3313_),
    .Y(_3441_));
 sky130_fd_sc_hd__nand2_1 _5820_ (.A(net558),
    .B(_3312_),
    .Y(_3314_));
 sky130_fd_sc_hd__nor2_1 _5821_ (.A(net557),
    .B(net401),
    .Y(_3315_));
 sky130_fd_sc_hd__a21oi_1 _5822_ (.A1(net557),
    .A2(net397),
    .B1(_3315_),
    .Y(_3316_));
 sky130_fd_sc_hd__mux2i_1 _5823_ (.A0(net557),
    .A1(_1864_),
    .S(net558),
    .Y(_3317_));
 sky130_fd_sc_hd__o22ai_1 _5824_ (.A1(_3314_),
    .A2(_3316_),
    .B1(_3317_),
    .B2(_3312_),
    .Y(_3318_));
 sky130_fd_sc_hd__nor2_1 _5825_ (.A(net557),
    .B(_3314_),
    .Y(_3319_));
 sky130_fd_sc_hd__nor3_1 _5826_ (.A(_3102_),
    .B(_3106_),
    .C(_3318_),
    .Y(_3320_));
 sky130_fd_sc_hd__a2bb2oi_1 _5827_ (.A1_N(_3318_),
    .A2_N(_3319_),
    .B1(_3320_),
    .B2(_3081_),
    .Y(_3442_));
 sky130_fd_sc_hd__a32oi_1 _5828_ (.A1(net400),
    .A2(net132),
    .A3(_1453_),
    .B1(_3215_),
    .B2(net555),
    .Y(_3321_));
 sky130_fd_sc_hd__o21a_1 _5829_ (.A1(net565),
    .A2(_3321_),
    .B1(net549),
    .X(_0011_));
 sky130_fd_sc_hd__a32oi_1 _5830_ (.A1(net399),
    .A2(net131),
    .A3(_1450_),
    .B1(_3270_),
    .B2(net563),
    .Y(_3322_));
 sky130_fd_sc_hd__o21a_1 _5831_ (.A1(net562),
    .A2(_3322_),
    .B1(net548),
    .X(_0010_));
 sky130_fd_sc_hd__o22a_1 _5832_ (.A1(net540),
    .A2(_1604_),
    .B1(net1266),
    .B2(net1227),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _5833_ (.A(net130),
    .B(_1731_),
    .Y(_3323_));
 sky130_fd_sc_hd__nor2_1 _5834_ (.A(net1271),
    .B(_3323_),
    .Y(_3324_));
 sky130_fd_sc_hd__a21oi_1 _5835_ (.A1(net1271),
    .A2(_3302_),
    .B1(_3324_),
    .Y(_3325_));
 sky130_fd_sc_hd__o21a_1 _5836_ (.A1(net1273),
    .A2(_3325_),
    .B1(net547),
    .X(_0009_));
 sky130_fd_sc_hd__o21a_1 _5837_ (.A1(net539),
    .A2(_1733_),
    .B1(_3162_),
    .X(_0005_));
 sky130_fd_sc_hd__o22a_1 _5838_ (.A1(net541),
    .A2(net1251),
    .B1(net1268),
    .B2(_3213_),
    .X(_0007_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(net129),
    .B(_1864_),
    .Y(_3326_));
 sky130_fd_sc_hd__nor2_1 _5840_ (.A(net558),
    .B(_3326_),
    .Y(_3327_));
 sky130_fd_sc_hd__a31oi_1 _5841_ (.A1(net558),
    .A2(net557),
    .A3(_3082_),
    .B1(_3327_),
    .Y(_3328_));
 sky130_fd_sc_hd__o21a_1 _5842_ (.A1(net554),
    .A2(_3328_),
    .B1(net546),
    .X(_0008_));
 sky130_fd_sc_hd__nor2_1 _5843_ (.A(net538),
    .B(_1866_),
    .Y(_3329_));
 sky130_fd_sc_hd__nor3_1 _5844_ (.A(_3102_),
    .B(_3106_),
    .C(_3329_),
    .Y(_3330_));
 sky130_fd_sc_hd__o2bb2ai_1 _5845_ (.A1_N(_3081_),
    .A2_N(_3330_),
    .B1(_3329_),
    .B2(net1263),
    .Y(_0004_));
 sky130_fd_sc_hd__nor2_1 _5846_ (.A(\active_channel_count[2] ),
    .B(\active_channel_count[3] ),
    .Y(_3331_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_0407_),
    .B(_3331_),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_1 _5848_ (.A(net185),
    .Y(_0410_));
 sky130_fd_sc_hd__inv_1 _5849_ (.A(net184),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_1 _5850_ (.A(net182),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_1 _5851_ (.A(net181),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_1 _5852_ (.A(net180),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_1 _5853_ (.A(net179),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_1 _5854_ (.A(net178),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_1 _5855_ (.A(net177),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_1 _5856_ (.A(net176),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_1 _5857_ (.A(net175),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_1 _5858_ (.A(net174),
    .Y(_0450_));
 sky130_fd_sc_hd__inv_1 _5859_ (.A(net173),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_1 _5860_ (.A(net171),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_1 _5861_ (.A(net170),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_1 _5862_ (.A(net169),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_1 _5863_ (.A(net168),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_1 _5864_ (.A(net167),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_1 _5865_ (.A(net166),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_1 _5866_ (.A(net165),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_1 _5867_ (.A(net164),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_1 _5868_ (.A(net155),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_1 _5869_ (.A(net144),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_1 _5870_ (.A(net260),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_1 _5871_ (.A(net249),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_1 _5872_ (.A(net227),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_1 _5873_ (.A(net216),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_1 _5874_ (.A(net205),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_1 _5875_ (.A(net194),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_1 _5876_ (.A(net183),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_1 _5877_ (.A(net172),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_1 _5878_ (.A(net187),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_1 _5879_ (.A(net189),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_1 _5880_ (.A(net188),
    .Y(_0544_));
 sky130_fd_sc_hd__inv_1 _5881_ (.A(net193),
    .Y(_0548_));
 sky130_fd_sc_hd__inv_1 _5882_ (.A(net192),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_1 _5883_ (.A(net191),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_1 _5884_ (.A(net190),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_1 _5885_ (.A(net202),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_1 _5886_ (.A(net201),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_1 _5887_ (.A(net200),
    .Y(_0572_));
 sky130_fd_sc_hd__inv_1 _5888_ (.A(net199),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_1 _5889_ (.A(net198),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_1 _5890_ (.A(net197),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_1 _5891_ (.A(net196),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_1 _5892_ (.A(net195),
    .Y(_0592_));
 sky130_fd_sc_hd__inv_1 _5893_ (.A(net220),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_1 _5894_ (.A(net218),
    .Y(_0604_));
 sky130_fd_sc_hd__inv_1 _5895_ (.A(net217),
    .Y(_0608_));
 sky130_fd_sc_hd__inv_1 _5896_ (.A(net215),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_1 _5897_ (.A(net214),
    .Y(_0616_));
 sky130_fd_sc_hd__inv_1 _5898_ (.A(net213),
    .Y(_0620_));
 sky130_fd_sc_hd__inv_1 _5899_ (.A(net210),
    .Y(_0632_));
 sky130_fd_sc_hd__inv_1 _5900_ (.A(net209),
    .Y(_0636_));
 sky130_fd_sc_hd__inv_1 _5901_ (.A(net208),
    .Y(_0640_));
 sky130_fd_sc_hd__inv_1 _5902_ (.A(net207),
    .Y(_0644_));
 sky130_fd_sc_hd__inv_1 _5903_ (.A(net206),
    .Y(_0648_));
 sky130_fd_sc_hd__inv_1 _5904_ (.A(net204),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_1 _5905_ (.A(net203),
    .Y(_0656_));
 sky130_fd_sc_hd__inv_1 _5906_ (.A(net257),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_1 _5907_ (.A(net259),
    .Y(_0665_));
 sky130_fd_sc_hd__inv_1 _5908_ (.A(net258),
    .Y(_0669_));
 sky130_fd_sc_hd__inv_1 _5909_ (.A(net137),
    .Y(_0673_));
 sky130_fd_sc_hd__inv_1 _5910_ (.A(net136),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_1 _5911_ (.A(net135),
    .Y(_0681_));
 sky130_fd_sc_hd__inv_1 _5912_ (.A(net134),
    .Y(_0685_));
 sky130_fd_sc_hd__inv_1 _5913_ (.A(net146),
    .Y(_0689_));
 sky130_fd_sc_hd__inv_1 _5914_ (.A(net145),
    .Y(_0693_));
 sky130_fd_sc_hd__inv_1 _5915_ (.A(net143),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_1 _5916_ (.A(net142),
    .Y(_0701_));
 sky130_fd_sc_hd__inv_1 _5917_ (.A(net141),
    .Y(_0705_));
 sky130_fd_sc_hd__inv_1 _5918_ (.A(net140),
    .Y(_0709_));
 sky130_fd_sc_hd__inv_1 _5919_ (.A(net139),
    .Y(_0713_));
 sky130_fd_sc_hd__inv_1 _5920_ (.A(net138),
    .Y(_0717_));
 sky130_fd_sc_hd__inv_1 _5921_ (.A(net163),
    .Y(_0721_));
 sky130_fd_sc_hd__inv_1 _5922_ (.A(net162),
    .Y(_0725_));
 sky130_fd_sc_hd__inv_1 _5923_ (.A(net161),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_1 _5924_ (.A(net160),
    .Y(_0733_));
 sky130_fd_sc_hd__inv_1 _5925_ (.A(net159),
    .Y(_0737_));
 sky130_fd_sc_hd__inv_1 _5926_ (.A(net158),
    .Y(_0741_));
 sky130_fd_sc_hd__inv_1 _5927_ (.A(net157),
    .Y(_0745_));
 sky130_fd_sc_hd__inv_1 _5928_ (.A(net156),
    .Y(_0749_));
 sky130_fd_sc_hd__inv_1 _5929_ (.A(net154),
    .Y(_0753_));
 sky130_fd_sc_hd__inv_1 _5930_ (.A(net153),
    .Y(_0757_));
 sky130_fd_sc_hd__inv_1 _5931_ (.A(net152),
    .Y(_0761_));
 sky130_fd_sc_hd__inv_1 _5932_ (.A(net151),
    .Y(_0765_));
 sky130_fd_sc_hd__inv_1 _5933_ (.A(net150),
    .Y(_0769_));
 sky130_fd_sc_hd__inv_1 _5934_ (.A(net149),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_1 _5935_ (.A(net148),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_1 _5936_ (.A(net147),
    .Y(_0781_));
 sky130_fd_sc_hd__inv_1 _5937_ (.A(net222),
    .Y(_0787_));
 sky130_fd_sc_hd__inv_1 _5938_ (.A(net224),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_1 _5939_ (.A(net223),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_1 _5940_ (.A(net229),
    .Y(_0798_));
 sky130_fd_sc_hd__inv_1 _5941_ (.A(net228),
    .Y(_0802_));
 sky130_fd_sc_hd__inv_1 _5942_ (.A(net226),
    .Y(_0806_));
 sky130_fd_sc_hd__inv_1 _5943_ (.A(net225),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_1 _5944_ (.A(net237),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_1 _5945_ (.A(net236),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_1 _5946_ (.A(net235),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_1 _5947_ (.A(net234),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_1 _5948_ (.A(net233),
    .Y(_0830_));
 sky130_fd_sc_hd__inv_1 _5949_ (.A(net232),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_1 _5950_ (.A(net231),
    .Y(_0838_));
 sky130_fd_sc_hd__inv_1 _5951_ (.A(net230),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_1 _5952_ (.A(net255),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_1 _5953_ (.A(net254),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_1 _5954_ (.A(net253),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_1 _5955_ (.A(net252),
    .Y(_0858_));
 sky130_fd_sc_hd__inv_1 _5956_ (.A(net251),
    .Y(_0862_));
 sky130_fd_sc_hd__inv_1 _5957_ (.A(net250),
    .Y(_0866_));
 sky130_fd_sc_hd__inv_1 _5958_ (.A(net248),
    .Y(_0870_));
 sky130_fd_sc_hd__inv_1 _5959_ (.A(net247),
    .Y(_0874_));
 sky130_fd_sc_hd__inv_1 _5960_ (.A(net246),
    .Y(_0878_));
 sky130_fd_sc_hd__inv_1 _5961_ (.A(net245),
    .Y(_0882_));
 sky130_fd_sc_hd__inv_1 _5962_ (.A(net244),
    .Y(_0886_));
 sky130_fd_sc_hd__inv_1 _5963_ (.A(net243),
    .Y(_0890_));
 sky130_fd_sc_hd__inv_1 _5964_ (.A(net242),
    .Y(_0894_));
 sky130_fd_sc_hd__inv_1 _5965_ (.A(net241),
    .Y(_0898_));
 sky130_fd_sc_hd__inv_1 _5966_ (.A(net240),
    .Y(_0902_));
 sky130_fd_sc_hd__inv_1 _5967_ (.A(net239),
    .Y(_0906_));
 sky130_fd_sc_hd__inv_1 _5968_ (.A(\active_channel_count[1] ),
    .Y(_0406_));
 sky130_fd_sc_hd__inv_1 _5969_ (.A(net238),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_1 _5970_ (.A(net219),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_1 _5971_ (.A(net212),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_1 _5972_ (.A(net211),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _5973_ (.A(net1),
    .B(_1866_),
    .Y(_3332_));
 sky130_fd_sc_hd__nand2_1 _5974_ (.A(\current_dst_addr[0][0] ),
    .B(_1880_),
    .Y(_3333_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_3332_),
    .B(_3333_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2_1 _5976_ (.A(net40),
    .B(_1866_),
    .Y(_3334_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(\current_dst_addr[0][1] ),
    .B(_1880_),
    .Y(_3335_));
 sky130_fd_sc_hd__nand2_1 _5978_ (.A(_3334_),
    .B(_3335_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _5979_ (.A(net54),
    .B(_1733_),
    .Y(_3336_));
 sky130_fd_sc_hd__nand2_1 _5980_ (.A(\current_dst_addr[1][0] ),
    .B(_1748_),
    .Y(_3337_));
 sky130_fd_sc_hd__nand2_1 _5981_ (.A(_3336_),
    .B(_3337_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(net55),
    .B(_1733_),
    .Y(_3338_));
 sky130_fd_sc_hd__nand2_1 _5983_ (.A(\current_dst_addr[1][1] ),
    .B(_1748_),
    .Y(_3339_));
 sky130_fd_sc_hd__nand2_1 _5984_ (.A(_3338_),
    .B(_3339_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(net89),
    .B(_1604_),
    .Y(_3340_));
 sky130_fd_sc_hd__nand2_1 _5986_ (.A(\current_dst_addr[2][0] ),
    .B(net1248),
    .Y(_3341_));
 sky130_fd_sc_hd__nand2_1 _5987_ (.A(_3340_),
    .B(_3341_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _5988_ (.A(net90),
    .B(net1249),
    .Y(_3342_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(\current_dst_addr[2][1] ),
    .B(net1248),
    .Y(_3343_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(_3342_),
    .B(_3343_),
    .Y(_0915_));
 sky130_fd_sc_hd__nand2_1 _5991_ (.A(net124),
    .B(net1251),
    .Y(_3344_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(\current_dst_addr[3][0] ),
    .B(net1250),
    .Y(_3345_));
 sky130_fd_sc_hd__nand2_1 _5993_ (.A(_3344_),
    .B(_3345_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _5994_ (.A(net125),
    .B(net1251),
    .Y(_3346_));
 sky130_fd_sc_hd__nand2_1 _5995_ (.A(\current_dst_addr[3][1] ),
    .B(net1250),
    .Y(_3347_));
 sky130_fd_sc_hd__nand2_1 _5996_ (.A(_3346_),
    .B(_3347_),
    .Y(_0917_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(net269),
    .B(_1866_),
    .Y(_3348_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(\current_src_addr[0][0] ),
    .B(net1243),
    .Y(_3349_));
 sky130_fd_sc_hd__nand2_1 _5999_ (.A(_3348_),
    .B(_3349_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _6000_ (.A(net308),
    .B(_1866_),
    .Y(_3350_));
 sky130_fd_sc_hd__nand2_1 _6001_ (.A(\current_src_addr[0][1] ),
    .B(net1243),
    .Y(_3351_));
 sky130_fd_sc_hd__nand2_1 _6002_ (.A(_3350_),
    .B(_3351_),
    .Y(_0919_));
 sky130_fd_sc_hd__nand2_1 _6003_ (.A(net322),
    .B(net1247),
    .Y(_3352_));
 sky130_fd_sc_hd__nand2_1 _6004_ (.A(\current_src_addr[1][0] ),
    .B(net1245),
    .Y(_3353_));
 sky130_fd_sc_hd__nand2_1 _6005_ (.A(_3352_),
    .B(_3353_),
    .Y(_0920_));
 sky130_fd_sc_hd__nand2_1 _6006_ (.A(net323),
    .B(net1247),
    .Y(_3354_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(\current_src_addr[1][1] ),
    .B(net1245),
    .Y(_3355_));
 sky130_fd_sc_hd__nand2_1 _6008_ (.A(_3354_),
    .B(_3355_),
    .Y(_0921_));
 sky130_fd_sc_hd__nand2_1 _6009_ (.A(net357),
    .B(_1604_),
    .Y(_3356_));
 sky130_fd_sc_hd__nand2_1 _6010_ (.A(\current_src_addr[2][0] ),
    .B(net1248),
    .Y(_3357_));
 sky130_fd_sc_hd__nand2_1 _6011_ (.A(_3356_),
    .B(_3357_),
    .Y(_0922_));
 sky130_fd_sc_hd__nand2_1 _6012_ (.A(net358),
    .B(net1249),
    .Y(_3358_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(\current_src_addr[2][1] ),
    .B(net1248),
    .Y(_3359_));
 sky130_fd_sc_hd__nand2_1 _6014_ (.A(_3358_),
    .B(_3359_),
    .Y(_0923_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(net392),
    .B(net1251),
    .Y(_3360_));
 sky130_fd_sc_hd__nand2_1 _6016_ (.A(\current_src_addr[3][0] ),
    .B(net1250),
    .Y(_3361_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(_3360_),
    .B(_3361_),
    .Y(_0924_));
 sky130_fd_sc_hd__nand2_1 _6018_ (.A(net393),
    .B(net1251),
    .Y(_3362_));
 sky130_fd_sc_hd__nand2_1 _6019_ (.A(\current_src_addr[3][1] ),
    .B(net1250),
    .Y(_3363_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_3362_),
    .B(_3363_),
    .Y(_0925_));
 sky130_fd_sc_hd__mux2_2 _6021_ (.A0(\data_buffer[0][0] ),
    .A1(net406),
    .S(net1237),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_2 _6022_ (.A0(\data_buffer[0][10] ),
    .A1(net417),
    .S(net1237),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_2 _6023_ (.A0(\data_buffer[0][11] ),
    .A1(net428),
    .S(net1237),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_2 _6024_ (.A0(\data_buffer[0][12] ),
    .A1(net437),
    .S(net1237),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_2 _6025_ (.A0(\data_buffer[0][13] ),
    .A1(net438),
    .S(net1237),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_2 _6026_ (.A0(\data_buffer[0][14] ),
    .A1(net439),
    .S(net1237),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_2 _6027_ (.A0(\data_buffer[0][15] ),
    .A1(net440),
    .S(net1237),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_2 _6028_ (.A0(\data_buffer[0][16] ),
    .A1(net441),
    .S(net1237),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_2 _6029_ (.A0(\data_buffer[0][17] ),
    .A1(net442),
    .S(net1237),
    .X(_0934_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input42 (.A(net1539),
    .X(net42));
 sky130_fd_sc_hd__mux2_2 _6031_ (.A0(\data_buffer[0][18] ),
    .A1(net443),
    .S(net1237),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_2 _6032_ (.A0(\data_buffer[0][19] ),
    .A1(net444),
    .S(net1237),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_2 _6033_ (.A0(\data_buffer[0][1] ),
    .A1(net445),
    .S(net1237),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_2 _6034_ (.A0(\data_buffer[0][20] ),
    .A1(net446),
    .S(net1237),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_2 _6035_ (.A0(\data_buffer[0][21] ),
    .A1(net447),
    .S(net1237),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_2 _6036_ (.A0(\data_buffer[0][22] ),
    .A1(net448),
    .S(net1237),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_2 _6037_ (.A0(\data_buffer[0][23] ),
    .A1(net449),
    .S(net1237),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_2 _6038_ (.A0(\data_buffer[0][24] ),
    .A1(net450),
    .S(net1237),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_2 _6039_ (.A0(\data_buffer[0][25] ),
    .A1(net451),
    .S(net1237),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_2 _6040_ (.A0(\data_buffer[0][26] ),
    .A1(net452),
    .S(net1237),
    .X(_0944_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input41 (.A(net1579),
    .X(net41));
 sky130_fd_sc_hd__mux2_2 _6042_ (.A0(\data_buffer[0][27] ),
    .A1(net453),
    .S(net1237),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_2 _6043_ (.A0(\data_buffer[0][28] ),
    .A1(net454),
    .S(net1237),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_2 _6044_ (.A0(\data_buffer[0][29] ),
    .A1(net455),
    .S(net1237),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_2 _6045_ (.A0(\data_buffer[0][2] ),
    .A1(net456),
    .S(net1237),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_2 _6046_ (.A0(\data_buffer[0][30] ),
    .A1(net457),
    .S(net1237),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_2 _6047_ (.A0(\data_buffer[0][31] ),
    .A1(net458),
    .S(net1237),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_2 _6048_ (.A0(\data_buffer[0][3] ),
    .A1(net467),
    .S(net1237),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_2 _6049_ (.A0(\data_buffer[0][4] ),
    .A1(net478),
    .S(net1237),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_2 _6050_ (.A0(\data_buffer[0][5] ),
    .A1(net489),
    .S(net1237),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_2 _6051_ (.A0(\data_buffer[0][6] ),
    .A1(net500),
    .S(net1237),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_2 _6052_ (.A0(\data_buffer[0][7] ),
    .A1(net511),
    .S(net1237),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_2 _6053_ (.A0(\data_buffer[0][8] ),
    .A1(net522),
    .S(net1237),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_2 _6054_ (.A0(\data_buffer[0][9] ),
    .A1(net533),
    .S(net1237),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_2 _6055_ (.A0(\data_buffer[1][0] ),
    .A1(net459),
    .S(net1238),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_2 _6056_ (.A0(\data_buffer[1][10] ),
    .A1(net470),
    .S(net1238),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_2 _6057_ (.A0(\data_buffer[1][11] ),
    .A1(net471),
    .S(net1238),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_2 _6058_ (.A0(\data_buffer[1][12] ),
    .A1(net472),
    .S(net1238),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_2 _6059_ (.A0(\data_buffer[1][13] ),
    .A1(net473),
    .S(net1238),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_2 _6060_ (.A0(\data_buffer[1][14] ),
    .A1(net474),
    .S(net1238),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_2 _6061_ (.A0(\data_buffer[1][15] ),
    .A1(net475),
    .S(net1238),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_2 _6062_ (.A0(\data_buffer[1][16] ),
    .A1(net476),
    .S(net1238),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_2 _6063_ (.A0(\data_buffer[1][17] ),
    .A1(net477),
    .S(net1238),
    .X(_0966_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input40 (.A(net1467),
    .X(net40));
 sky130_fd_sc_hd__mux2_2 _6065_ (.A0(\data_buffer[1][18] ),
    .A1(net479),
    .S(net1238),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_2 _6066_ (.A0(\data_buffer[1][19] ),
    .A1(net480),
    .S(net1238),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_2 _6067_ (.A0(\data_buffer[1][1] ),
    .A1(net460),
    .S(net1238),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_2 _6068_ (.A0(\data_buffer[1][20] ),
    .A1(net481),
    .S(net1238),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_2 _6069_ (.A0(\data_buffer[1][21] ),
    .A1(net482),
    .S(net1238),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_2 _6070_ (.A0(\data_buffer[1][22] ),
    .A1(net483),
    .S(net1238),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_2 _6071_ (.A0(\data_buffer[1][23] ),
    .A1(net484),
    .S(net1238),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_2 _6072_ (.A0(\data_buffer[1][24] ),
    .A1(net485),
    .S(net1238),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_2 _6073_ (.A0(\data_buffer[1][25] ),
    .A1(net486),
    .S(net1238),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_2 _6074_ (.A0(\data_buffer[1][26] ),
    .A1(net487),
    .S(net1238),
    .X(_0976_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input39 (.A(channel_dst_addr[19]),
    .X(net39));
 sky130_fd_sc_hd__mux2_2 _6076_ (.A0(\data_buffer[1][27] ),
    .A1(net488),
    .S(net1238),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_2 _6077_ (.A0(\data_buffer[1][28] ),
    .A1(net490),
    .S(net1238),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_2 _6078_ (.A0(\data_buffer[1][29] ),
    .A1(net491),
    .S(net1238),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_2 _6079_ (.A0(\data_buffer[1][2] ),
    .A1(net461),
    .S(net1238),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_2 _6080_ (.A0(\data_buffer[1][30] ),
    .A1(net492),
    .S(net1238),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_2 _6081_ (.A0(\data_buffer[1][31] ),
    .A1(net493),
    .S(net1238),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_2 _6082_ (.A0(\data_buffer[1][3] ),
    .A1(net462),
    .S(net1238),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_2 _6083_ (.A0(\data_buffer[1][4] ),
    .A1(net463),
    .S(net1238),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_2 _6084_ (.A0(\data_buffer[1][5] ),
    .A1(net464),
    .S(net1238),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_2 _6085_ (.A0(\data_buffer[1][6] ),
    .A1(net465),
    .S(net1238),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_2 _6086_ (.A0(\data_buffer[1][7] ),
    .A1(net466),
    .S(net1238),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_2 _6087_ (.A0(\data_buffer[1][8] ),
    .A1(net468),
    .S(net1238),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_2 _6088_ (.A0(\data_buffer[1][9] ),
    .A1(net469),
    .S(net1238),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_2 _6089_ (.A0(\data_buffer[2][0] ),
    .A1(net494),
    .S(net1260),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_2 _6090_ (.A0(\data_buffer[2][10] ),
    .A1(net505),
    .S(net1260),
    .X(_0991_));
 sky130_fd_sc_hd__mux2_2 _6091_ (.A0(\data_buffer[2][11] ),
    .A1(net506),
    .S(net1260),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_2 _6092_ (.A0(\data_buffer[2][12] ),
    .A1(net507),
    .S(net1260),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_2 _6093_ (.A0(\data_buffer[2][13] ),
    .A1(net508),
    .S(net1260),
    .X(_0994_));
 sky130_fd_sc_hd__mux2_2 _6094_ (.A0(\data_buffer[2][14] ),
    .A1(net509),
    .S(net1260),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_2 _6095_ (.A0(\data_buffer[2][15] ),
    .A1(net510),
    .S(net1260),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_2 _6096_ (.A0(\data_buffer[2][16] ),
    .A1(net512),
    .S(net1260),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_2 _6097_ (.A0(\data_buffer[2][17] ),
    .A1(net513),
    .S(net1260),
    .X(_0998_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input38 (.A(net1630),
    .X(net38));
 sky130_fd_sc_hd__mux2_2 _6099_ (.A0(\data_buffer[2][18] ),
    .A1(net514),
    .S(net1260),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_2 _6100_ (.A0(\data_buffer[2][19] ),
    .A1(net515),
    .S(net1260),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_2 _6101_ (.A0(\data_buffer[2][1] ),
    .A1(net495),
    .S(net1260),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_2 _6102_ (.A0(\data_buffer[2][20] ),
    .A1(net516),
    .S(net1260),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_2 _6103_ (.A0(\data_buffer[2][21] ),
    .A1(net517),
    .S(net1260),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_2 _6104_ (.A0(\data_buffer[2][22] ),
    .A1(net518),
    .S(net1260),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_2 _6105_ (.A0(\data_buffer[2][23] ),
    .A1(net519),
    .S(net1260),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_2 _6106_ (.A0(\data_buffer[2][24] ),
    .A1(net520),
    .S(net1260),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_2 _6107_ (.A0(\data_buffer[2][25] ),
    .A1(net521),
    .S(net1260),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_2 _6108_ (.A0(\data_buffer[2][26] ),
    .A1(net523),
    .S(net1260),
    .X(_1008_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input37 (.A(channel_dst_addr[17]),
    .X(net37));
 sky130_fd_sc_hd__mux2_2 _6110_ (.A0(\data_buffer[2][27] ),
    .A1(net524),
    .S(net1260),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_2 _6111_ (.A0(\data_buffer[2][28] ),
    .A1(net525),
    .S(net1260),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_2 _6112_ (.A0(\data_buffer[2][29] ),
    .A1(net526),
    .S(net1260),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_2 _6113_ (.A0(\data_buffer[2][2] ),
    .A1(net496),
    .S(net1260),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_2 _6114_ (.A0(\data_buffer[2][30] ),
    .A1(net527),
    .S(net1260),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_2 _6115_ (.A0(\data_buffer[2][31] ),
    .A1(net528),
    .S(net1260),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_2 _6116_ (.A0(\data_buffer[2][3] ),
    .A1(net497),
    .S(net1260),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_2 _6117_ (.A0(\data_buffer[2][4] ),
    .A1(net498),
    .S(net1260),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_2 _6118_ (.A0(\data_buffer[2][5] ),
    .A1(net499),
    .S(net1260),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_2 _6119_ (.A0(\data_buffer[2][6] ),
    .A1(net501),
    .S(net1260),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_2 _6120_ (.A0(\data_buffer[2][7] ),
    .A1(net502),
    .S(net1260),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_2 _6121_ (.A0(\data_buffer[2][8] ),
    .A1(net503),
    .S(net1260),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_2 _6122_ (.A0(\data_buffer[2][9] ),
    .A1(net504),
    .S(net1260),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_2 _6123_ (.A0(\data_buffer[3][0] ),
    .A1(net529),
    .S(net1261),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_2 _6124_ (.A0(\data_buffer[3][10] ),
    .A1(net413),
    .S(net1262),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_2 _6125_ (.A0(\data_buffer[3][11] ),
    .A1(net414),
    .S(net1261),
    .X(_1024_));
 sky130_fd_sc_hd__mux2_2 _6126_ (.A0(\data_buffer[3][12] ),
    .A1(net415),
    .S(net1261),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_2 _6127_ (.A0(\data_buffer[3][13] ),
    .A1(net416),
    .S(net1261),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_2 _6128_ (.A0(\data_buffer[3][14] ),
    .A1(net418),
    .S(net1261),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_2 _6129_ (.A0(\data_buffer[3][15] ),
    .A1(net419),
    .S(net1261),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_2 _6130_ (.A0(\data_buffer[3][16] ),
    .A1(net420),
    .S(net1261),
    .X(_1029_));
 sky130_fd_sc_hd__mux2_2 _6131_ (.A0(\data_buffer[3][17] ),
    .A1(net421),
    .S(net1261),
    .X(_1030_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input36 (.A(channel_dst_addr[16]),
    .X(net36));
 sky130_fd_sc_hd__mux2_2 _6133_ (.A0(\data_buffer[3][18] ),
    .A1(net422),
    .S(net1261),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_2 _6134_ (.A0(\data_buffer[3][19] ),
    .A1(net423),
    .S(net1261),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_2 _6135_ (.A0(\data_buffer[3][1] ),
    .A1(net530),
    .S(net1262),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_2 _6136_ (.A0(\data_buffer[3][20] ),
    .A1(net424),
    .S(net1261),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_2 _6137_ (.A0(\data_buffer[3][21] ),
    .A1(net425),
    .S(net1261),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_2 _6138_ (.A0(\data_buffer[3][22] ),
    .A1(net426),
    .S(net1261),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_2 _6139_ (.A0(\data_buffer[3][23] ),
    .A1(net427),
    .S(net1262),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_2 _6140_ (.A0(\data_buffer[3][24] ),
    .A1(net429),
    .S(net1261),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_2 _6141_ (.A0(\data_buffer[3][25] ),
    .A1(net430),
    .S(net1261),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_2 _6142_ (.A0(\data_buffer[3][26] ),
    .A1(net431),
    .S(net1261),
    .X(_1040_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input35 (.A(channel_dst_addr[15]),
    .X(net35));
 sky130_fd_sc_hd__mux2_2 _6144_ (.A0(\data_buffer[3][27] ),
    .A1(net432),
    .S(net1261),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_2 _6145_ (.A0(\data_buffer[3][28] ),
    .A1(net433),
    .S(net1261),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_2 _6146_ (.A0(\data_buffer[3][29] ),
    .A1(net434),
    .S(net1261),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_2 _6147_ (.A0(\data_buffer[3][2] ),
    .A1(net531),
    .S(net1261),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_2 _6148_ (.A0(\data_buffer[3][30] ),
    .A1(net435),
    .S(net1261),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_2 _6149_ (.A0(\data_buffer[3][31] ),
    .A1(net436),
    .S(net1261),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_2 _6150_ (.A0(\data_buffer[3][3] ),
    .A1(net532),
    .S(net1261),
    .X(_1047_));
 sky130_fd_sc_hd__mux2_2 _6151_ (.A0(\data_buffer[3][4] ),
    .A1(net407),
    .S(net1261),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_2 _6152_ (.A0(\data_buffer[3][5] ),
    .A1(net408),
    .S(net1262),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_2 _6153_ (.A0(\data_buffer[3][6] ),
    .A1(net409),
    .S(net1261),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_2 _6154_ (.A0(\data_buffer[3][7] ),
    .A1(net410),
    .S(net1262),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_2 _6155_ (.A0(\data_buffer[3][8] ),
    .A1(net411),
    .S(net1262),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_2 _6156_ (.A0(\data_buffer[3][9] ),
    .A1(net412),
    .S(net1262),
    .X(_1053_));
 sky130_fd_sc_hd__nand3b_1 _6157_ (.A_N(net558),
    .B(net554),
    .C(net557),
    .Y(_3372_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input34 (.A(net1597),
    .X(net34));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input33 (.A(channel_dst_addr[13]),
    .X(net33));
 sky130_fd_sc_hd__mux2_2 _6160_ (.A0(\current_dst_addr[0][0] ),
    .A1(net695),
    .S(net1255),
    .X(_1054_));
 sky130_fd_sc_hd__nand3_4 _6161_ (.A(_3214_),
    .B(net555),
    .C(net565),
    .Y(_3375_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input32 (.A(net1627),
    .X(net32));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input31 (.A(net1384),
    .X(net31));
 sky130_fd_sc_hd__nand2_1 _6164_ (.A(net696),
    .B(_3375_),
    .Y(_3378_));
 sky130_fd_sc_hd__o21ai_0 _6165_ (.A1(_1485_),
    .A2(_3375_),
    .B1(_3378_),
    .Y(_1055_));
 sky130_fd_sc_hd__mux2_2 _6166_ (.A0(\current_dst_addr[3][5] ),
    .A1(net697),
    .S(_3375_),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_2 _6167_ (.A0(\current_dst_addr[3][6] ),
    .A1(net698),
    .S(_3375_),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_2 _6168_ (.A0(\current_dst_addr[3][7] ),
    .A1(net699),
    .S(net1236),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_2 _6169_ (.A0(\current_dst_addr[3][8] ),
    .A1(net700),
    .S(net1236),
    .X(_1059_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input30 (.A(net1496),
    .X(net30));
 sky130_fd_sc_hd__mux2_2 _6171_ (.A0(\current_dst_addr[3][9] ),
    .A1(net701),
    .S(net1236),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_2 _6172_ (.A0(\current_dst_addr[3][10] ),
    .A1(net702),
    .S(net1236),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_2 _6173_ (.A0(\current_dst_addr[3][11] ),
    .A1(net703),
    .S(_3375_),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_2 _6174_ (.A0(\current_dst_addr[3][12] ),
    .A1(net704),
    .S(_3375_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_2 _6175_ (.A0(\current_dst_addr[3][13] ),
    .A1(net705),
    .S(_3375_),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_2 _6176_ (.A0(\current_dst_addr[0][10] ),
    .A1(net706),
    .S(net1255),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_2 _6177_ (.A0(\current_dst_addr[3][14] ),
    .A1(net707),
    .S(_3375_),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_2 _6178_ (.A0(\current_dst_addr[3][15] ),
    .A1(net708),
    .S(_3375_),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_2 _6179_ (.A0(\current_dst_addr[3][16] ),
    .A1(net709),
    .S(_3375_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_2 _6180_ (.A0(\current_dst_addr[3][17] ),
    .A1(net710),
    .S(_3375_),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_2 _6181_ (.A0(\current_dst_addr[3][18] ),
    .A1(net711),
    .S(_3375_),
    .X(_1070_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input29 (.A(net1418),
    .X(net29));
 sky130_fd_sc_hd__mux2_2 _6183_ (.A0(\current_dst_addr[3][19] ),
    .A1(net712),
    .S(_3375_),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_2 _6184_ (.A0(\current_dst_addr[3][20] ),
    .A1(net713),
    .S(_3375_),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_2 _6185_ (.A0(\current_dst_addr[3][21] ),
    .A1(net714),
    .S(_3375_),
    .X(_1073_));
 sky130_fd_sc_hd__mux2_2 _6186_ (.A0(\current_dst_addr[3][22] ),
    .A1(net715),
    .S(_3375_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_2 _6187_ (.A0(\current_dst_addr[3][23] ),
    .A1(net716),
    .S(_3375_),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_2 _6188_ (.A0(\current_dst_addr[0][11] ),
    .A1(net717),
    .S(net1256),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_2 _6189_ (.A0(\current_dst_addr[3][24] ),
    .A1(net718),
    .S(_3375_),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_2 _6190_ (.A0(\current_dst_addr[3][25] ),
    .A1(net719),
    .S(net1236),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_1 _6191_ (.A(net720),
    .B(_3375_),
    .Y(_3381_));
 sky130_fd_sc_hd__o21ai_0 _6192_ (.A1(_1583_),
    .A2(_3375_),
    .B1(_3381_),
    .Y(_1079_));
 sky130_fd_sc_hd__mux2_2 _6193_ (.A0(\current_dst_addr[3][27] ),
    .A1(net721),
    .S(_3375_),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_2 _6194_ (.A0(\current_dst_addr[3][28] ),
    .A1(net722),
    .S(_3375_),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_2 _6195_ (.A0(\current_dst_addr[3][29] ),
    .A1(net723),
    .S(_3375_),
    .X(_1082_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input28 (.A(net1444),
    .X(net28));
 sky130_fd_sc_hd__mux2_2 _6197_ (.A0(\current_dst_addr[3][30] ),
    .A1(net724),
    .S(net1236),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_2 _6198_ (.A0(\current_dst_addr[3][31] ),
    .A1(net725),
    .S(net1236),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_2 _6199_ (.A0(\current_dst_addr[0][12] ),
    .A1(net726),
    .S(net1256),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_2 _6200_ (.A0(\current_dst_addr[0][13] ),
    .A1(net727),
    .S(net1256),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_2 _6201_ (.A0(\current_dst_addr[0][14] ),
    .A1(net728),
    .S(net1255),
    .X(_1087_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input27 (.A(net1468),
    .X(net27));
 sky130_fd_sc_hd__mux2_2 _6203_ (.A0(\current_dst_addr[0][15] ),
    .A1(net729),
    .S(net1256),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_2 _6204_ (.A0(\current_dst_addr[0][16] ),
    .A1(net730),
    .S(net1255),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_2 _6205_ (.A0(\current_dst_addr[0][17] ),
    .A1(net731),
    .S(net1255),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_2 _6206_ (.A0(\current_dst_addr[0][18] ),
    .A1(net732),
    .S(net1256),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_2 _6207_ (.A0(\current_dst_addr[0][19] ),
    .A1(net733),
    .S(net1256),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_2 _6208_ (.A0(\current_dst_addr[0][1] ),
    .A1(net734),
    .S(net1255),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_2 _6209_ (.A0(\current_dst_addr[0][20] ),
    .A1(net735),
    .S(net1256),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_2 _6210_ (.A0(\current_dst_addr[0][21] ),
    .A1(net736),
    .S(net1255),
    .X(_1095_));
 sky130_fd_sc_hd__nand2_1 _6211_ (.A(net737),
    .B(net1255),
    .Y(_3384_));
 sky130_fd_sc_hd__o21ai_0 _6212_ (.A1(_1973_),
    .A2(net1255),
    .B1(_3384_),
    .Y(_1096_));
 sky130_fd_sc_hd__mux2_2 _6213_ (.A0(\current_dst_addr[0][23] ),
    .A1(net738),
    .S(net1255),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_2 _6214_ (.A0(\current_dst_addr[0][24] ),
    .A1(net739),
    .S(net1255),
    .X(_1098_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input26 (.A(net1631),
    .X(net26));
 sky130_fd_sc_hd__mux2_2 _6216_ (.A0(\current_dst_addr[0][25] ),
    .A1(net740),
    .S(net1256),
    .X(_1099_));
 sky130_fd_sc_hd__mux2_2 _6217_ (.A0(\current_dst_addr[0][26] ),
    .A1(net741),
    .S(net1256),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_2 _6218_ (.A0(\current_dst_addr[0][27] ),
    .A1(net742),
    .S(net1256),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_2 _6219_ (.A0(\current_dst_addr[0][28] ),
    .A1(net743),
    .S(net1256),
    .X(_1102_));
 sky130_fd_sc_hd__mux2_2 _6220_ (.A0(\current_dst_addr[0][29] ),
    .A1(net744),
    .S(net1255),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_2 _6221_ (.A0(\current_dst_addr[0][2] ),
    .A1(net745),
    .S(net1255),
    .X(_1104_));
 sky130_fd_sc_hd__mux2_2 _6222_ (.A0(\current_dst_addr[0][30] ),
    .A1(net746),
    .S(net1255),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_2 _6223_ (.A0(\current_dst_addr[0][31] ),
    .A1(net747),
    .S(net1255),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_2 _6224_ (.A0(\current_dst_addr[1][0] ),
    .A1(net748),
    .S(net1259),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_2 _6225_ (.A0(\current_dst_addr[1][1] ),
    .A1(net749),
    .S(net1259),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_2 _6226_ (.A0(\current_dst_addr[1][2] ),
    .A1(net750),
    .S(net1257),
    .X(_1109_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input25 (.A(net1586),
    .X(net25));
 sky130_fd_sc_hd__mux2_2 _6228_ (.A0(\current_dst_addr[1][3] ),
    .A1(net751),
    .S(net1257),
    .X(_1110_));
 sky130_fd_sc_hd__nand2_1 _6229_ (.A(net752),
    .B(net1257),
    .Y(_3387_));
 sky130_fd_sc_hd__o21ai_0 _6230_ (.A1(_1753_),
    .A2(net1257),
    .B1(_3387_),
    .Y(_1111_));
 sky130_fd_sc_hd__mux2_2 _6231_ (.A0(\current_dst_addr[1][5] ),
    .A1(net753),
    .S(net1257),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_2 _6232_ (.A0(\current_dst_addr[1][6] ),
    .A1(net754),
    .S(net1257),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_2 _6233_ (.A0(\current_dst_addr[1][7] ),
    .A1(net755),
    .S(net1257),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_2 _6234_ (.A0(\current_dst_addr[0][3] ),
    .A1(net756),
    .S(net1256),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_2 _6235_ (.A0(\current_dst_addr[1][8] ),
    .A1(net757),
    .S(net1257),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_2 _6236_ (.A0(\current_dst_addr[1][9] ),
    .A1(net758),
    .S(net1257),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_2 _6237_ (.A0(\current_dst_addr[1][10] ),
    .A1(net759),
    .S(net1258),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_2 _6238_ (.A0(\current_dst_addr[1][11] ),
    .A1(net760),
    .S(net1258),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_2 _6239_ (.A0(\current_dst_addr[1][12] ),
    .A1(net761),
    .S(net1258),
    .X(_1120_));
 sky130_fd_sc_hd__mux2_2 _6240_ (.A0(\current_dst_addr[1][13] ),
    .A1(net762),
    .S(net1257),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_1 _6241_ (.A(net763),
    .B(net1258),
    .Y(_3388_));
 sky130_fd_sc_hd__o21ai_0 _6242_ (.A1(_1801_),
    .A2(net1258),
    .B1(_3388_),
    .Y(_1122_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input24 (.A(net1622),
    .X(net24));
 sky130_fd_sc_hd__mux2_2 _6244_ (.A0(\current_dst_addr[1][15] ),
    .A1(net764),
    .S(net1257),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_2 _6245_ (.A0(\current_dst_addr[1][16] ),
    .A1(net765),
    .S(net1257),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_2 _6246_ (.A0(\current_dst_addr[1][17] ),
    .A1(net766),
    .S(net1258),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_2 _6247_ (.A0(\current_dst_addr[0][4] ),
    .A1(net767),
    .S(net1256),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_2 _6248_ (.A0(\current_dst_addr[1][18] ),
    .A1(net768),
    .S(net1257),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_2 _6249_ (.A0(\current_dst_addr[1][19] ),
    .A1(net769),
    .S(net1257),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_2 _6250_ (.A0(\current_dst_addr[1][20] ),
    .A1(net770),
    .S(net1257),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_2 _6251_ (.A0(\current_dst_addr[1][21] ),
    .A1(net771),
    .S(net1257),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_2 _6252_ (.A0(\current_dst_addr[1][22] ),
    .A1(net772),
    .S(net1257),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_2 _6253_ (.A0(\current_dst_addr[1][23] ),
    .A1(net773),
    .S(net1257),
    .X(_1132_));
 sky130_fd_sc_hd__mux2_2 _6254_ (.A0(\current_dst_addr[1][24] ),
    .A1(net774),
    .S(net1257),
    .X(_1133_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input23 (.A(net1638),
    .X(net23));
 sky130_fd_sc_hd__mux2_2 _6256_ (.A0(\current_dst_addr[1][25] ),
    .A1(net775),
    .S(net1257),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_2 _6257_ (.A0(\current_dst_addr[1][26] ),
    .A1(net776),
    .S(net1257),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_2 _6258_ (.A0(\current_dst_addr[1][27] ),
    .A1(net777),
    .S(net1257),
    .X(_1136_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input22 (.A(net1580),
    .X(net22));
 sky130_fd_sc_hd__mux2_2 _6260_ (.A0(\current_dst_addr[0][5] ),
    .A1(net778),
    .S(net1255),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_2 _6261_ (.A0(\current_dst_addr[1][28] ),
    .A1(net779),
    .S(net1257),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_2 _6262_ (.A0(\current_dst_addr[1][29] ),
    .A1(net780),
    .S(net1257),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_2 _6263_ (.A0(\current_dst_addr[1][30] ),
    .A1(net781),
    .S(net1257),
    .X(_1140_));
 sky130_fd_sc_hd__mux2_2 _6264_ (.A0(\current_dst_addr[1][31] ),
    .A1(net782),
    .S(net1257),
    .X(_1141_));
 sky130_fd_sc_hd__nand3_4 _6265_ (.A(_3269_),
    .B(net563),
    .C(net562),
    .Y(_3392_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input21 (.A(net1572),
    .X(net21));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input20 (.A(net1542),
    .X(net20));
 sky130_fd_sc_hd__mux2_2 _6268_ (.A0(\current_dst_addr[2][0] ),
    .A1(net783),
    .S(_3392_),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_2 _6269_ (.A0(\current_dst_addr[2][1] ),
    .A1(net784),
    .S(_3392_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_2 _6270_ (.A0(\current_dst_addr[2][2] ),
    .A1(net785),
    .S(_3392_),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_2 _6271_ (.A0(\current_dst_addr[2][3] ),
    .A1(net786),
    .S(_3392_),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_2 _6272_ (.A0(\current_dst_addr[2][4] ),
    .A1(net787),
    .S(_3392_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_2 _6273_ (.A0(\current_dst_addr[2][5] ),
    .A1(net788),
    .S(_3392_),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_2 _6274_ (.A0(\current_dst_addr[0][6] ),
    .A1(net789),
    .S(net1255),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_2 _6275_ (.A0(\current_dst_addr[2][6] ),
    .A1(net790),
    .S(_3392_),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_2 _6276_ (.A0(\current_dst_addr[2][7] ),
    .A1(net791),
    .S(_3392_),
    .X(_1150_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input19 (.A(net1618),
    .X(net19));
 sky130_fd_sc_hd__mux2_2 _6278_ (.A0(\current_dst_addr[2][8] ),
    .A1(net792),
    .S(_3392_),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_2 _6279_ (.A0(\current_dst_addr[2][9] ),
    .A1(net793),
    .S(_3392_),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_2 _6280_ (.A0(\current_dst_addr[2][10] ),
    .A1(net794),
    .S(_3392_),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_2 _6281_ (.A0(\current_dst_addr[2][11] ),
    .A1(net795),
    .S(_3392_),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_2 _6282_ (.A0(\current_dst_addr[2][12] ),
    .A1(net796),
    .S(_3392_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_2 _6283_ (.A0(\current_dst_addr[2][13] ),
    .A1(net797),
    .S(_3392_),
    .X(_1156_));
 sky130_fd_sc_hd__mux2_2 _6284_ (.A0(\current_dst_addr[2][14] ),
    .A1(net798),
    .S(_3392_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_2 _6285_ (.A0(\current_dst_addr[2][15] ),
    .A1(net799),
    .S(_3392_),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_2 _6286_ (.A0(\current_dst_addr[0][7] ),
    .A1(net800),
    .S(net1255),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_2 _6287_ (.A0(\current_dst_addr[2][16] ),
    .A1(net801),
    .S(_3392_),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_2 _6288_ (.A0(\current_dst_addr[2][17] ),
    .A1(net802),
    .S(_3392_),
    .X(_1161_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input18 (.A(net1499),
    .X(net18));
 sky130_fd_sc_hd__mux2_2 _6290_ (.A0(\current_dst_addr[2][18] ),
    .A1(net803),
    .S(_3392_),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_2 _6291_ (.A0(\current_dst_addr[2][19] ),
    .A1(net804),
    .S(_3392_),
    .X(_1163_));
 sky130_fd_sc_hd__mux2_2 _6292_ (.A0(\current_dst_addr[2][20] ),
    .A1(net805),
    .S(_3392_),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_2 _6293_ (.A0(\current_dst_addr[2][21] ),
    .A1(net806),
    .S(_3392_),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_2 _6294_ (.A0(\current_dst_addr[2][22] ),
    .A1(net807),
    .S(_3392_),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_2 _6295_ (.A0(\current_dst_addr[2][23] ),
    .A1(net808),
    .S(_3392_),
    .X(_1167_));
 sky130_fd_sc_hd__mux2_2 _6296_ (.A0(\current_dst_addr[2][24] ),
    .A1(net809),
    .S(_3392_),
    .X(_1168_));
 sky130_fd_sc_hd__mux2_2 _6297_ (.A0(\current_dst_addr[2][25] ),
    .A1(net810),
    .S(net1235),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_2 _6298_ (.A0(\current_dst_addr[0][8] ),
    .A1(net811),
    .S(net1255),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_2 _6299_ (.A0(\current_dst_addr[2][26] ),
    .A1(net812),
    .S(net1235),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_2 _6300_ (.A0(\current_dst_addr[2][27] ),
    .A1(net813),
    .S(net1235),
    .X(_1172_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input17 (.A(net1372),
    .X(net17));
 sky130_fd_sc_hd__mux2_2 _6302_ (.A0(\current_dst_addr[2][28] ),
    .A1(net814),
    .S(net1235),
    .X(_1173_));
 sky130_fd_sc_hd__mux2_2 _6303_ (.A0(\current_dst_addr[2][29] ),
    .A1(net815),
    .S(net1235),
    .X(_1174_));
 sky130_fd_sc_hd__mux2_2 _6304_ (.A0(\current_dst_addr[2][30] ),
    .A1(net816),
    .S(_3392_),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_2 _6305_ (.A0(\current_dst_addr[2][31] ),
    .A1(net817),
    .S(_3392_),
    .X(_1176_));
 sky130_fd_sc_hd__mux2_2 _6306_ (.A0(\current_dst_addr[3][0] ),
    .A1(net818),
    .S(_3375_),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_2 _6307_ (.A0(\current_dst_addr[3][1] ),
    .A1(net819),
    .S(_3375_),
    .X(_1178_));
 sky130_fd_sc_hd__mux2_2 _6308_ (.A0(\current_dst_addr[3][2] ),
    .A1(net820),
    .S(net1236),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_2 _6309_ (.A0(\current_dst_addr[3][3] ),
    .A1(net821),
    .S(_3375_),
    .X(_1180_));
 sky130_fd_sc_hd__mux2_2 _6310_ (.A0(\current_dst_addr[0][9] ),
    .A1(net822),
    .S(net1256),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_2 _6311_ (.A0(\data_buffer[0][0] ),
    .A1(net823),
    .S(net1255),
    .X(_1182_));
 sky130_fd_sc_hd__mux2_2 _6312_ (.A0(\data_buffer[3][4] ),
    .A1(net824),
    .S(net1236),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_2 _6313_ (.A0(\data_buffer[3][5] ),
    .A1(net825),
    .S(_3375_),
    .X(_1184_));
 sky130_fd_sc_hd__mux2_2 _6314_ (.A0(\data_buffer[3][6] ),
    .A1(net826),
    .S(net1236),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_2 _6315_ (.A0(\data_buffer[3][7] ),
    .A1(net827),
    .S(_3375_),
    .X(_1186_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input16 (.A(net1483),
    .X(net16));
 sky130_fd_sc_hd__mux2_2 _6317_ (.A0(\data_buffer[3][8] ),
    .A1(net828),
    .S(_3375_),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_2 _6318_ (.A0(\data_buffer[3][9] ),
    .A1(net829),
    .S(_3375_),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_2 _6319_ (.A0(\data_buffer[3][10] ),
    .A1(net830),
    .S(_3375_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_2 _6320_ (.A0(\data_buffer[3][11] ),
    .A1(net831),
    .S(net1236),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_2 _6321_ (.A0(\data_buffer[3][12] ),
    .A1(net832),
    .S(net1236),
    .X(_1191_));
 sky130_fd_sc_hd__mux2_2 _6322_ (.A0(\data_buffer[3][13] ),
    .A1(net833),
    .S(net1236),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_2 _6323_ (.A0(\data_buffer[0][10] ),
    .A1(net834),
    .S(net1255),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_2 _6324_ (.A0(\data_buffer[3][14] ),
    .A1(net835),
    .S(net1236),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_2 _6325_ (.A0(\data_buffer[3][15] ),
    .A1(net836),
    .S(net1236),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_2 _6326_ (.A0(\data_buffer[3][16] ),
    .A1(net837),
    .S(net1236),
    .X(_1196_));
 sky130_fd_sc_hd__mux2_2 _6327_ (.A0(\data_buffer[3][17] ),
    .A1(net838),
    .S(net1236),
    .X(_1197_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input15 (.A(net1605),
    .X(net15));
 sky130_fd_sc_hd__mux2_2 _6329_ (.A0(\data_buffer[3][18] ),
    .A1(net839),
    .S(net1236),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_2 _6330_ (.A0(\data_buffer[3][19] ),
    .A1(net840),
    .S(net1236),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_2 _6331_ (.A0(\data_buffer[3][20] ),
    .A1(net841),
    .S(net1236),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_2 _6332_ (.A0(\data_buffer[3][21] ),
    .A1(net842),
    .S(net1236),
    .X(_1201_));
 sky130_fd_sc_hd__mux2_2 _6333_ (.A0(\data_buffer[3][22] ),
    .A1(net843),
    .S(net1236),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_2 _6334_ (.A0(\data_buffer[3][23] ),
    .A1(net844),
    .S(_3375_),
    .X(_1203_));
 sky130_fd_sc_hd__mux2_2 _6335_ (.A0(\data_buffer[0][11] ),
    .A1(net845),
    .S(net1255),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_2 _6336_ (.A0(\data_buffer[3][24] ),
    .A1(net846),
    .S(net1236),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_2 _6337_ (.A0(\data_buffer[3][25] ),
    .A1(net847),
    .S(net1236),
    .X(_1206_));
 sky130_fd_sc_hd__mux2_2 _6338_ (.A0(\data_buffer[3][26] ),
    .A1(net848),
    .S(net1236),
    .X(_1207_));
 sky130_fd_sc_hd__mux2_2 _6339_ (.A0(\data_buffer[3][27] ),
    .A1(net849),
    .S(net1236),
    .X(_1208_));
 sky130_fd_sc_hd__mux2_2 _6340_ (.A0(\data_buffer[3][28] ),
    .A1(net850),
    .S(net1236),
    .X(_1209_));
 sky130_fd_sc_hd__mux2_2 _6341_ (.A0(\data_buffer[3][29] ),
    .A1(net851),
    .S(net1236),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_2 _6342_ (.A0(\data_buffer[3][30] ),
    .A1(net852),
    .S(net1236),
    .X(_1211_));
 sky130_fd_sc_hd__mux2_2 _6343_ (.A0(\data_buffer[3][31] ),
    .A1(net853),
    .S(net1236),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_2 _6344_ (.A0(\data_buffer[0][12] ),
    .A1(net854),
    .S(net1255),
    .X(_1213_));
 sky130_fd_sc_hd__mux2_2 _6345_ (.A0(\data_buffer[0][13] ),
    .A1(net855),
    .S(net1255),
    .X(_1214_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input14 (.A(net1492),
    .X(net14));
 sky130_fd_sc_hd__mux2_2 _6347_ (.A0(\data_buffer[0][14] ),
    .A1(net856),
    .S(net1255),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_2 _6348_ (.A0(\data_buffer[0][15] ),
    .A1(net857),
    .S(net1255),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_2 _6349_ (.A0(\data_buffer[0][16] ),
    .A1(net858),
    .S(net1255),
    .X(_1217_));
 sky130_fd_sc_hd__mux2_2 _6350_ (.A0(\data_buffer[0][17] ),
    .A1(net859),
    .S(net1255),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_2 _6351_ (.A0(\data_buffer[0][18] ),
    .A1(net860),
    .S(net1255),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_2 _6352_ (.A0(\data_buffer[0][19] ),
    .A1(net861),
    .S(net1255),
    .X(_1220_));
 sky130_fd_sc_hd__mux2_2 _6353_ (.A0(\data_buffer[0][1] ),
    .A1(net862),
    .S(net1255),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_2 _6354_ (.A0(\data_buffer[0][20] ),
    .A1(net863),
    .S(net1255),
    .X(_1222_));
 sky130_fd_sc_hd__mux2_2 _6355_ (.A0(\data_buffer[0][21] ),
    .A1(net864),
    .S(net1255),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_2 _6356_ (.A0(\data_buffer[0][22] ),
    .A1(net865),
    .S(net1255),
    .X(_1224_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input13 (.A(net1528),
    .X(net13));
 sky130_fd_sc_hd__mux2_2 _6358_ (.A0(\data_buffer[0][23] ),
    .A1(net866),
    .S(net1255),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_2 _6359_ (.A0(\data_buffer[0][24] ),
    .A1(net867),
    .S(net1255),
    .X(_1226_));
 sky130_fd_sc_hd__mux2_2 _6360_ (.A0(\data_buffer[0][25] ),
    .A1(net868),
    .S(net1255),
    .X(_1227_));
 sky130_fd_sc_hd__mux2_2 _6361_ (.A0(\data_buffer[0][26] ),
    .A1(net869),
    .S(net1255),
    .X(_1228_));
 sky130_fd_sc_hd__mux2_2 _6362_ (.A0(\data_buffer[0][27] ),
    .A1(net870),
    .S(net1255),
    .X(_1229_));
 sky130_fd_sc_hd__mux2_2 _6363_ (.A0(\data_buffer[0][28] ),
    .A1(net871),
    .S(net1255),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_2 _6364_ (.A0(\data_buffer[0][29] ),
    .A1(net872),
    .S(net1255),
    .X(_1231_));
 sky130_fd_sc_hd__mux2_2 _6365_ (.A0(\data_buffer[0][2] ),
    .A1(net873),
    .S(net1255),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_2 _6366_ (.A0(\data_buffer[0][30] ),
    .A1(net874),
    .S(net1255),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_2 _6367_ (.A0(\data_buffer[0][31] ),
    .A1(net875),
    .S(net1255),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_2 _6368_ (.A0(\data_buffer[1][0] ),
    .A1(net876),
    .S(net1259),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_2 _6369_ (.A0(\data_buffer[1][1] ),
    .A1(net877),
    .S(net1259),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_2 _6370_ (.A0(\data_buffer[1][2] ),
    .A1(net878),
    .S(net1259),
    .X(_1237_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input12 (.A(channel_dst_addr[10]),
    .X(net12));
 sky130_fd_sc_hd__mux2_2 _6372_ (.A0(\data_buffer[1][3] ),
    .A1(net879),
    .S(net1259),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_2 _6373_ (.A0(\data_buffer[1][4] ),
    .A1(net880),
    .S(net1259),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_2 _6374_ (.A0(\data_buffer[1][5] ),
    .A1(net881),
    .S(net1259),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_2 _6375_ (.A0(\data_buffer[1][6] ),
    .A1(net882),
    .S(net1259),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_2 _6376_ (.A0(\data_buffer[1][7] ),
    .A1(net883),
    .S(net1259),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_2 _6377_ (.A0(\data_buffer[0][3] ),
    .A1(net884),
    .S(net1255),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_2 _6378_ (.A0(\data_buffer[1][8] ),
    .A1(net885),
    .S(net1259),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_2 _6379_ (.A0(\data_buffer[1][9] ),
    .A1(net886),
    .S(net1259),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_2 _6380_ (.A0(\data_buffer[1][10] ),
    .A1(net887),
    .S(net1259),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_2 _6381_ (.A0(\data_buffer[1][11] ),
    .A1(net888),
    .S(net1259),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_2 _6382_ (.A0(\data_buffer[1][12] ),
    .A1(net889),
    .S(net1259),
    .X(_1248_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input11 (.A(net1485),
    .X(net11));
 sky130_fd_sc_hd__mux2_2 _6384_ (.A0(\data_buffer[1][13] ),
    .A1(net890),
    .S(net1259),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_2 _6385_ (.A0(\data_buffer[1][14] ),
    .A1(net891),
    .S(net1259),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_2 _6386_ (.A0(\data_buffer[1][15] ),
    .A1(net892),
    .S(net1259),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_2 _6387_ (.A0(\data_buffer[1][16] ),
    .A1(net893),
    .S(net1259),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_2 _6388_ (.A0(\data_buffer[1][17] ),
    .A1(net894),
    .S(net1259),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_2 _6389_ (.A0(\data_buffer[0][4] ),
    .A1(net895),
    .S(net1255),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_2 _6390_ (.A0(\data_buffer[1][18] ),
    .A1(net896),
    .S(net1259),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_2 _6391_ (.A0(\data_buffer[1][19] ),
    .A1(net897),
    .S(net1259),
    .X(_1256_));
 sky130_fd_sc_hd__mux2_2 _6392_ (.A0(\data_buffer[1][20] ),
    .A1(net898),
    .S(net1259),
    .X(_1257_));
 sky130_fd_sc_hd__mux2_2 _6393_ (.A0(\data_buffer[1][21] ),
    .A1(net899),
    .S(net1259),
    .X(_1258_));
 sky130_fd_sc_hd__mux2_2 _6394_ (.A0(\data_buffer[1][22] ),
    .A1(net900),
    .S(net1259),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_2 _6395_ (.A0(\data_buffer[1][23] ),
    .A1(net901),
    .S(net1259),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_2 _6396_ (.A0(\data_buffer[1][24] ),
    .A1(net902),
    .S(net1259),
    .X(_1261_));
 sky130_fd_sc_hd__mux2_2 _6397_ (.A0(\data_buffer[1][25] ),
    .A1(net903),
    .S(net1259),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_2 _6398_ (.A0(\data_buffer[1][26] ),
    .A1(net904),
    .S(net1259),
    .X(_1263_));
 sky130_fd_sc_hd__mux2_2 _6399_ (.A0(\data_buffer[1][27] ),
    .A1(net905),
    .S(net1259),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_2 _6400_ (.A0(\data_buffer[0][5] ),
    .A1(net906),
    .S(net1255),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_2 _6401_ (.A0(\data_buffer[1][28] ),
    .A1(net907),
    .S(net1259),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_2 _6402_ (.A0(\data_buffer[1][29] ),
    .A1(net908),
    .S(net1259),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_2 _6403_ (.A0(\data_buffer[1][30] ),
    .A1(net909),
    .S(net1259),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_2 _6404_ (.A0(\data_buffer[1][31] ),
    .A1(net910),
    .S(net1259),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_2 _6405_ (.A0(\data_buffer[2][0] ),
    .A1(net911),
    .S(net1235),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_2 _6406_ (.A0(\data_buffer[2][1] ),
    .A1(net912),
    .S(net1235),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_2 _6407_ (.A0(\data_buffer[2][2] ),
    .A1(net913),
    .S(net1235),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_2 _6408_ (.A0(\data_buffer[2][3] ),
    .A1(net914),
    .S(net1235),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_2 _6409_ (.A0(\data_buffer[2][4] ),
    .A1(net915),
    .S(net1235),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_2 _6410_ (.A0(\data_buffer[2][5] ),
    .A1(net916),
    .S(net1235),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_2 _6411_ (.A0(\data_buffer[0][6] ),
    .A1(net917),
    .S(net1255),
    .X(_1276_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input10 (.A(net1498),
    .X(net10));
 sky130_fd_sc_hd__mux2_2 _6413_ (.A0(\data_buffer[2][6] ),
    .A1(net918),
    .S(net1235),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_2 _6414_ (.A0(\data_buffer[2][7] ),
    .A1(net919),
    .S(net1235),
    .X(_1278_));
 sky130_fd_sc_hd__mux2_2 _6415_ (.A0(\data_buffer[2][8] ),
    .A1(net920),
    .S(net1235),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_2 _6416_ (.A0(\data_buffer[2][9] ),
    .A1(net921),
    .S(net1235),
    .X(_1280_));
 sky130_fd_sc_hd__mux2_2 _6417_ (.A0(\data_buffer[2][10] ),
    .A1(net922),
    .S(net1235),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_2 _6418_ (.A0(\data_buffer[2][11] ),
    .A1(net923),
    .S(net1235),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_2 _6419_ (.A0(\data_buffer[2][12] ),
    .A1(net924),
    .S(net1235),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_2 _6420_ (.A0(\data_buffer[2][13] ),
    .A1(net925),
    .S(net1235),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_2 _6421_ (.A0(\data_buffer[2][14] ),
    .A1(net926),
    .S(net1235),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_2 _6422_ (.A0(\data_buffer[2][15] ),
    .A1(net927),
    .S(net1235),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_2 _6423_ (.A0(\data_buffer[0][7] ),
    .A1(net928),
    .S(net1255),
    .X(_1287_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input9 (.A(net1634),
    .X(net9));
 sky130_fd_sc_hd__mux2_2 _6425_ (.A0(\data_buffer[2][16] ),
    .A1(net929),
    .S(net1235),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_2 _6426_ (.A0(\data_buffer[2][17] ),
    .A1(net930),
    .S(net1235),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_2 _6427_ (.A0(\data_buffer[2][18] ),
    .A1(net931),
    .S(net1235),
    .X(_1290_));
 sky130_fd_sc_hd__mux2_2 _6428_ (.A0(\data_buffer[2][19] ),
    .A1(net932),
    .S(net1235),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_2 _6429_ (.A0(\data_buffer[2][20] ),
    .A1(net933),
    .S(net1235),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_2 _6430_ (.A0(\data_buffer[2][21] ),
    .A1(net934),
    .S(net1235),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_2 _6431_ (.A0(\data_buffer[2][22] ),
    .A1(net935),
    .S(net1235),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_2 _6432_ (.A0(\data_buffer[2][23] ),
    .A1(net936),
    .S(net1235),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_2 _6433_ (.A0(\data_buffer[2][24] ),
    .A1(net937),
    .S(net1235),
    .X(_1296_));
 sky130_fd_sc_hd__mux2_2 _6434_ (.A0(\data_buffer[2][25] ),
    .A1(net938),
    .S(net1235),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_2 _6435_ (.A0(\data_buffer[0][8] ),
    .A1(net939),
    .S(net1255),
    .X(_1298_));
 sky130_fd_sc_hd__mux2_2 _6436_ (.A0(\data_buffer[2][26] ),
    .A1(net940),
    .S(net1235),
    .X(_1299_));
 sky130_fd_sc_hd__mux2_2 _6437_ (.A0(\data_buffer[2][27] ),
    .A1(net941),
    .S(net1235),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_2 _6438_ (.A0(\data_buffer[2][28] ),
    .A1(net942),
    .S(net1235),
    .X(_1301_));
 sky130_fd_sc_hd__mux2_2 _6439_ (.A0(\data_buffer[2][29] ),
    .A1(net943),
    .S(net1235),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_2 _6440_ (.A0(\data_buffer[2][30] ),
    .A1(net944),
    .S(net1235),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_2 _6441_ (.A0(\data_buffer[2][31] ),
    .A1(net945),
    .S(net1235),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_2 _6442_ (.A0(\data_buffer[3][0] ),
    .A1(net946),
    .S(net1236),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_2 _6443_ (.A0(\data_buffer[3][1] ),
    .A1(net947),
    .S(_3375_),
    .X(_1306_));
 sky130_fd_sc_hd__mux2_2 _6444_ (.A0(\data_buffer[3][2] ),
    .A1(net948),
    .S(net1236),
    .X(_1307_));
 sky130_fd_sc_hd__mux2_2 _6445_ (.A0(\data_buffer[3][3] ),
    .A1(net949),
    .S(net1236),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_2 _6446_ (.A0(\data_buffer[0][9] ),
    .A1(net950),
    .S(net1255),
    .X(_1309_));
 sky130_fd_sc_hd__o21ai_0 _6447_ (.A1(net557),
    .A2(_3314_),
    .B1(net1256),
    .Y(_1310_));
 sky130_fd_sc_hd__nand2b_1 _6448_ (.A_N(net1273),
    .B(net1271),
    .Y(_3406_));
 sky130_fd_sc_hd__o21ai_0 _6449_ (.A1(net1272),
    .A2(_3406_),
    .B1(net1257),
    .Y(_1311_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(_3287_),
    .B(_3392_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _6451_ (.A(_3277_),
    .B(_3375_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2b_1 _6452_ (.A_N(net957),
    .B(net1235),
    .Y(_1314_));
 sky130_fd_sc_hd__nand2b_1 _6453_ (.A_N(net961),
    .B(_3375_),
    .Y(_1315_));
 sky130_fd_sc_hd__nand2b_1 _6454_ (.A_N(net964),
    .B(net1255),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2b_1 _6455_ (.A_N(net968),
    .B(net1259),
    .Y(_1317_));
 sky130_fd_sc_hd__mux2_2 _6456_ (.A0(net971),
    .A1(\current_src_addr[0][0] ),
    .S(net1252),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_2 _6457_ (.A0(net972),
    .A1(\current_src_addr[3][4] ),
    .S(net1253),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_2 _6458_ (.A0(net973),
    .A1(\current_src_addr[3][5] ),
    .S(net1253),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_2 _6459_ (.A0(net974),
    .A1(\current_src_addr[3][6] ),
    .S(net1253),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_2 _6460_ (.A0(net975),
    .A1(\current_src_addr[3][7] ),
    .S(net1253),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_2 _6461_ (.A0(net976),
    .A1(\current_src_addr[3][8] ),
    .S(net1253),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_2 _6462_ (.A0(net977),
    .A1(\current_src_addr[3][9] ),
    .S(net1253),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_2 _6463_ (.A0(net978),
    .A1(\current_src_addr[3][10] ),
    .S(net1253),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_2 _6464_ (.A0(net979),
    .A1(\current_src_addr[3][11] ),
    .S(net1253),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_2 _6465_ (.A0(net980),
    .A1(\current_src_addr[3][12] ),
    .S(net1253),
    .X(_1327_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input8 (.A(net1472),
    .X(net8));
 sky130_fd_sc_hd__mux2_2 _6467_ (.A0(net981),
    .A1(\current_src_addr[3][13] ),
    .S(net1253),
    .X(_1328_));
 sky130_fd_sc_hd__mux2_2 _6468_ (.A0(net982),
    .A1(\current_src_addr[0][10] ),
    .S(net1252),
    .X(_1329_));
 sky130_fd_sc_hd__mux2_2 _6469_ (.A0(net983),
    .A1(\current_src_addr[3][14] ),
    .S(net1253),
    .X(_1330_));
 sky130_fd_sc_hd__mux2_2 _6470_ (.A0(net984),
    .A1(\current_src_addr[3][15] ),
    .S(net1253),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_2 _6471_ (.A0(net985),
    .A1(\current_src_addr[3][16] ),
    .S(net1253),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_2 _6472_ (.A0(net986),
    .A1(\current_src_addr[3][17] ),
    .S(net1253),
    .X(_1333_));
 sky130_fd_sc_hd__mux2_2 _6473_ (.A0(net987),
    .A1(\current_src_addr[3][18] ),
    .S(net1253),
    .X(_1334_));
 sky130_fd_sc_hd__mux2_2 _6474_ (.A0(net988),
    .A1(\current_src_addr[3][19] ),
    .S(net1253),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_2 _6475_ (.A0(net989),
    .A1(\current_src_addr[3][20] ),
    .S(net1253),
    .X(_1336_));
 sky130_fd_sc_hd__mux2_2 _6476_ (.A0(net990),
    .A1(\current_src_addr[3][21] ),
    .S(net1253),
    .X(_1337_));
 sky130_fd_sc_hd__mux2_2 _6477_ (.A0(net991),
    .A1(\current_src_addr[3][22] ),
    .S(net1253),
    .X(_1338_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input7 (.A(net1417),
    .X(net7));
 sky130_fd_sc_hd__mux2_2 _6479_ (.A0(net992),
    .A1(\current_src_addr[3][23] ),
    .S(net1253),
    .X(_1339_));
 sky130_fd_sc_hd__mux2_2 _6480_ (.A0(net993),
    .A1(\current_src_addr[0][11] ),
    .S(net1252),
    .X(_1340_));
 sky130_fd_sc_hd__mux2_2 _6481_ (.A0(net994),
    .A1(\current_src_addr[3][24] ),
    .S(net1253),
    .X(_1341_));
 sky130_fd_sc_hd__mux2_2 _6482_ (.A0(net995),
    .A1(\current_src_addr[3][25] ),
    .S(net1253),
    .X(_1342_));
 sky130_fd_sc_hd__mux2_2 _6483_ (.A0(net996),
    .A1(\current_src_addr[3][26] ),
    .S(net1253),
    .X(_1343_));
 sky130_fd_sc_hd__mux2_2 _6484_ (.A0(net997),
    .A1(\current_src_addr[3][27] ),
    .S(net1253),
    .X(_1344_));
 sky130_fd_sc_hd__mux2_2 _6485_ (.A0(net998),
    .A1(\current_src_addr[3][28] ),
    .S(net1253),
    .X(_1345_));
 sky130_fd_sc_hd__mux2_2 _6486_ (.A0(net999),
    .A1(\current_src_addr[3][29] ),
    .S(net1253),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_2 _6487_ (.A0(net1000),
    .A1(\current_src_addr[3][30] ),
    .S(net1253),
    .X(_1347_));
 sky130_fd_sc_hd__mux2_2 _6488_ (.A0(net1001),
    .A1(\current_src_addr[3][31] ),
    .S(net1253),
    .X(_1348_));
 sky130_fd_sc_hd__mux2_2 _6489_ (.A0(net1002),
    .A1(\current_src_addr[0][12] ),
    .S(net1252),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_2 _6490_ (.A0(net1003),
    .A1(\current_src_addr[0][13] ),
    .S(net1252),
    .X(_1350_));
 sky130_fd_sc_hd__mux2_2 _6491_ (.A0(net1004),
    .A1(\current_src_addr[0][14] ),
    .S(net1252),
    .X(_1351_));
 sky130_fd_sc_hd__mux2_2 _6492_ (.A0(net1005),
    .A1(\current_src_addr[0][15] ),
    .S(net1252),
    .X(_1352_));
 sky130_fd_sc_hd__mux2_2 _6493_ (.A0(net1006),
    .A1(\current_src_addr[0][16] ),
    .S(net1252),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_2 _6494_ (.A0(net1007),
    .A1(\current_src_addr[0][17] ),
    .S(net1252),
    .X(_1354_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input6 (.A(net1507),
    .X(net6));
 sky130_fd_sc_hd__mux2_2 _6496_ (.A0(net1008),
    .A1(\current_src_addr[0][18] ),
    .S(net1252),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_2 _6497_ (.A0(net1009),
    .A1(\current_src_addr[0][19] ),
    .S(net1252),
    .X(_1356_));
 sky130_fd_sc_hd__mux2_2 _6498_ (.A0(net1010),
    .A1(\current_src_addr[0][1] ),
    .S(net1252),
    .X(_1357_));
 sky130_fd_sc_hd__mux2_2 _6499_ (.A0(net1011),
    .A1(\current_src_addr[0][20] ),
    .S(net1252),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_2 _6500_ (.A0(net1012),
    .A1(\current_src_addr[0][21] ),
    .S(net1252),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_2 _6501_ (.A0(net1013),
    .A1(\current_src_addr[0][22] ),
    .S(net1252),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_2 _6502_ (.A0(net1014),
    .A1(\current_src_addr[0][23] ),
    .S(net1252),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_2 _6503_ (.A0(net1015),
    .A1(\current_src_addr[0][24] ),
    .S(net1252),
    .X(_1362_));
 sky130_fd_sc_hd__mux2_2 _6504_ (.A0(net1016),
    .A1(\current_src_addr[0][25] ),
    .S(net1252),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_2 _6505_ (.A0(net1017),
    .A1(\current_src_addr[0][26] ),
    .S(net1252),
    .X(_1364_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input5 (.A(net1590),
    .X(net5));
 sky130_fd_sc_hd__mux2_2 _6507_ (.A0(net1018),
    .A1(\current_src_addr[0][27] ),
    .S(net1252),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_2 _6508_ (.A0(net1019),
    .A1(\current_src_addr[0][28] ),
    .S(net1252),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_2 _6509_ (.A0(net1020),
    .A1(\current_src_addr[0][29] ),
    .S(net1252),
    .X(_1367_));
 sky130_fd_sc_hd__mux2_2 _6510_ (.A0(net1021),
    .A1(\current_src_addr[0][2] ),
    .S(net1252),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_2 _6511_ (.A0(net1022),
    .A1(\current_src_addr[0][30] ),
    .S(net1252),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_2 _6512_ (.A0(net1023),
    .A1(\current_src_addr[0][31] ),
    .S(net1252),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_2 _6513_ (.A0(net1024),
    .A1(\current_src_addr[1][0] ),
    .S(net1269),
    .X(_1371_));
 sky130_fd_sc_hd__mux2_2 _6514_ (.A0(net1025),
    .A1(\current_src_addr[1][1] ),
    .S(net1269),
    .X(_1372_));
 sky130_fd_sc_hd__mux2_2 _6515_ (.A0(net1026),
    .A1(\current_src_addr[1][2] ),
    .S(net1269),
    .X(_1373_));
 sky130_fd_sc_hd__mux2_2 _6516_ (.A0(net1027),
    .A1(\current_src_addr[1][3] ),
    .S(net1269),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_2 _6517_ (.A0(net1028),
    .A1(\current_src_addr[1][4] ),
    .S(net1269),
    .X(_1375_));
 sky130_fd_sc_hd__mux2_2 _6518_ (.A0(net1029),
    .A1(\current_src_addr[1][5] ),
    .S(net1269),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_2 _6519_ (.A0(net1030),
    .A1(\current_src_addr[1][6] ),
    .S(net1269),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_2 _6520_ (.A0(net1031),
    .A1(\current_src_addr[1][7] ),
    .S(net1269),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_2 _6521_ (.A0(net1032),
    .A1(\current_src_addr[0][3] ),
    .S(net1252),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_2 _6522_ (.A0(net1033),
    .A1(\current_src_addr[1][8] ),
    .S(net1269),
    .X(_1380_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input4 (.A(net1453),
    .X(net4));
 sky130_fd_sc_hd__mux2_2 _6524_ (.A0(net1034),
    .A1(\current_src_addr[1][9] ),
    .S(net1269),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_2 _6525_ (.A0(net1035),
    .A1(\current_src_addr[1][10] ),
    .S(net1269),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_2 _6526_ (.A0(net1036),
    .A1(\current_src_addr[1][11] ),
    .S(net1269),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_2 _6527_ (.A0(net1037),
    .A1(\current_src_addr[1][12] ),
    .S(net1269),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_2 _6528_ (.A0(net1038),
    .A1(\current_src_addr[1][13] ),
    .S(net1269),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_2 _6529_ (.A0(net1039),
    .A1(\current_src_addr[1][14] ),
    .S(net1269),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_2 _6530_ (.A0(net1040),
    .A1(\current_src_addr[1][15] ),
    .S(net1269),
    .X(_1387_));
 sky130_fd_sc_hd__mux2_2 _6531_ (.A0(net1041),
    .A1(\current_src_addr[1][16] ),
    .S(net1269),
    .X(_1388_));
 sky130_fd_sc_hd__mux2_2 _6532_ (.A0(net1042),
    .A1(\current_src_addr[1][17] ),
    .S(net1269),
    .X(_1389_));
 sky130_fd_sc_hd__mux2_2 _6533_ (.A0(net1043),
    .A1(\current_src_addr[0][4] ),
    .S(net1252),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_2 _6534_ (.A0(net1044),
    .A1(\current_src_addr[1][18] ),
    .S(net1269),
    .X(_1391_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input3 (.A(net1501),
    .X(net3));
 sky130_fd_sc_hd__mux2_2 _6536_ (.A0(net1045),
    .A1(\current_src_addr[1][19] ),
    .S(net1269),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_2 _6537_ (.A0(net1046),
    .A1(\current_src_addr[1][20] ),
    .S(net1269),
    .X(_1393_));
 sky130_fd_sc_hd__mux2_2 _6538_ (.A0(net1047),
    .A1(\current_src_addr[1][21] ),
    .S(net1269),
    .X(_1394_));
 sky130_fd_sc_hd__mux2_2 _6539_ (.A0(net1048),
    .A1(\current_src_addr[1][22] ),
    .S(net1269),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_2 _6540_ (.A0(net1049),
    .A1(\current_src_addr[1][23] ),
    .S(net1269),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_2 _6541_ (.A0(net1050),
    .A1(\current_src_addr[1][24] ),
    .S(net1269),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_2 _6542_ (.A0(net1051),
    .A1(\current_src_addr[1][25] ),
    .S(net1269),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_2 _6543_ (.A0(net1052),
    .A1(\current_src_addr[1][26] ),
    .S(net1269),
    .X(_1399_));
 sky130_fd_sc_hd__mux2_2 _6544_ (.A0(net1053),
    .A1(\current_src_addr[1][27] ),
    .S(net1269),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_2 _6545_ (.A0(net1054),
    .A1(\current_src_addr[0][5] ),
    .S(net1252),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_2 _6546_ (.A0(net1055),
    .A1(\current_src_addr[1][28] ),
    .S(net1269),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_2 _6547_ (.A0(net1056),
    .A1(\current_src_addr[1][29] ),
    .S(net1269),
    .X(_1403_));
 sky130_fd_sc_hd__mux2_2 _6548_ (.A0(net1057),
    .A1(\current_src_addr[1][30] ),
    .S(net1269),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_2 _6549_ (.A0(net1058),
    .A1(\current_src_addr[1][31] ),
    .S(net1269),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_2 _6550_ (.A0(net1059),
    .A1(\current_src_addr[2][0] ),
    .S(net1254),
    .X(_1406_));
 sky130_fd_sc_hd__mux2_2 _6551_ (.A0(net1060),
    .A1(\current_src_addr[2][1] ),
    .S(net1254),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_2 _6552_ (.A0(net1061),
    .A1(\current_src_addr[2][2] ),
    .S(net1254),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_2 _6553_ (.A0(net1062),
    .A1(\current_src_addr[2][3] ),
    .S(net1254),
    .X(_1409_));
 sky130_fd_sc_hd__mux2_2 _6554_ (.A0(net1063),
    .A1(\current_src_addr[2][4] ),
    .S(net1254),
    .X(_1410_));
 sky130_fd_sc_hd__mux2_2 _6555_ (.A0(net1064),
    .A1(\current_src_addr[2][5] ),
    .S(net1254),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_2 _6556_ (.A0(net1065),
    .A1(\current_src_addr[0][6] ),
    .S(net1252),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_2 _6557_ (.A0(net1066),
    .A1(\current_src_addr[2][6] ),
    .S(net1254),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_2 _6558_ (.A0(net1067),
    .A1(\current_src_addr[2][7] ),
    .S(net1254),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_2 _6559_ (.A0(net1068),
    .A1(\current_src_addr[2][8] ),
    .S(net1254),
    .X(_1415_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input2 (.A(net1497),
    .X(net2));
 sky130_fd_sc_hd__mux2_2 _6561_ (.A0(net1069),
    .A1(\current_src_addr[2][9] ),
    .S(net1254),
    .X(_1416_));
 sky130_fd_sc_hd__mux2_2 _6562_ (.A0(net1070),
    .A1(\current_src_addr[2][10] ),
    .S(net1254),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_2 _6563_ (.A0(net1071),
    .A1(\current_src_addr[2][11] ),
    .S(net1254),
    .X(_1418_));
 sky130_fd_sc_hd__mux2_2 _6564_ (.A0(net1072),
    .A1(\current_src_addr[2][12] ),
    .S(net1254),
    .X(_1419_));
 sky130_fd_sc_hd__mux2_2 _6565_ (.A0(net1073),
    .A1(\current_src_addr[2][13] ),
    .S(net1254),
    .X(_1420_));
 sky130_fd_sc_hd__mux2_2 _6566_ (.A0(net1074),
    .A1(\current_src_addr[2][14] ),
    .S(net1254),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_2 _6567_ (.A0(net1075),
    .A1(\current_src_addr[2][15] ),
    .S(net1254),
    .X(_1422_));
 sky130_fd_sc_hd__mux2_2 _6568_ (.A0(net1076),
    .A1(\current_src_addr[0][7] ),
    .S(net1252),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_2 _6569_ (.A0(net1077),
    .A1(\current_src_addr[2][16] ),
    .S(net1254),
    .X(_1424_));
 sky130_fd_sc_hd__mux2_2 _6570_ (.A0(net1078),
    .A1(\current_src_addr[2][17] ),
    .S(net1254),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_2 _6571_ (.A0(net1079),
    .A1(\current_src_addr[2][18] ),
    .S(net1254),
    .X(_1426_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input1 (.A(net1374),
    .X(net1));
 sky130_fd_sc_hd__mux2_2 _6573_ (.A0(net1080),
    .A1(\current_src_addr[2][19] ),
    .S(net1254),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_2 _6574_ (.A0(net1081),
    .A1(\current_src_addr[2][20] ),
    .S(net1254),
    .X(_1428_));
 sky130_fd_sc_hd__mux2_2 _6575_ (.A0(net1082),
    .A1(\current_src_addr[2][21] ),
    .S(net1254),
    .X(_1429_));
 sky130_fd_sc_hd__mux2_2 _6576_ (.A0(net1083),
    .A1(\current_src_addr[2][22] ),
    .S(net1254),
    .X(_1430_));
 sky130_fd_sc_hd__mux2_2 _6577_ (.A0(net1084),
    .A1(\current_src_addr[2][23] ),
    .S(net1254),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_2 _6578_ (.A0(net1085),
    .A1(\current_src_addr[2][24] ),
    .S(net1254),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_2 _6579_ (.A0(net1086),
    .A1(\current_src_addr[2][25] ),
    .S(net1254),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_2 _6580_ (.A0(net1087),
    .A1(\current_src_addr[0][8] ),
    .S(net1252),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_2 _6581_ (.A0(net1088),
    .A1(\current_src_addr[2][26] ),
    .S(net1254),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_2 _6582_ (.A0(net1089),
    .A1(\current_src_addr[2][27] ),
    .S(net1254),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_2 _6583_ (.A0(net1090),
    .A1(\current_src_addr[2][28] ),
    .S(net1254),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_2 _6584_ (.A0(net1091),
    .A1(\current_src_addr[2][29] ),
    .S(net1254),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_2 _6585_ (.A0(net1092),
    .A1(\current_src_addr[2][30] ),
    .S(net1254),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_2 _6586_ (.A0(net1093),
    .A1(\current_src_addr[2][31] ),
    .S(net1254),
    .X(_1440_));
 sky130_fd_sc_hd__mux2_2 _6587_ (.A0(net1094),
    .A1(\current_src_addr[3][0] ),
    .S(net1253),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_2 _6588_ (.A0(net1095),
    .A1(\current_src_addr[3][1] ),
    .S(net1253),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_2 _6589_ (.A0(net1096),
    .A1(\current_src_addr[3][2] ),
    .S(net1253),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_2 _6590_ (.A0(net1097),
    .A1(\current_src_addr[3][3] ),
    .S(net1253),
    .X(_1444_));
 sky130_fd_sc_hd__mux2_2 _6591_ (.A0(net1098),
    .A1(\current_src_addr[0][9] ),
    .S(net1252),
    .X(_1445_));
 sky130_fd_sc_hd__inv_1 _6592_ (.A(net534),
    .Y(_3415_));
 sky130_fd_sc_hd__nand3_1 _6593_ (.A(_3312_),
    .B(net557),
    .C(_3415_),
    .Y(_3416_));
 sky130_fd_sc_hd__a21oi_1 _6594_ (.A1(_1458_),
    .A2(_3416_),
    .B1(net558),
    .Y(_1446_));
 sky130_fd_sc_hd__nor3_1 _6595_ (.A(net1273),
    .B(_3301_),
    .C(net535),
    .Y(_3417_));
 sky130_fd_sc_hd__a21oi_1 _6596_ (.A1(net1273),
    .A2(_3301_),
    .B1(_3417_),
    .Y(_3418_));
 sky130_fd_sc_hd__nor2_1 _6597_ (.A(net1271),
    .B(_3418_),
    .Y(_1447_));
 sky130_fd_sc_hd__nor2_1 _6598_ (.A(net562),
    .B(net536),
    .Y(_3419_));
 sky130_fd_sc_hd__mux2i_1 _6599_ (.A0(net562),
    .A1(_3419_),
    .S(net563),
    .Y(_3420_));
 sky130_fd_sc_hd__nor2_1 _6600_ (.A(net564),
    .B(_3420_),
    .Y(_1448_));
 sky130_fd_sc_hd__nor2_1 _6601_ (.A(net565),
    .B(net537),
    .Y(_3421_));
 sky130_fd_sc_hd__mux2i_1 _6602_ (.A0(net565),
    .A1(_3421_),
    .S(net555),
    .Y(_3422_));
 sky130_fd_sc_hd__nor2_1 _6603_ (.A(net556),
    .B(_3422_),
    .Y(_1449_));
 sky130_fd_sc_hd__ha_1 _6604_ (.A(\current_dst_addr[3][2] ),
    .B(\current_dst_addr[3][3] ),
    .COUT(_0381_),
    .SUM(_0382_));
 sky130_fd_sc_hd__ha_1 _6605_ (.A(\current_dst_addr[2][2] ),
    .B(\current_dst_addr[2][3] ),
    .COUT(_0383_),
    .SUM(_0384_));
 sky130_fd_sc_hd__ha_1 _6606_ (.A(\current_dst_addr[1][2] ),
    .B(\current_dst_addr[1][3] ),
    .COUT(_0385_),
    .SUM(_0386_));
 sky130_fd_sc_hd__ha_1 _6607_ (.A(\current_dst_addr[0][2] ),
    .B(\current_dst_addr[0][3] ),
    .COUT(_0387_),
    .SUM(_0388_));
 sky130_fd_sc_hd__ha_1 _6608_ (.A(\current_src_addr[3][2] ),
    .B(\current_src_addr[3][3] ),
    .COUT(_0389_),
    .SUM(_0390_));
 sky130_fd_sc_hd__ha_1 _6609_ (.A(\current_src_addr[2][2] ),
    .B(\current_src_addr[2][3] ),
    .COUT(_0391_),
    .SUM(_0392_));
 sky130_fd_sc_hd__ha_1 _6610_ (.A(\current_src_addr[1][2] ),
    .B(\current_src_addr[1][3] ),
    .COUT(_0393_),
    .SUM(_0394_));
 sky130_fd_sc_hd__ha_1 _6611_ (.A(\current_src_addr[0][2] ),
    .B(\current_src_addr[0][3] ),
    .COUT(_0395_),
    .SUM(_0396_));
 sky130_fd_sc_hd__ha_1 _6612_ (.A(net690),
    .B(net691),
    .COUT(_0397_),
    .SUM(_0398_));
 sky130_fd_sc_hd__ha_1 _6613_ (.A(net655),
    .B(net656),
    .COUT(_0399_),
    .SUM(_0400_));
 sky130_fd_sc_hd__ha_1 _6614_ (.A(net620),
    .B(net621),
    .COUT(_0401_),
    .SUM(_0402_));
 sky130_fd_sc_hd__ha_1 _6615_ (.A(net567),
    .B(net606),
    .COUT(_0403_),
    .SUM(_0404_));
 sky130_fd_sc_hd__ha_1 _6616_ (.A(_0405_),
    .B(_0406_),
    .COUT(_0407_),
    .SUM(_0408_));
 sky130_fd_sc_hd__ha_1 _6617_ (.A(\active_channel_count[0] ),
    .B(\active_channel_count[1] ),
    .COUT(_0409_),
    .SUM(_3443_));
 sky130_fd_sc_hd__ha_1 _6618_ (.A(_0410_),
    .B(_0411_),
    .COUT(_0412_),
    .SUM(_0413_));
 sky130_fd_sc_hd__ha_1 _6619_ (.A(_0414_),
    .B(_0415_),
    .COUT(_0416_),
    .SUM(_0417_));
 sky130_fd_sc_hd__ha_1 _6620_ (.A(_0418_),
    .B(_0419_),
    .COUT(_0420_),
    .SUM(_0421_));
 sky130_fd_sc_hd__ha_1 _6621_ (.A(_0422_),
    .B(_0423_),
    .COUT(_0424_),
    .SUM(_0425_));
 sky130_fd_sc_hd__ha_1 _6622_ (.A(_0426_),
    .B(_0427_),
    .COUT(_0428_),
    .SUM(_0429_));
 sky130_fd_sc_hd__ha_1 _6623_ (.A(_0430_),
    .B(_0431_),
    .COUT(_0432_),
    .SUM(_0433_));
 sky130_fd_sc_hd__ha_1 _6624_ (.A(_0434_),
    .B(_0435_),
    .COUT(_0436_),
    .SUM(_0437_));
 sky130_fd_sc_hd__ha_1 _6625_ (.A(_0438_),
    .B(_0439_),
    .COUT(_0440_),
    .SUM(_0441_));
 sky130_fd_sc_hd__ha_1 _6626_ (.A(_0442_),
    .B(_0443_),
    .COUT(_0444_),
    .SUM(_0445_));
 sky130_fd_sc_hd__ha_1 _6627_ (.A(_0446_),
    .B(_0447_),
    .COUT(_0448_),
    .SUM(_0449_));
 sky130_fd_sc_hd__ha_1 _6628_ (.A(_0450_),
    .B(_0451_),
    .COUT(_0452_),
    .SUM(_0453_));
 sky130_fd_sc_hd__ha_1 _6629_ (.A(_0454_),
    .B(_0455_),
    .COUT(_0456_),
    .SUM(_0457_));
 sky130_fd_sc_hd__ha_1 _6630_ (.A(_0458_),
    .B(_0459_),
    .COUT(_0460_),
    .SUM(_0461_));
 sky130_fd_sc_hd__ha_1 _6631_ (.A(_0462_),
    .B(_0463_),
    .COUT(_0464_),
    .SUM(_0465_));
 sky130_fd_sc_hd__ha_1 _6632_ (.A(_0466_),
    .B(_0467_),
    .COUT(_0468_),
    .SUM(_0469_));
 sky130_fd_sc_hd__ha_1 _6633_ (.A(_0470_),
    .B(_0471_),
    .COUT(_0472_),
    .SUM(_0473_));
 sky130_fd_sc_hd__ha_1 _6634_ (.A(_0474_),
    .B(_0475_),
    .COUT(_0476_),
    .SUM(_0477_));
 sky130_fd_sc_hd__ha_1 _6635_ (.A(_0478_),
    .B(_0479_),
    .COUT(_0480_),
    .SUM(_0481_));
 sky130_fd_sc_hd__ha_1 _6636_ (.A(_0482_),
    .B(_0483_),
    .COUT(_0484_),
    .SUM(_0485_));
 sky130_fd_sc_hd__ha_1 _6637_ (.A(_0486_),
    .B(_0487_),
    .COUT(_0488_),
    .SUM(_0489_));
 sky130_fd_sc_hd__ha_1 _6638_ (.A(_0490_),
    .B(_0491_),
    .COUT(_0492_),
    .SUM(_0493_));
 sky130_fd_sc_hd__ha_1 _6639_ (.A(_0494_),
    .B(_0495_),
    .COUT(_0496_),
    .SUM(_0497_));
 sky130_fd_sc_hd__ha_1 _6640_ (.A(_0498_),
    .B(_0499_),
    .COUT(_0500_),
    .SUM(_0501_));
 sky130_fd_sc_hd__ha_1 _6641_ (.A(_0502_),
    .B(_0503_),
    .COUT(_0504_),
    .SUM(_0505_));
 sky130_fd_sc_hd__ha_1 _6642_ (.A(_0506_),
    .B(_0507_),
    .COUT(_0508_),
    .SUM(_0509_));
 sky130_fd_sc_hd__ha_1 _6643_ (.A(_0510_),
    .B(_0511_),
    .COUT(_0512_),
    .SUM(_0513_));
 sky130_fd_sc_hd__ha_1 _6644_ (.A(_0514_),
    .B(_0515_),
    .COUT(_0516_),
    .SUM(_0517_));
 sky130_fd_sc_hd__ha_1 _6645_ (.A(_0518_),
    .B(_0519_),
    .COUT(_0520_),
    .SUM(_0521_));
 sky130_fd_sc_hd__ha_1 _6646_ (.A(_0522_),
    .B(_0523_),
    .COUT(_0524_),
    .SUM(_0525_));
 sky130_fd_sc_hd__ha_1 _6647_ (.A(_0526_),
    .B(_0527_),
    .COUT(_0528_),
    .SUM(_0529_));
 sky130_fd_sc_hd__ha_1 _6648_ (.A(_0530_),
    .B(_0404_),
    .COUT(_0531_),
    .SUM(_0532_));
 sky130_fd_sc_hd__ha_1 _6649_ (.A(net133),
    .B(net567),
    .COUT(_0533_),
    .SUM(_0534_));
 sky130_fd_sc_hd__ha_1 _6650_ (.A(net186),
    .B(net620),
    .COUT(_0535_),
    .SUM(_0536_));
 sky130_fd_sc_hd__ha_1 _6651_ (.A(_0537_),
    .B(_0402_),
    .COUT(_0538_),
    .SUM(_0539_));
 sky130_fd_sc_hd__ha_1 _6652_ (.A(_0540_),
    .B(_0541_),
    .COUT(_0542_),
    .SUM(_0543_));
 sky130_fd_sc_hd__ha_1 _6653_ (.A(_0544_),
    .B(_0545_),
    .COUT(_0546_),
    .SUM(_0547_));
 sky130_fd_sc_hd__ha_1 _6654_ (.A(_0548_),
    .B(_0549_),
    .COUT(_0550_),
    .SUM(_0551_));
 sky130_fd_sc_hd__ha_1 _6655_ (.A(_0552_),
    .B(_0553_),
    .COUT(_0554_),
    .SUM(_0555_));
 sky130_fd_sc_hd__ha_1 _6656_ (.A(_0556_),
    .B(_0557_),
    .COUT(_0558_),
    .SUM(_0559_));
 sky130_fd_sc_hd__ha_1 _6657_ (.A(_0560_),
    .B(_0561_),
    .COUT(_0562_),
    .SUM(_0563_));
 sky130_fd_sc_hd__ha_1 _6658_ (.A(_0564_),
    .B(_0565_),
    .COUT(_0566_),
    .SUM(_0567_));
 sky130_fd_sc_hd__ha_1 _6659_ (.A(_0568_),
    .B(_0569_),
    .COUT(_0570_),
    .SUM(_0571_));
 sky130_fd_sc_hd__ha_1 _6660_ (.A(_0572_),
    .B(_0573_),
    .COUT(_0574_),
    .SUM(_0575_));
 sky130_fd_sc_hd__ha_1 _6661_ (.A(_0576_),
    .B(_0577_),
    .COUT(_0578_),
    .SUM(_0579_));
 sky130_fd_sc_hd__ha_1 _6662_ (.A(_0580_),
    .B(_0581_),
    .COUT(_0582_),
    .SUM(_0583_));
 sky130_fd_sc_hd__ha_1 _6663_ (.A(_0584_),
    .B(_0585_),
    .COUT(_0586_),
    .SUM(_0587_));
 sky130_fd_sc_hd__ha_1 _6664_ (.A(_0588_),
    .B(_0589_),
    .COUT(_0590_),
    .SUM(_0591_));
 sky130_fd_sc_hd__ha_1 _6665_ (.A(_0592_),
    .B(_0593_),
    .COUT(_0594_),
    .SUM(_0595_));
 sky130_fd_sc_hd__ha_1 _6666_ (.A(_0596_),
    .B(_0597_),
    .COUT(_0598_),
    .SUM(_0599_));
 sky130_fd_sc_hd__ha_1 _6667_ (.A(_0600_),
    .B(_0601_),
    .COUT(_0602_),
    .SUM(_0603_));
 sky130_fd_sc_hd__ha_1 _6668_ (.A(_0604_),
    .B(_0605_),
    .COUT(_0606_),
    .SUM(_0607_));
 sky130_fd_sc_hd__ha_1 _6669_ (.A(_0608_),
    .B(_0609_),
    .COUT(_0610_),
    .SUM(_0611_));
 sky130_fd_sc_hd__ha_1 _6670_ (.A(_0612_),
    .B(_0613_),
    .COUT(_0614_),
    .SUM(_0615_));
 sky130_fd_sc_hd__ha_1 _6671_ (.A(_0616_),
    .B(_0617_),
    .COUT(_0618_),
    .SUM(_0619_));
 sky130_fd_sc_hd__ha_1 _6672_ (.A(_0620_),
    .B(_0621_),
    .COUT(_0622_),
    .SUM(_0623_));
 sky130_fd_sc_hd__ha_1 _6673_ (.A(_0624_),
    .B(_0625_),
    .COUT(_0626_),
    .SUM(_0627_));
 sky130_fd_sc_hd__ha_1 _6674_ (.A(_0628_),
    .B(_0629_),
    .COUT(_0630_),
    .SUM(_0631_));
 sky130_fd_sc_hd__ha_1 _6675_ (.A(_0632_),
    .B(_0633_),
    .COUT(_0634_),
    .SUM(_0635_));
 sky130_fd_sc_hd__ha_1 _6676_ (.A(_0636_),
    .B(_0637_),
    .COUT(_0638_),
    .SUM(_0639_));
 sky130_fd_sc_hd__ha_1 _6677_ (.A(_0640_),
    .B(_0641_),
    .COUT(_0642_),
    .SUM(_0643_));
 sky130_fd_sc_hd__ha_1 _6678_ (.A(_0644_),
    .B(_0645_),
    .COUT(_0646_),
    .SUM(_0647_));
 sky130_fd_sc_hd__ha_1 _6679_ (.A(_0648_),
    .B(_0649_),
    .COUT(_0650_),
    .SUM(_0651_));
 sky130_fd_sc_hd__ha_1 _6680_ (.A(_0652_),
    .B(_0653_),
    .COUT(_0654_),
    .SUM(_0655_));
 sky130_fd_sc_hd__ha_1 _6681_ (.A(_0656_),
    .B(_0657_),
    .COUT(_0658_),
    .SUM(_0659_));
 sky130_fd_sc_hd__ha_1 _6682_ (.A(net256),
    .B(net690),
    .COUT(_0660_),
    .SUM(_0661_));
 sky130_fd_sc_hd__ha_1 _6683_ (.A(_0662_),
    .B(_0398_),
    .COUT(_0663_),
    .SUM(_0664_));
 sky130_fd_sc_hd__ha_1 _6684_ (.A(_0665_),
    .B(_0666_),
    .COUT(_0667_),
    .SUM(_0668_));
 sky130_fd_sc_hd__ha_1 _6685_ (.A(_0669_),
    .B(_0670_),
    .COUT(_0671_),
    .SUM(_0672_));
 sky130_fd_sc_hd__ha_1 _6686_ (.A(_0673_),
    .B(_0674_),
    .COUT(_0675_),
    .SUM(_0676_));
 sky130_fd_sc_hd__ha_1 _6687_ (.A(_0677_),
    .B(_0678_),
    .COUT(_0679_),
    .SUM(_0680_));
 sky130_fd_sc_hd__ha_1 _6688_ (.A(_0681_),
    .B(_0682_),
    .COUT(_0683_),
    .SUM(_0684_));
 sky130_fd_sc_hd__ha_1 _6689_ (.A(_0685_),
    .B(_0686_),
    .COUT(_0687_),
    .SUM(_0688_));
 sky130_fd_sc_hd__ha_1 _6690_ (.A(_0689_),
    .B(_0690_),
    .COUT(_0691_),
    .SUM(_0692_));
 sky130_fd_sc_hd__ha_1 _6691_ (.A(_0693_),
    .B(_0694_),
    .COUT(_0695_),
    .SUM(_0696_));
 sky130_fd_sc_hd__ha_1 _6692_ (.A(_0697_),
    .B(_0698_),
    .COUT(_0699_),
    .SUM(_0700_));
 sky130_fd_sc_hd__ha_1 _6693_ (.A(_0701_),
    .B(_0702_),
    .COUT(_0703_),
    .SUM(_0704_));
 sky130_fd_sc_hd__ha_1 _6694_ (.A(_0705_),
    .B(_0706_),
    .COUT(_0707_),
    .SUM(_0708_));
 sky130_fd_sc_hd__ha_1 _6695_ (.A(_0709_),
    .B(_0710_),
    .COUT(_0711_),
    .SUM(_0712_));
 sky130_fd_sc_hd__ha_1 _6696_ (.A(_0713_),
    .B(_0714_),
    .COUT(_0715_),
    .SUM(_0716_));
 sky130_fd_sc_hd__ha_1 _6697_ (.A(_0717_),
    .B(_0718_),
    .COUT(_0719_),
    .SUM(_0720_));
 sky130_fd_sc_hd__ha_1 _6698_ (.A(_0721_),
    .B(_0722_),
    .COUT(_0723_),
    .SUM(_0724_));
 sky130_fd_sc_hd__ha_1 _6699_ (.A(_0725_),
    .B(_0726_),
    .COUT(_0727_),
    .SUM(_0728_));
 sky130_fd_sc_hd__ha_1 _6700_ (.A(_0729_),
    .B(_0730_),
    .COUT(_0731_),
    .SUM(_0732_));
 sky130_fd_sc_hd__ha_1 _6701_ (.A(_0733_),
    .B(_0734_),
    .COUT(_0735_),
    .SUM(_0736_));
 sky130_fd_sc_hd__ha_1 _6702_ (.A(_0737_),
    .B(_0738_),
    .COUT(_0739_),
    .SUM(_0740_));
 sky130_fd_sc_hd__ha_1 _6703_ (.A(_0741_),
    .B(_0742_),
    .COUT(_0743_),
    .SUM(_0744_));
 sky130_fd_sc_hd__ha_1 _6704_ (.A(_0745_),
    .B(_0746_),
    .COUT(_0747_),
    .SUM(_0748_));
 sky130_fd_sc_hd__ha_1 _6705_ (.A(_0749_),
    .B(_0750_),
    .COUT(_0751_),
    .SUM(_0752_));
 sky130_fd_sc_hd__ha_1 _6706_ (.A(_0753_),
    .B(_0754_),
    .COUT(_0755_),
    .SUM(_0756_));
 sky130_fd_sc_hd__ha_1 _6707_ (.A(_0757_),
    .B(_0758_),
    .COUT(_0759_),
    .SUM(_0760_));
 sky130_fd_sc_hd__ha_1 _6708_ (.A(_0761_),
    .B(_0762_),
    .COUT(_0763_),
    .SUM(_0764_));
 sky130_fd_sc_hd__ha_1 _6709_ (.A(_0765_),
    .B(_0766_),
    .COUT(_0767_),
    .SUM(_0768_));
 sky130_fd_sc_hd__ha_1 _6710_ (.A(_0769_),
    .B(_0770_),
    .COUT(_0771_),
    .SUM(_0772_));
 sky130_fd_sc_hd__ha_1 _6711_ (.A(_0773_),
    .B(_0774_),
    .COUT(_0775_),
    .SUM(_0776_));
 sky130_fd_sc_hd__ha_1 _6712_ (.A(_0777_),
    .B(_0778_),
    .COUT(_0779_),
    .SUM(_0780_));
 sky130_fd_sc_hd__ha_1 _6713_ (.A(_0781_),
    .B(_0782_),
    .COUT(_0783_),
    .SUM(_0784_));
 sky130_fd_sc_hd__ha_1 _6714_ (.A(net221),
    .B(net655),
    .COUT(_0785_),
    .SUM(_0786_));
 sky130_fd_sc_hd__ha_1 _6715_ (.A(_0787_),
    .B(_0400_),
    .COUT(_0788_),
    .SUM(_0789_));
 sky130_fd_sc_hd__ha_1 _6716_ (.A(_0790_),
    .B(_0791_),
    .COUT(_0792_),
    .SUM(_0793_));
 sky130_fd_sc_hd__ha_1 _6717_ (.A(_0794_),
    .B(_0795_),
    .COUT(_0796_),
    .SUM(_0797_));
 sky130_fd_sc_hd__ha_1 _6718_ (.A(_0798_),
    .B(_0799_),
    .COUT(_0800_),
    .SUM(_0801_));
 sky130_fd_sc_hd__ha_1 _6719_ (.A(_0802_),
    .B(_0803_),
    .COUT(_0804_),
    .SUM(_0805_));
 sky130_fd_sc_hd__ha_1 _6720_ (.A(_0806_),
    .B(_0807_),
    .COUT(_0808_),
    .SUM(_0809_));
 sky130_fd_sc_hd__ha_1 _6721_ (.A(_0810_),
    .B(_0811_),
    .COUT(_0812_),
    .SUM(_0813_));
 sky130_fd_sc_hd__ha_1 _6722_ (.A(_0814_),
    .B(_0815_),
    .COUT(_0816_),
    .SUM(_0817_));
 sky130_fd_sc_hd__ha_1 _6723_ (.A(_0818_),
    .B(_0819_),
    .COUT(_0820_),
    .SUM(_0821_));
 sky130_fd_sc_hd__ha_1 _6724_ (.A(_0822_),
    .B(_0823_),
    .COUT(_0824_),
    .SUM(_0825_));
 sky130_fd_sc_hd__ha_1 _6725_ (.A(_0826_),
    .B(_0827_),
    .COUT(_0828_),
    .SUM(_0829_));
 sky130_fd_sc_hd__ha_1 _6726_ (.A(_0830_),
    .B(_0831_),
    .COUT(_0832_),
    .SUM(_0833_));
 sky130_fd_sc_hd__ha_1 _6727_ (.A(_0834_),
    .B(_0835_),
    .COUT(_0836_),
    .SUM(_0837_));
 sky130_fd_sc_hd__ha_1 _6728_ (.A(_0838_),
    .B(_0839_),
    .COUT(_0840_),
    .SUM(_0841_));
 sky130_fd_sc_hd__ha_1 _6729_ (.A(_0842_),
    .B(_0843_),
    .COUT(_0844_),
    .SUM(_0845_));
 sky130_fd_sc_hd__ha_1 _6730_ (.A(_0846_),
    .B(_0847_),
    .COUT(_0848_),
    .SUM(_0849_));
 sky130_fd_sc_hd__ha_1 _6731_ (.A(_0850_),
    .B(_0851_),
    .COUT(_0852_),
    .SUM(_0853_));
 sky130_fd_sc_hd__ha_1 _6732_ (.A(_0854_),
    .B(_0855_),
    .COUT(_0856_),
    .SUM(_0857_));
 sky130_fd_sc_hd__ha_1 _6733_ (.A(_0858_),
    .B(_0859_),
    .COUT(_0860_),
    .SUM(_0861_));
 sky130_fd_sc_hd__ha_1 _6734_ (.A(_0862_),
    .B(_0863_),
    .COUT(_0864_),
    .SUM(_0865_));
 sky130_fd_sc_hd__ha_1 _6735_ (.A(_0866_),
    .B(_0867_),
    .COUT(_0868_),
    .SUM(_0869_));
 sky130_fd_sc_hd__ha_1 _6736_ (.A(_0870_),
    .B(_0871_),
    .COUT(_0872_),
    .SUM(_0873_));
 sky130_fd_sc_hd__ha_1 _6737_ (.A(_0874_),
    .B(_0875_),
    .COUT(_0876_),
    .SUM(_0877_));
 sky130_fd_sc_hd__ha_1 _6738_ (.A(_0878_),
    .B(_0879_),
    .COUT(_0880_),
    .SUM(_0881_));
 sky130_fd_sc_hd__ha_1 _6739_ (.A(_0882_),
    .B(_0883_),
    .COUT(_0884_),
    .SUM(_0885_));
 sky130_fd_sc_hd__ha_1 _6740_ (.A(_0886_),
    .B(_0887_),
    .COUT(_0888_),
    .SUM(_0889_));
 sky130_fd_sc_hd__ha_1 _6741_ (.A(_0890_),
    .B(_0891_),
    .COUT(_0892_),
    .SUM(_0893_));
 sky130_fd_sc_hd__ha_1 _6742_ (.A(_0894_),
    .B(_0895_),
    .COUT(_0896_),
    .SUM(_0897_));
 sky130_fd_sc_hd__ha_1 _6743_ (.A(_0898_),
    .B(_0899_),
    .COUT(_0900_),
    .SUM(_0901_));
 sky130_fd_sc_hd__ha_1 _6744_ (.A(_0902_),
    .B(_0903_),
    .COUT(_0904_),
    .SUM(_0905_));
 sky130_fd_sc_hd__ha_1 _6745_ (.A(_0906_),
    .B(_0907_),
    .COUT(_0908_),
    .SUM(_0909_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_4 place1274 (.A(net405),
    .X(net1274));
 sky130_fd_sc_hd__buf_4 place1271 (.A(net561),
    .X(net1271));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[0]$_DFF_PN0_  (.D(_0000_),
    .Q(\active_channel_count[0] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[1]$_DFF_PN0_  (.D(_0001_),
    .Q(\active_channel_count[1] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[2]$_DFF_PN0_  (.D(_0002_),
    .Q(\active_channel_count[2] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \active_channel_count[3]$_DFF_PN0_  (.D(_0003_),
    .Q(\active_channel_count[3] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[0]$_DFF_PN0_  (.D(_0004_),
    .Q(net538),
    .RESET_B(net1279),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[1]$_DFF_PN0_  (.D(_0005_),
    .Q(net539),
    .RESET_B(net1290),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[2]$_DFF_PN0_  (.D(_0006_),
    .Q(net540),
    .RESET_B(net1275),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_busy[3]$_DFF_PN0_  (.D(_0007_),
    .Q(net541),
    .RESET_B(net1283),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[0]$_DFF_PN0_  (.D(_3428_),
    .Q(net542),
    .RESET_B(net1279),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[1]$_DFF_PN0_  (.D(_3426_),
    .Q(net543),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[2]$_DFF_PN0_  (.D(_3423_),
    .Q(net544),
    .RESET_B(net1275),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_done[3]$_DFF_PN0_  (.D(_3425_),
    .Q(net545),
    .RESET_B(net1283),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[0]$_DFF_PN0_  (.D(_0008_),
    .Q(net546),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[1]$_DFF_PN0_  (.D(_0009_),
    .Q(net547),
    .RESET_B(net1290),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[2]$_DFF_PN0_  (.D(_0010_),
    .Q(net548),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_error[3]$_DFF_PN0_  (.D(_0011_),
    .Q(net549),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[0][0]$_DFF_PN0_  (.D(_3440_),
    .Q(net554),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[0][1]$_DFF_PN0_  (.D(_3441_),
    .Q(net557),
    .RESET_B(net1279),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[0][2]$_DFF_PN0_  (.D(_3442_),
    .Q(net558),
    .RESET_B(net1279),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[1][0]$_DFF_PN0_  (.D(_3437_),
    .Q(net559),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[1][1]$_DFF_PN0_  (.D(_3438_),
    .Q(net560),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[1][2]$_DFF_PN0_  (.D(_3439_),
    .Q(net561),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[2][0]$_DFF_PN0_  (.D(_3434_),
    .Q(net562),
    .RESET_B(net1276),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[2][1]$_DFF_PN0_  (.D(_3435_),
    .Q(net563),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[2][2]$_DFF_PN0_  (.D(_3436_),
    .Q(net564),
    .RESET_B(net1275),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[3][0]$_DFF_PN0_  (.D(_3431_),
    .Q(net565),
    .RESET_B(net1283),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[3][1]$_DFF_PN0_  (.D(_3432_),
    .Q(net555),
    .RESET_B(net1283),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \channel_state[3][2]$_DFF_PN0_  (.D(_3433_),
    .Q(net556),
    .RESET_B(net1283),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][0]$_DFFE_PN0P_  (.D(_0910_),
    .Q(\current_dst_addr[0][0] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][10]$_DFF_PN0_  (.D(_0012_),
    .Q(\current_dst_addr[0][10] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][11]$_DFF_PN0_  (.D(_0013_),
    .Q(\current_dst_addr[0][11] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][12]$_DFF_PN0_  (.D(_0014_),
    .Q(\current_dst_addr[0][12] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][13]$_DFF_PN0_  (.D(_0015_),
    .Q(\current_dst_addr[0][13] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][14]$_DFF_PN0_  (.D(_0016_),
    .Q(\current_dst_addr[0][14] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][15]$_DFF_PN0_  (.D(_0017_),
    .Q(\current_dst_addr[0][15] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][16]$_DFF_PN0_  (.D(_0018_),
    .Q(\current_dst_addr[0][16] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][17]$_DFF_PN0_  (.D(_0019_),
    .Q(\current_dst_addr[0][17] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][18]$_DFF_PN0_  (.D(_0020_),
    .Q(\current_dst_addr[0][18] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][19]$_DFF_PN0_  (.D(_0021_),
    .Q(\current_dst_addr[0][19] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][1]$_DFFE_PN0P_  (.D(_0911_),
    .Q(\current_dst_addr[0][1] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][20]$_DFF_PN0_  (.D(_0022_),
    .Q(\current_dst_addr[0][20] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][21]$_DFF_PN0_  (.D(_0023_),
    .Q(\current_dst_addr[0][21] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][22]$_DFF_PN0_  (.D(_0024_),
    .Q(\current_dst_addr[0][22] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][23]$_DFF_PN0_  (.D(_0025_),
    .Q(\current_dst_addr[0][23] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][24]$_DFF_PN0_  (.D(_0026_),
    .Q(\current_dst_addr[0][24] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][25]$_DFF_PN0_  (.D(_0027_),
    .Q(\current_dst_addr[0][25] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][26]$_DFF_PN0_  (.D(_0028_),
    .Q(\current_dst_addr[0][26] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][27]$_DFF_PN0_  (.D(_0029_),
    .Q(\current_dst_addr[0][27] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][28]$_DFF_PN0_  (.D(_0030_),
    .Q(\current_dst_addr[0][28] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][29]$_DFF_PN0_  (.D(_0031_),
    .Q(\current_dst_addr[0][29] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][2]$_DFF_PN0_  (.D(_0032_),
    .Q(\current_dst_addr[0][2] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][30]$_DFF_PN0_  (.D(_0033_),
    .Q(\current_dst_addr[0][30] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][31]$_DFF_PN0_  (.D(_0034_),
    .Q(\current_dst_addr[0][31] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][3]$_DFF_PN0_  (.D(_0035_),
    .Q(\current_dst_addr[0][3] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][4]$_DFF_PN0_  (.D(_0036_),
    .Q(\current_dst_addr[0][4] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][5]$_DFF_PN0_  (.D(_0037_),
    .Q(\current_dst_addr[0][5] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][6]$_DFF_PN0_  (.D(_0038_),
    .Q(\current_dst_addr[0][6] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][7]$_DFF_PN0_  (.D(_0039_),
    .Q(\current_dst_addr[0][7] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][8]$_DFF_PN0_  (.D(_0040_),
    .Q(\current_dst_addr[0][8] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[0][9]$_DFF_PN0_  (.D(_0041_),
    .Q(\current_dst_addr[0][9] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][0]$_DFFE_PN0P_  (.D(_0912_),
    .Q(\current_dst_addr[1][0] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][10]$_DFF_PN0_  (.D(_0042_),
    .Q(\current_dst_addr[1][10] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][11]$_DFF_PN0_  (.D(_0043_),
    .Q(\current_dst_addr[1][11] ),
    .RESET_B(net1290),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][12]$_DFF_PN0_  (.D(_0044_),
    .Q(\current_dst_addr[1][12] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][13]$_DFF_PN0_  (.D(_0045_),
    .Q(\current_dst_addr[1][13] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][14]$_DFF_PN0_  (.D(_0046_),
    .Q(\current_dst_addr[1][14] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][15]$_DFF_PN0_  (.D(_0047_),
    .Q(\current_dst_addr[1][15] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][16]$_DFF_PN0_  (.D(_0048_),
    .Q(\current_dst_addr[1][16] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][17]$_DFF_PN0_  (.D(_0049_),
    .Q(\current_dst_addr[1][17] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][18]$_DFF_PN0_  (.D(_0050_),
    .Q(\current_dst_addr[1][18] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][19]$_DFF_PN0_  (.D(_0051_),
    .Q(\current_dst_addr[1][19] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][1]$_DFFE_PN0P_  (.D(_0913_),
    .Q(\current_dst_addr[1][1] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][20]$_DFF_PN0_  (.D(_0052_),
    .Q(\current_dst_addr[1][20] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][21]$_DFF_PN0_  (.D(_0053_),
    .Q(\current_dst_addr[1][21] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][22]$_DFF_PN0_  (.D(_0054_),
    .Q(\current_dst_addr[1][22] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][23]$_DFF_PN0_  (.D(_0055_),
    .Q(\current_dst_addr[1][23] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][24]$_DFF_PN0_  (.D(_0056_),
    .Q(\current_dst_addr[1][24] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][25]$_DFF_PN0_  (.D(_0057_),
    .Q(\current_dst_addr[1][25] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][26]$_DFF_PN0_  (.D(_0058_),
    .Q(\current_dst_addr[1][26] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][27]$_DFF_PN0_  (.D(_0059_),
    .Q(\current_dst_addr[1][27] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][28]$_DFF_PN0_  (.D(_0060_),
    .Q(\current_dst_addr[1][28] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][29]$_DFF_PN0_  (.D(_0061_),
    .Q(\current_dst_addr[1][29] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][2]$_DFF_PN0_  (.D(_0062_),
    .Q(\current_dst_addr[1][2] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][30]$_DFF_PN0_  (.D(_0063_),
    .Q(\current_dst_addr[1][30] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][31]$_DFF_PN0_  (.D(_0064_),
    .Q(\current_dst_addr[1][31] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][3]$_DFF_PN0_  (.D(_0065_),
    .Q(\current_dst_addr[1][3] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][4]$_DFF_PN0_  (.D(_0066_),
    .Q(\current_dst_addr[1][4] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][5]$_DFF_PN0_  (.D(_0067_),
    .Q(\current_dst_addr[1][5] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][6]$_DFF_PN0_  (.D(_0068_),
    .Q(\current_dst_addr[1][6] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][7]$_DFF_PN0_  (.D(_0069_),
    .Q(\current_dst_addr[1][7] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][8]$_DFF_PN0_  (.D(_0070_),
    .Q(\current_dst_addr[1][8] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[1][9]$_DFF_PN0_  (.D(_0071_),
    .Q(\current_dst_addr[1][9] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][0]$_DFFE_PN0P_  (.D(_0914_),
    .Q(\current_dst_addr[2][0] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][10]$_DFF_PN0_  (.D(_0072_),
    .Q(\current_dst_addr[2][10] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][11]$_DFF_PN0_  (.D(_0073_),
    .Q(\current_dst_addr[2][11] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][12]$_DFF_PN0_  (.D(_0074_),
    .Q(\current_dst_addr[2][12] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][13]$_DFF_PN0_  (.D(_0075_),
    .Q(\current_dst_addr[2][13] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][14]$_DFF_PN0_  (.D(_0076_),
    .Q(\current_dst_addr[2][14] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][15]$_DFF_PN0_  (.D(_0077_),
    .Q(\current_dst_addr[2][15] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][16]$_DFF_PN0_  (.D(_0078_),
    .Q(\current_dst_addr[2][16] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][17]$_DFF_PN0_  (.D(_0079_),
    .Q(\current_dst_addr[2][17] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][18]$_DFF_PN0_  (.D(_0080_),
    .Q(\current_dst_addr[2][18] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][19]$_DFF_PN0_  (.D(_0081_),
    .Q(\current_dst_addr[2][19] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][1]$_DFFE_PN0P_  (.D(_0915_),
    .Q(\current_dst_addr[2][1] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][20]$_DFF_PN0_  (.D(_0082_),
    .Q(\current_dst_addr[2][20] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][21]$_DFF_PN0_  (.D(_0083_),
    .Q(\current_dst_addr[2][21] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][22]$_DFF_PN0_  (.D(_0084_),
    .Q(\current_dst_addr[2][22] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][23]$_DFF_PN0_  (.D(_0085_),
    .Q(\current_dst_addr[2][23] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][24]$_DFF_PN0_  (.D(_0086_),
    .Q(\current_dst_addr[2][24] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][25]$_DFF_PN0_  (.D(_0087_),
    .Q(\current_dst_addr[2][25] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][26]$_DFF_PN0_  (.D(_0088_),
    .Q(\current_dst_addr[2][26] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][27]$_DFF_PN0_  (.D(_0089_),
    .Q(\current_dst_addr[2][27] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][28]$_DFF_PN0_  (.D(_0090_),
    .Q(\current_dst_addr[2][28] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][29]$_DFF_PN0_  (.D(_0091_),
    .Q(\current_dst_addr[2][29] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][2]$_DFF_PN0_  (.D(_0092_),
    .Q(\current_dst_addr[2][2] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][30]$_DFF_PN0_  (.D(_0093_),
    .Q(\current_dst_addr[2][30] ),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][31]$_DFF_PN0_  (.D(_0094_),
    .Q(\current_dst_addr[2][31] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][3]$_DFF_PN0_  (.D(_0095_),
    .Q(\current_dst_addr[2][3] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][4]$_DFF_PN0_  (.D(_0096_),
    .Q(\current_dst_addr[2][4] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][5]$_DFF_PN0_  (.D(_0097_),
    .Q(\current_dst_addr[2][5] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][6]$_DFF_PN0_  (.D(_0098_),
    .Q(\current_dst_addr[2][6] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][7]$_DFF_PN0_  (.D(_0099_),
    .Q(\current_dst_addr[2][7] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][8]$_DFF_PN0_  (.D(_0100_),
    .Q(\current_dst_addr[2][8] ),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[2][9]$_DFF_PN0_  (.D(_0101_),
    .Q(\current_dst_addr[2][9] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][0]$_DFFE_PN0P_  (.D(_0916_),
    .Q(\current_dst_addr[3][0] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][10]$_DFF_PN0_  (.D(_0102_),
    .Q(\current_dst_addr[3][10] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][11]$_DFF_PN0_  (.D(_0103_),
    .Q(\current_dst_addr[3][11] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][12]$_DFF_PN0_  (.D(_0104_),
    .Q(\current_dst_addr[3][12] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][13]$_DFF_PN0_  (.D(_0105_),
    .Q(\current_dst_addr[3][13] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][14]$_DFF_PN0_  (.D(_0106_),
    .Q(\current_dst_addr[3][14] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][15]$_DFF_PN0_  (.D(_0107_),
    .Q(\current_dst_addr[3][15] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][16]$_DFF_PN0_  (.D(_0108_),
    .Q(\current_dst_addr[3][16] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][17]$_DFF_PN0_  (.D(_0109_),
    .Q(\current_dst_addr[3][17] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][18]$_DFF_PN0_  (.D(_0110_),
    .Q(\current_dst_addr[3][18] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][19]$_DFF_PN0_  (.D(_0111_),
    .Q(\current_dst_addr[3][19] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][1]$_DFFE_PN0P_  (.D(_0917_),
    .Q(\current_dst_addr[3][1] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][20]$_DFF_PN0_  (.D(_0112_),
    .Q(\current_dst_addr[3][20] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][21]$_DFF_PN0_  (.D(_0113_),
    .Q(\current_dst_addr[3][21] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][22]$_DFF_PN0_  (.D(_0114_),
    .Q(\current_dst_addr[3][22] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][23]$_DFF_PN0_  (.D(_0115_),
    .Q(\current_dst_addr[3][23] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][24]$_DFF_PN0_  (.D(_0116_),
    .Q(\current_dst_addr[3][24] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][25]$_DFF_PN0_  (.D(_0117_),
    .Q(\current_dst_addr[3][25] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][26]$_DFF_PN0_  (.D(_0118_),
    .Q(\current_dst_addr[3][26] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][27]$_DFF_PN0_  (.D(_0119_),
    .Q(\current_dst_addr[3][27] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][28]$_DFF_PN0_  (.D(_0120_),
    .Q(\current_dst_addr[3][28] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][29]$_DFF_PN0_  (.D(_0121_),
    .Q(\current_dst_addr[3][29] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][2]$_DFF_PN0_  (.D(_0122_),
    .Q(\current_dst_addr[3][2] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][30]$_DFF_PN0_  (.D(_0123_),
    .Q(\current_dst_addr[3][30] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][31]$_DFF_PN0_  (.D(_0124_),
    .Q(\current_dst_addr[3][31] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][3]$_DFF_PN0_  (.D(_0125_),
    .Q(\current_dst_addr[3][3] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][4]$_DFF_PN0_  (.D(_0126_),
    .Q(\current_dst_addr[3][4] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][5]$_DFF_PN0_  (.D(_0127_),
    .Q(\current_dst_addr[3][5] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][6]$_DFF_PN0_  (.D(_0128_),
    .Q(\current_dst_addr[3][6] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][7]$_DFF_PN0_  (.D(_0129_),
    .Q(\current_dst_addr[3][7] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][8]$_DFF_PN0_  (.D(_0130_),
    .Q(\current_dst_addr[3][8] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_dst_addr[3][9]$_DFF_PN0_  (.D(_0131_),
    .Q(\current_dst_addr[3][9] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][0]$_DFFE_PN0P_  (.D(_0918_),
    .Q(\current_src_addr[0][0] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][10]$_DFF_PN0_  (.D(_0132_),
    .Q(\current_src_addr[0][10] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][11]$_DFF_PN0_  (.D(_0133_),
    .Q(\current_src_addr[0][11] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][12]$_DFF_PN0_  (.D(_0134_),
    .Q(\current_src_addr[0][12] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][13]$_DFF_PN0_  (.D(_0135_),
    .Q(\current_src_addr[0][13] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][14]$_DFF_PN0_  (.D(_0136_),
    .Q(\current_src_addr[0][14] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][15]$_DFF_PN0_  (.D(_0137_),
    .Q(\current_src_addr[0][15] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][16]$_DFF_PN0_  (.D(_0138_),
    .Q(\current_src_addr[0][16] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][17]$_DFF_PN0_  (.D(_0139_),
    .Q(\current_src_addr[0][17] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][18]$_DFF_PN0_  (.D(_0140_),
    .Q(\current_src_addr[0][18] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][19]$_DFF_PN0_  (.D(_0141_),
    .Q(\current_src_addr[0][19] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][1]$_DFFE_PN0P_  (.D(_0919_),
    .Q(\current_src_addr[0][1] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][20]$_DFF_PN0_  (.D(_0142_),
    .Q(\current_src_addr[0][20] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][21]$_DFF_PN0_  (.D(_0143_),
    .Q(\current_src_addr[0][21] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][22]$_DFF_PN0_  (.D(_0144_),
    .Q(\current_src_addr[0][22] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][23]$_DFF_PN0_  (.D(_0145_),
    .Q(\current_src_addr[0][23] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][24]$_DFF_PN0_  (.D(_0146_),
    .Q(\current_src_addr[0][24] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][25]$_DFF_PN0_  (.D(_0147_),
    .Q(\current_src_addr[0][25] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][26]$_DFF_PN0_  (.D(_0148_),
    .Q(\current_src_addr[0][26] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][27]$_DFF_PN0_  (.D(_0149_),
    .Q(\current_src_addr[0][27] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][28]$_DFF_PN0_  (.D(_0150_),
    .Q(\current_src_addr[0][28] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][29]$_DFF_PN0_  (.D(_0151_),
    .Q(\current_src_addr[0][29] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][2]$_DFF_PN0_  (.D(_0152_),
    .Q(\current_src_addr[0][2] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][30]$_DFF_PN0_  (.D(_0153_),
    .Q(\current_src_addr[0][30] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][31]$_DFF_PN0_  (.D(_0154_),
    .Q(\current_src_addr[0][31] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][3]$_DFF_PN0_  (.D(_0155_),
    .Q(\current_src_addr[0][3] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][4]$_DFF_PN0_  (.D(_0156_),
    .Q(\current_src_addr[0][4] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][5]$_DFF_PN0_  (.D(_0157_),
    .Q(\current_src_addr[0][5] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][6]$_DFF_PN0_  (.D(_0158_),
    .Q(\current_src_addr[0][6] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][7]$_DFF_PN0_  (.D(_0159_),
    .Q(\current_src_addr[0][7] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][8]$_DFF_PN0_  (.D(_0160_),
    .Q(\current_src_addr[0][8] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[0][9]$_DFF_PN0_  (.D(_0161_),
    .Q(\current_src_addr[0][9] ),
    .RESET_B(net1279),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][0]$_DFFE_PN0P_  (.D(_0920_),
    .Q(\current_src_addr[1][0] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][10]$_DFF_PN0_  (.D(_0162_),
    .Q(\current_src_addr[1][10] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][11]$_DFF_PN0_  (.D(_0163_),
    .Q(\current_src_addr[1][11] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][12]$_DFF_PN0_  (.D(_0164_),
    .Q(\current_src_addr[1][12] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][13]$_DFF_PN0_  (.D(_0165_),
    .Q(\current_src_addr[1][13] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][14]$_DFF_PN0_  (.D(_0166_),
    .Q(\current_src_addr[1][14] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][15]$_DFF_PN0_  (.D(_0167_),
    .Q(\current_src_addr[1][15] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][16]$_DFF_PN0_  (.D(_0168_),
    .Q(\current_src_addr[1][16] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][17]$_DFF_PN0_  (.D(_0169_),
    .Q(\current_src_addr[1][17] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][18]$_DFF_PN0_  (.D(_0170_),
    .Q(\current_src_addr[1][18] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][19]$_DFF_PN0_  (.D(_0171_),
    .Q(\current_src_addr[1][19] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][1]$_DFFE_PN0P_  (.D(_0921_),
    .Q(\current_src_addr[1][1] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][20]$_DFF_PN0_  (.D(_0172_),
    .Q(\current_src_addr[1][20] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][21]$_DFF_PN0_  (.D(_0173_),
    .Q(\current_src_addr[1][21] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][22]$_DFF_PN0_  (.D(_0174_),
    .Q(\current_src_addr[1][22] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][23]$_DFF_PN0_  (.D(_0175_),
    .Q(\current_src_addr[1][23] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][24]$_DFF_PN0_  (.D(_0176_),
    .Q(\current_src_addr[1][24] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][25]$_DFF_PN0_  (.D(_0177_),
    .Q(\current_src_addr[1][25] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][26]$_DFF_PN0_  (.D(_0178_),
    .Q(\current_src_addr[1][26] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][27]$_DFF_PN0_  (.D(_0179_),
    .Q(\current_src_addr[1][27] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][28]$_DFF_PN0_  (.D(_0180_),
    .Q(\current_src_addr[1][28] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][29]$_DFF_PN0_  (.D(_0181_),
    .Q(\current_src_addr[1][29] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][2]$_DFF_PN0_  (.D(_0182_),
    .Q(\current_src_addr[1][2] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][30]$_DFF_PN0_  (.D(_0183_),
    .Q(\current_src_addr[1][30] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][31]$_DFF_PN0_  (.D(_0184_),
    .Q(\current_src_addr[1][31] ),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][3]$_DFF_PN0_  (.D(_0185_),
    .Q(\current_src_addr[1][3] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][4]$_DFF_PN0_  (.D(_0186_),
    .Q(\current_src_addr[1][4] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][5]$_DFF_PN0_  (.D(_0187_),
    .Q(\current_src_addr[1][5] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][6]$_DFF_PN0_  (.D(_0188_),
    .Q(\current_src_addr[1][6] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][7]$_DFF_PN0_  (.D(_0189_),
    .Q(\current_src_addr[1][7] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][8]$_DFF_PN0_  (.D(_0190_),
    .Q(\current_src_addr[1][8] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[1][9]$_DFF_PN0_  (.D(_0191_),
    .Q(\current_src_addr[1][9] ),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][0]$_DFFE_PN0P_  (.D(_0922_),
    .Q(\current_src_addr[2][0] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][10]$_DFF_PN0_  (.D(_0192_),
    .Q(\current_src_addr[2][10] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][11]$_DFF_PN0_  (.D(_0193_),
    .Q(\current_src_addr[2][11] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][12]$_DFF_PN0_  (.D(_0194_),
    .Q(\current_src_addr[2][12] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][13]$_DFF_PN0_  (.D(_0195_),
    .Q(\current_src_addr[2][13] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][14]$_DFF_PN0_  (.D(_0196_),
    .Q(\current_src_addr[2][14] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][15]$_DFF_PN0_  (.D(_0197_),
    .Q(\current_src_addr[2][15] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][16]$_DFF_PN0_  (.D(_0198_),
    .Q(\current_src_addr[2][16] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][17]$_DFF_PN0_  (.D(_0199_),
    .Q(\current_src_addr[2][17] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][18]$_DFF_PN0_  (.D(_0200_),
    .Q(\current_src_addr[2][18] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][19]$_DFF_PN0_  (.D(_0201_),
    .Q(\current_src_addr[2][19] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][1]$_DFFE_PN0P_  (.D(_0923_),
    .Q(\current_src_addr[2][1] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][20]$_DFF_PN0_  (.D(_0202_),
    .Q(\current_src_addr[2][20] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][21]$_DFF_PN0_  (.D(_0203_),
    .Q(\current_src_addr[2][21] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][22]$_DFF_PN0_  (.D(_0204_),
    .Q(\current_src_addr[2][22] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][23]$_DFF_PN0_  (.D(_0205_),
    .Q(\current_src_addr[2][23] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][24]$_DFF_PN0_  (.D(_0206_),
    .Q(\current_src_addr[2][24] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][25]$_DFF_PN0_  (.D(_0207_),
    .Q(\current_src_addr[2][25] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][26]$_DFF_PN0_  (.D(_0208_),
    .Q(\current_src_addr[2][26] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][27]$_DFF_PN0_  (.D(_0209_),
    .Q(\current_src_addr[2][27] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][28]$_DFF_PN0_  (.D(_0210_),
    .Q(\current_src_addr[2][28] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][29]$_DFF_PN0_  (.D(_0211_),
    .Q(\current_src_addr[2][29] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][2]$_DFF_PN0_  (.D(_0212_),
    .Q(\current_src_addr[2][2] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][30]$_DFF_PN0_  (.D(_0213_),
    .Q(\current_src_addr[2][30] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][31]$_DFF_PN0_  (.D(_0214_),
    .Q(\current_src_addr[2][31] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][3]$_DFF_PN0_  (.D(_0215_),
    .Q(\current_src_addr[2][3] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][4]$_DFF_PN0_  (.D(_0216_),
    .Q(\current_src_addr[2][4] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][5]$_DFF_PN0_  (.D(_0217_),
    .Q(\current_src_addr[2][5] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][6]$_DFF_PN0_  (.D(_0218_),
    .Q(\current_src_addr[2][6] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][7]$_DFF_PN0_  (.D(_0219_),
    .Q(\current_src_addr[2][7] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][8]$_DFF_PN0_  (.D(_0220_),
    .Q(\current_src_addr[2][8] ),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[2][9]$_DFF_PN0_  (.D(_0221_),
    .Q(\current_src_addr[2][9] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][0]$_DFFE_PN0P_  (.D(_0924_),
    .Q(\current_src_addr[3][0] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][10]$_DFF_PN0_  (.D(_0222_),
    .Q(\current_src_addr[3][10] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][11]$_DFF_PN0_  (.D(_0223_),
    .Q(\current_src_addr[3][11] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][12]$_DFF_PN0_  (.D(_0224_),
    .Q(\current_src_addr[3][12] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][13]$_DFF_PN0_  (.D(_0225_),
    .Q(\current_src_addr[3][13] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][14]$_DFF_PN0_  (.D(_0226_),
    .Q(\current_src_addr[3][14] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][15]$_DFF_PN0_  (.D(_0227_),
    .Q(\current_src_addr[3][15] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][16]$_DFF_PN0_  (.D(_0228_),
    .Q(\current_src_addr[3][16] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][17]$_DFF_PN0_  (.D(_0229_),
    .Q(\current_src_addr[3][17] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][18]$_DFF_PN0_  (.D(_0230_),
    .Q(\current_src_addr[3][18] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][19]$_DFF_PN0_  (.D(_0231_),
    .Q(\current_src_addr[3][19] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][1]$_DFFE_PN0P_  (.D(_0925_),
    .Q(\current_src_addr[3][1] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][20]$_DFF_PN0_  (.D(_0232_),
    .Q(\current_src_addr[3][20] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][21]$_DFF_PN0_  (.D(_0233_),
    .Q(\current_src_addr[3][21] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][22]$_DFF_PN0_  (.D(_0234_),
    .Q(\current_src_addr[3][22] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][23]$_DFF_PN0_  (.D(_0235_),
    .Q(\current_src_addr[3][23] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][24]$_DFF_PN0_  (.D(_0236_),
    .Q(\current_src_addr[3][24] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][25]$_DFF_PN0_  (.D(_0237_),
    .Q(\current_src_addr[3][25] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][26]$_DFF_PN0_  (.D(_0238_),
    .Q(\current_src_addr[3][26] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][27]$_DFF_PN0_  (.D(_0239_),
    .Q(\current_src_addr[3][27] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][28]$_DFF_PN0_  (.D(_0240_),
    .Q(\current_src_addr[3][28] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][29]$_DFF_PN0_  (.D(_0241_),
    .Q(\current_src_addr[3][29] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][2]$_DFF_PN0_  (.D(_0242_),
    .Q(\current_src_addr[3][2] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][30]$_DFF_PN0_  (.D(_0243_),
    .Q(\current_src_addr[3][30] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][31]$_DFF_PN0_  (.D(_0244_),
    .Q(\current_src_addr[3][31] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][3]$_DFF_PN0_  (.D(_0245_),
    .Q(\current_src_addr[3][3] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][4]$_DFF_PN0_  (.D(_0246_),
    .Q(\current_src_addr[3][4] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][5]$_DFF_PN0_  (.D(_0247_),
    .Q(\current_src_addr[3][5] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][6]$_DFF_PN0_  (.D(_0248_),
    .Q(\current_src_addr[3][6] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][7]$_DFF_PN0_  (.D(_0249_),
    .Q(\current_src_addr[3][7] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][8]$_DFF_PN0_  (.D(_0250_),
    .Q(\current_src_addr[3][8] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \current_src_addr[3][9]$_DFF_PN0_  (.D(_0251_),
    .Q(\current_src_addr[3][9] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][0]$_DFFE_PN0P_  (.D(_0926_),
    .Q(\data_buffer[0][0] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][10]$_DFFE_PN0P_  (.D(_0927_),
    .Q(\data_buffer[0][10] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][11]$_DFFE_PN0P_  (.D(_0928_),
    .Q(\data_buffer[0][11] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][12]$_DFFE_PN0P_  (.D(_0929_),
    .Q(\data_buffer[0][12] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][13]$_DFFE_PN0P_  (.D(_0930_),
    .Q(\data_buffer[0][13] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][14]$_DFFE_PN0P_  (.D(_0931_),
    .Q(\data_buffer[0][14] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][15]$_DFFE_PN0P_  (.D(_0932_),
    .Q(\data_buffer[0][15] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][16]$_DFFE_PN0P_  (.D(_0933_),
    .Q(\data_buffer[0][16] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][17]$_DFFE_PN0P_  (.D(_0934_),
    .Q(\data_buffer[0][17] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][18]$_DFFE_PN0P_  (.D(_0935_),
    .Q(\data_buffer[0][18] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][19]$_DFFE_PN0P_  (.D(_0936_),
    .Q(\data_buffer[0][19] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][1]$_DFFE_PN0P_  (.D(_0937_),
    .Q(\data_buffer[0][1] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][20]$_DFFE_PN0P_  (.D(_0938_),
    .Q(\data_buffer[0][20] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][21]$_DFFE_PN0P_  (.D(_0939_),
    .Q(\data_buffer[0][21] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][22]$_DFFE_PN0P_  (.D(_0940_),
    .Q(\data_buffer[0][22] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][23]$_DFFE_PN0P_  (.D(_0941_),
    .Q(\data_buffer[0][23] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][24]$_DFFE_PN0P_  (.D(_0942_),
    .Q(\data_buffer[0][24] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][25]$_DFFE_PN0P_  (.D(_0943_),
    .Q(\data_buffer[0][25] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][26]$_DFFE_PN0P_  (.D(_0944_),
    .Q(\data_buffer[0][26] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][27]$_DFFE_PN0P_  (.D(_0945_),
    .Q(\data_buffer[0][27] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][28]$_DFFE_PN0P_  (.D(_0946_),
    .Q(\data_buffer[0][28] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][29]$_DFFE_PN0P_  (.D(_0947_),
    .Q(\data_buffer[0][29] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][2]$_DFFE_PN0P_  (.D(_0948_),
    .Q(\data_buffer[0][2] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][30]$_DFFE_PN0P_  (.D(_0949_),
    .Q(\data_buffer[0][30] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][31]$_DFFE_PN0P_  (.D(_0950_),
    .Q(\data_buffer[0][31] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][3]$_DFFE_PN0P_  (.D(_0951_),
    .Q(\data_buffer[0][3] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][4]$_DFFE_PN0P_  (.D(_0952_),
    .Q(\data_buffer[0][4] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][5]$_DFFE_PN0P_  (.D(_0953_),
    .Q(\data_buffer[0][5] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][6]$_DFFE_PN0P_  (.D(_0954_),
    .Q(\data_buffer[0][6] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][7]$_DFFE_PN0P_  (.D(_0955_),
    .Q(\data_buffer[0][7] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][8]$_DFFE_PN0P_  (.D(_0956_),
    .Q(\data_buffer[0][8] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[0][9]$_DFFE_PN0P_  (.D(_0957_),
    .Q(\data_buffer[0][9] ),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][0]$_DFFE_PN0P_  (.D(_0958_),
    .Q(\data_buffer[1][0] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][10]$_DFFE_PN0P_  (.D(_0959_),
    .Q(\data_buffer[1][10] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][11]$_DFFE_PN0P_  (.D(_0960_),
    .Q(\data_buffer[1][11] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][12]$_DFFE_PN0P_  (.D(_0961_),
    .Q(\data_buffer[1][12] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][13]$_DFFE_PN0P_  (.D(_0962_),
    .Q(\data_buffer[1][13] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][14]$_DFFE_PN0P_  (.D(_0963_),
    .Q(\data_buffer[1][14] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][15]$_DFFE_PN0P_  (.D(_0964_),
    .Q(\data_buffer[1][15] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][16]$_DFFE_PN0P_  (.D(_0965_),
    .Q(\data_buffer[1][16] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][17]$_DFFE_PN0P_  (.D(_0966_),
    .Q(\data_buffer[1][17] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][18]$_DFFE_PN0P_  (.D(_0967_),
    .Q(\data_buffer[1][18] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][19]$_DFFE_PN0P_  (.D(_0968_),
    .Q(\data_buffer[1][19] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][1]$_DFFE_PN0P_  (.D(_0969_),
    .Q(\data_buffer[1][1] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][20]$_DFFE_PN0P_  (.D(_0970_),
    .Q(\data_buffer[1][20] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][21]$_DFFE_PN0P_  (.D(_0971_),
    .Q(\data_buffer[1][21] ),
    .RESET_B(net1286),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][22]$_DFFE_PN0P_  (.D(_0972_),
    .Q(\data_buffer[1][22] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][23]$_DFFE_PN0P_  (.D(_0973_),
    .Q(\data_buffer[1][23] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][24]$_DFFE_PN0P_  (.D(_0974_),
    .Q(\data_buffer[1][24] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][25]$_DFFE_PN0P_  (.D(_0975_),
    .Q(\data_buffer[1][25] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][26]$_DFFE_PN0P_  (.D(_0976_),
    .Q(\data_buffer[1][26] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][27]$_DFFE_PN0P_  (.D(_0977_),
    .Q(\data_buffer[1][27] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][28]$_DFFE_PN0P_  (.D(_0978_),
    .Q(\data_buffer[1][28] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][29]$_DFFE_PN0P_  (.D(_0979_),
    .Q(\data_buffer[1][29] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][2]$_DFFE_PN0P_  (.D(_0980_),
    .Q(\data_buffer[1][2] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][30]$_DFFE_PN0P_  (.D(_0981_),
    .Q(\data_buffer[1][30] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][31]$_DFFE_PN0P_  (.D(_0982_),
    .Q(\data_buffer[1][31] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][3]$_DFFE_PN0P_  (.D(_0983_),
    .Q(\data_buffer[1][3] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][4]$_DFFE_PN0P_  (.D(_0984_),
    .Q(\data_buffer[1][4] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][5]$_DFFE_PN0P_  (.D(_0985_),
    .Q(\data_buffer[1][5] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][6]$_DFFE_PN0P_  (.D(_0986_),
    .Q(\data_buffer[1][6] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][7]$_DFFE_PN0P_  (.D(_0987_),
    .Q(\data_buffer[1][7] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][8]$_DFFE_PN0P_  (.D(_0988_),
    .Q(\data_buffer[1][8] ),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[1][9]$_DFFE_PN0P_  (.D(_0989_),
    .Q(\data_buffer[1][9] ),
    .RESET_B(net1288),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][0]$_DFFE_PN0P_  (.D(_0990_),
    .Q(\data_buffer[2][0] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][10]$_DFFE_PN0P_  (.D(_0991_),
    .Q(\data_buffer[2][10] ),
    .RESET_B(net1276),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][11]$_DFFE_PN0P_  (.D(_0992_),
    .Q(\data_buffer[2][11] ),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][12]$_DFFE_PN0P_  (.D(_0993_),
    .Q(\data_buffer[2][12] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][13]$_DFFE_PN0P_  (.D(_0994_),
    .Q(\data_buffer[2][13] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][14]$_DFFE_PN0P_  (.D(_0995_),
    .Q(\data_buffer[2][14] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][15]$_DFFE_PN0P_  (.D(_0996_),
    .Q(\data_buffer[2][15] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][16]$_DFFE_PN0P_  (.D(_0997_),
    .Q(\data_buffer[2][16] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][17]$_DFFE_PN0P_  (.D(_0998_),
    .Q(\data_buffer[2][17] ),
    .RESET_B(net1276),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][18]$_DFFE_PN0P_  (.D(_0999_),
    .Q(\data_buffer[2][18] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][19]$_DFFE_PN0P_  (.D(_1000_),
    .Q(\data_buffer[2][19] ),
    .RESET_B(net1276),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][1]$_DFFE_PN0P_  (.D(_1001_),
    .Q(\data_buffer[2][1] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][20]$_DFFE_PN0P_  (.D(_1002_),
    .Q(\data_buffer[2][20] ),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][21]$_DFFE_PN0P_  (.D(_1003_),
    .Q(\data_buffer[2][21] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][22]$_DFFE_PN0P_  (.D(_1004_),
    .Q(\data_buffer[2][22] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][23]$_DFFE_PN0P_  (.D(_1005_),
    .Q(\data_buffer[2][23] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][24]$_DFFE_PN0P_  (.D(_1006_),
    .Q(\data_buffer[2][24] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][25]$_DFFE_PN0P_  (.D(_1007_),
    .Q(\data_buffer[2][25] ),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][26]$_DFFE_PN0P_  (.D(_1008_),
    .Q(\data_buffer[2][26] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][27]$_DFFE_PN0P_  (.D(_1009_),
    .Q(\data_buffer[2][27] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][28]$_DFFE_PN0P_  (.D(_1010_),
    .Q(\data_buffer[2][28] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][29]$_DFFE_PN0P_  (.D(_1011_),
    .Q(\data_buffer[2][29] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][2]$_DFFE_PN0P_  (.D(_1012_),
    .Q(\data_buffer[2][2] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][30]$_DFFE_PN0P_  (.D(_1013_),
    .Q(\data_buffer[2][30] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][31]$_DFFE_PN0P_  (.D(_1014_),
    .Q(\data_buffer[2][31] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][3]$_DFFE_PN0P_  (.D(_1015_),
    .Q(\data_buffer[2][3] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][4]$_DFFE_PN0P_  (.D(_1016_),
    .Q(\data_buffer[2][4] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][5]$_DFFE_PN0P_  (.D(_1017_),
    .Q(\data_buffer[2][5] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][6]$_DFFE_PN0P_  (.D(_1018_),
    .Q(\data_buffer[2][6] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][7]$_DFFE_PN0P_  (.D(_1019_),
    .Q(\data_buffer[2][7] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][8]$_DFFE_PN0P_  (.D(_1020_),
    .Q(\data_buffer[2][8] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[2][9]$_DFFE_PN0P_  (.D(_1021_),
    .Q(\data_buffer[2][9] ),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][0]$_DFFE_PN0P_  (.D(_1022_),
    .Q(\data_buffer[3][0] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][10]$_DFFE_PN0P_  (.D(_1023_),
    .Q(\data_buffer[3][10] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][11]$_DFFE_PN0P_  (.D(_1024_),
    .Q(\data_buffer[3][11] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][12]$_DFFE_PN0P_  (.D(_1025_),
    .Q(\data_buffer[3][12] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][13]$_DFFE_PN0P_  (.D(_1026_),
    .Q(\data_buffer[3][13] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][14]$_DFFE_PN0P_  (.D(_1027_),
    .Q(\data_buffer[3][14] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][15]$_DFFE_PN0P_  (.D(_1028_),
    .Q(\data_buffer[3][15] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][16]$_DFFE_PN0P_  (.D(_1029_),
    .Q(\data_buffer[3][16] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][17]$_DFFE_PN0P_  (.D(_1030_),
    .Q(\data_buffer[3][17] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][18]$_DFFE_PN0P_  (.D(_1031_),
    .Q(\data_buffer[3][18] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][19]$_DFFE_PN0P_  (.D(_1032_),
    .Q(\data_buffer[3][19] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][1]$_DFFE_PN0P_  (.D(_1033_),
    .Q(\data_buffer[3][1] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][20]$_DFFE_PN0P_  (.D(_1034_),
    .Q(\data_buffer[3][20] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][21]$_DFFE_PN0P_  (.D(_1035_),
    .Q(\data_buffer[3][21] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][22]$_DFFE_PN0P_  (.D(_1036_),
    .Q(\data_buffer[3][22] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][23]$_DFFE_PN0P_  (.D(_1037_),
    .Q(\data_buffer[3][23] ),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][24]$_DFFE_PN0P_  (.D(_1038_),
    .Q(\data_buffer[3][24] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][25]$_DFFE_PN0P_  (.D(_1039_),
    .Q(\data_buffer[3][25] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][26]$_DFFE_PN0P_  (.D(_1040_),
    .Q(\data_buffer[3][26] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][27]$_DFFE_PN0P_  (.D(_1041_),
    .Q(\data_buffer[3][27] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][28]$_DFFE_PN0P_  (.D(_1042_),
    .Q(\data_buffer[3][28] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][29]$_DFFE_PN0P_  (.D(_1043_),
    .Q(\data_buffer[3][29] ),
    .RESET_B(net1281),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][2]$_DFFE_PN0P_  (.D(_1044_),
    .Q(\data_buffer[3][2] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][30]$_DFFE_PN0P_  (.D(_1045_),
    .Q(\data_buffer[3][30] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][31]$_DFFE_PN0P_  (.D(_1046_),
    .Q(\data_buffer[3][31] ),
    .RESET_B(net1282),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][3]$_DFFE_PN0P_  (.D(_1047_),
    .Q(\data_buffer[3][3] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][4]$_DFFE_PN0P_  (.D(_1048_),
    .Q(\data_buffer[3][4] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][5]$_DFFE_PN0P_  (.D(_1049_),
    .Q(\data_buffer[3][5] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][6]$_DFFE_PN0P_  (.D(_1050_),
    .Q(\data_buffer[3][6] ),
    .RESET_B(net1283),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][7]$_DFFE_PN0P_  (.D(_1051_),
    .Q(\data_buffer[3][7] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][8]$_DFFE_PN0P_  (.D(_1052_),
    .Q(\data_buffer[3][8] ),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_buffer[3][9]$_DFFE_PN0P_  (.D(_1053_),
    .Q(\data_buffer[3][9] ),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[0]$_DFF_PN0_  (.D(\active_channel_count[0] ),
    .Q(net550),
    .RESET_B(net1287),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[1]$_DFF_PN0_  (.D(\active_channel_count[1] ),
    .Q(net551),
    .RESET_B(net1287),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[2]$_DFF_PN0_  (.D(\active_channel_count[2] ),
    .Q(net552),
    .RESET_B(net1287),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_active_channels[3]$_DFF_PN0_  (.D(\active_channel_count[3] ),
    .Q(net553),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \debug_has_active_channels$_DFF_PN0_  (.D(_0252_),
    .Q(net566),
    .RESET_B(net1287),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[0]$_DFFE_PN0P_  (.D(_1054_),
    .Q(net695),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[100]$_DFFE_PN0P_  (.D(_1055_),
    .Q(net696),
    .RESET_B(net1295),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[101]$_DFFE_PN0P_  (.D(_1056_),
    .Q(net697),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[102]$_DFFE_PN0P_  (.D(_1057_),
    .Q(net698),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[103]$_DFFE_PN0P_  (.D(_1058_),
    .Q(net699),
    .RESET_B(net1284),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[104]$_DFFE_PN0P_  (.D(_1059_),
    .Q(net700),
    .RESET_B(net1283),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[105]$_DFFE_PN0P_  (.D(_1060_),
    .Q(net701),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[106]$_DFFE_PN0P_  (.D(_1061_),
    .Q(net702),
    .RESET_B(net1283),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[107]$_DFFE_PN0P_  (.D(_1062_),
    .Q(net703),
    .RESET_B(net1283),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[108]$_DFFE_PN0P_  (.D(_1063_),
    .Q(net704),
    .RESET_B(net1295),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[109]$_DFFE_PN0P_  (.D(_1064_),
    .Q(net705),
    .RESET_B(net1285),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[10]$_DFFE_PN0P_  (.D(_1065_),
    .Q(net706),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[110]$_DFFE_PN0P_  (.D(_1066_),
    .Q(net707),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[111]$_DFFE_PN0P_  (.D(_1067_),
    .Q(net708),
    .RESET_B(net1284),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[112]$_DFFE_PN0P_  (.D(_1068_),
    .Q(net709),
    .RESET_B(net1295),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[113]$_DFFE_PN0P_  (.D(_1069_),
    .Q(net710),
    .RESET_B(net1295),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[114]$_DFFE_PN0P_  (.D(_1070_),
    .Q(net711),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[115]$_DFFE_PN0P_  (.D(_1071_),
    .Q(net712),
    .RESET_B(net1284),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[116]$_DFFE_PN0P_  (.D(_1072_),
    .Q(net713),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[117]$_DFFE_PN0P_  (.D(_1073_),
    .Q(net714),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[118]$_DFFE_PN0P_  (.D(_1074_),
    .Q(net715),
    .RESET_B(net1295),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[119]$_DFFE_PN0P_  (.D(_1075_),
    .Q(net716),
    .RESET_B(net1285),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[11]$_DFFE_PN0P_  (.D(_1076_),
    .Q(net717),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[120]$_DFFE_PN0P_  (.D(_1077_),
    .Q(net718),
    .RESET_B(net1295),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[121]$_DFFE_PN0P_  (.D(_1078_),
    .Q(net719),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[122]$_DFFE_PN0P_  (.D(_1079_),
    .Q(net720),
    .RESET_B(net1285),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[123]$_DFFE_PN0P_  (.D(_1080_),
    .Q(net721),
    .RESET_B(net1295),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[124]$_DFFE_PN0P_  (.D(_1081_),
    .Q(net722),
    .RESET_B(net1283),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[125]$_DFFE_PN0P_  (.D(_1082_),
    .Q(net723),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[126]$_DFFE_PN0P_  (.D(_1083_),
    .Q(net724),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[127]$_DFFE_PN0P_  (.D(_1084_),
    .Q(net725),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[12]$_DFFE_PN0P_  (.D(_1085_),
    .Q(net726),
    .RESET_B(net1278),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[13]$_DFFE_PN0P_  (.D(_1086_),
    .Q(net727),
    .RESET_B(net1278),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[14]$_DFFE_PN0P_  (.D(_1087_),
    .Q(net728),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[15]$_DFFE_PN0P_  (.D(_1088_),
    .Q(net729),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[16]$_DFFE_PN0P_  (.D(_1089_),
    .Q(net730),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[17]$_DFFE_PN0P_  (.D(_1090_),
    .Q(net731),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[18]$_DFFE_PN0P_  (.D(_1091_),
    .Q(net732),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[19]$_DFFE_PN0P_  (.D(_1092_),
    .Q(net733),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[1]$_DFFE_PN0P_  (.D(_1093_),
    .Q(net734),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[20]$_DFFE_PN0P_  (.D(_1094_),
    .Q(net735),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[21]$_DFFE_PN0P_  (.D(_1095_),
    .Q(net736),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[22]$_DFFE_PN0P_  (.D(_1096_),
    .Q(net737),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[23]$_DFFE_PN0P_  (.D(_1097_),
    .Q(net738),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[24]$_DFFE_PN0P_  (.D(_1098_),
    .Q(net739),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[25]$_DFFE_PN0P_  (.D(_1099_),
    .Q(net740),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[26]$_DFFE_PN0P_  (.D(_1100_),
    .Q(net741),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[27]$_DFFE_PN0P_  (.D(_1101_),
    .Q(net742),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[28]$_DFFE_PN0P_  (.D(_1102_),
    .Q(net743),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[29]$_DFFE_PN0P_  (.D(_1103_),
    .Q(net744),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[2]$_DFFE_PN0P_  (.D(_1104_),
    .Q(net745),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[30]$_DFFE_PN0P_  (.D(_1105_),
    .Q(net746),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[31]$_DFFE_PN0P_  (.D(_1106_),
    .Q(net747),
    .RESET_B(net1278),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[32]$_DFFE_PN0P_  (.D(_1107_),
    .Q(net748),
    .RESET_B(net1287),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[33]$_DFFE_PN0P_  (.D(_1108_),
    .Q(net749),
    .RESET_B(net1287),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[34]$_DFFE_PN0P_  (.D(_1109_),
    .Q(net750),
    .RESET_B(net1292),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[35]$_DFFE_PN0P_  (.D(_1110_),
    .Q(net751),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[36]$_DFFE_PN0P_  (.D(_1111_),
    .Q(net752),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[37]$_DFFE_PN0P_  (.D(_1112_),
    .Q(net753),
    .RESET_B(net1291),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[38]$_DFFE_PN0P_  (.D(_1113_),
    .Q(net754),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[39]$_DFFE_PN0P_  (.D(_1114_),
    .Q(net755),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[3]$_DFFE_PN0P_  (.D(_1115_),
    .Q(net756),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[40]$_DFFE_PN0P_  (.D(_1116_),
    .Q(net757),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[41]$_DFFE_PN0P_  (.D(_1117_),
    .Q(net758),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[42]$_DFFE_PN0P_  (.D(_1118_),
    .Q(net759),
    .RESET_B(net1290),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[43]$_DFFE_PN0P_  (.D(_1119_),
    .Q(net760),
    .RESET_B(net1290),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[44]$_DFFE_PN0P_  (.D(_1120_),
    .Q(net761),
    .RESET_B(net1290),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[45]$_DFFE_PN0P_  (.D(_1121_),
    .Q(net762),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[46]$_DFFE_PN0P_  (.D(_1122_),
    .Q(net763),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[47]$_DFFE_PN0P_  (.D(_1123_),
    .Q(net764),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[48]$_DFFE_PN0P_  (.D(_1124_),
    .Q(net765),
    .RESET_B(net1291),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[49]$_DFFE_PN0P_  (.D(_1125_),
    .Q(net766),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[4]$_DFFE_PN0P_  (.D(_1126_),
    .Q(net767),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[50]$_DFFE_PN0P_  (.D(_1127_),
    .Q(net768),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[51]$_DFFE_PN0P_  (.D(_1128_),
    .Q(net769),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[52]$_DFFE_PN0P_  (.D(_1129_),
    .Q(net770),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[53]$_DFFE_PN0P_  (.D(_1130_),
    .Q(net771),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[54]$_DFFE_PN0P_  (.D(_1131_),
    .Q(net772),
    .RESET_B(net1292),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[55]$_DFFE_PN0P_  (.D(_1132_),
    .Q(net773),
    .RESET_B(net1292),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[56]$_DFFE_PN0P_  (.D(_1133_),
    .Q(net774),
    .RESET_B(net1292),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[57]$_DFFE_PN0P_  (.D(_1134_),
    .Q(net775),
    .RESET_B(net1292),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[58]$_DFFE_PN0P_  (.D(_1135_),
    .Q(net776),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[59]$_DFFE_PN0P_  (.D(_1136_),
    .Q(net777),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[5]$_DFFE_PN0P_  (.D(_1137_),
    .Q(net778),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[60]$_DFFE_PN0P_  (.D(_1138_),
    .Q(net779),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[61]$_DFFE_PN0P_  (.D(_1139_),
    .Q(net780),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[62]$_DFFE_PN0P_  (.D(_1140_),
    .Q(net781),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[63]$_DFFE_PN0P_  (.D(_1141_),
    .Q(net782),
    .RESET_B(net1292),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[64]$_DFFE_PN0P_  (.D(_1142_),
    .Q(net783),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[65]$_DFFE_PN0P_  (.D(_1143_),
    .Q(net784),
    .RESET_B(net1281),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[66]$_DFFE_PN0P_  (.D(_1144_),
    .Q(net785),
    .RESET_B(net1275),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[67]$_DFFE_PN0P_  (.D(_1145_),
    .Q(net786),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[68]$_DFFE_PN0P_  (.D(_1146_),
    .Q(net787),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[69]$_DFFE_PN0P_  (.D(_1147_),
    .Q(net788),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[6]$_DFFE_PN0P_  (.D(_1148_),
    .Q(net789),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[70]$_DFFE_PN0P_  (.D(_1149_),
    .Q(net790),
    .RESET_B(net1274),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[71]$_DFFE_PN0P_  (.D(_1150_),
    .Q(net791),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[72]$_DFFE_PN0P_  (.D(_1151_),
    .Q(net792),
    .RESET_B(net1275),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[73]$_DFFE_PN0P_  (.D(_1152_),
    .Q(net793),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[74]$_DFFE_PN0P_  (.D(_1153_),
    .Q(net794),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[75]$_DFFE_PN0P_  (.D(_1154_),
    .Q(net795),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[76]$_DFFE_PN0P_  (.D(_1155_),
    .Q(net796),
    .RESET_B(net1275),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[77]$_DFFE_PN0P_  (.D(_1156_),
    .Q(net797),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[78]$_DFFE_PN0P_  (.D(_1157_),
    .Q(net798),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[79]$_DFFE_PN0P_  (.D(_1158_),
    .Q(net799),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[7]$_DFFE_PN0P_  (.D(_1159_),
    .Q(net800),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[80]$_DFFE_PN0P_  (.D(_1160_),
    .Q(net801),
    .RESET_B(net1274),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[81]$_DFFE_PN0P_  (.D(_1161_),
    .Q(net802),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[82]$_DFFE_PN0P_  (.D(_1162_),
    .Q(net803),
    .RESET_B(net1274),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[83]$_DFFE_PN0P_  (.D(_1163_),
    .Q(net804),
    .RESET_B(net1281),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[84]$_DFFE_PN0P_  (.D(_1164_),
    .Q(net805),
    .RESET_B(net1280),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[85]$_DFFE_PN0P_  (.D(_1165_),
    .Q(net806),
    .RESET_B(net1274),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[86]$_DFFE_PN0P_  (.D(_1166_),
    .Q(net807),
    .RESET_B(net1280),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[87]$_DFFE_PN0P_  (.D(_1167_),
    .Q(net808),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[88]$_DFFE_PN0P_  (.D(_1168_),
    .Q(net809),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[89]$_DFFE_PN0P_  (.D(_1169_),
    .Q(net810),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[8]$_DFFE_PN0P_  (.D(_1170_),
    .Q(net811),
    .RESET_B(net1278),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[90]$_DFFE_PN0P_  (.D(_1171_),
    .Q(net812),
    .RESET_B(net1274),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[91]$_DFFE_PN0P_  (.D(_1172_),
    .Q(net813),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[92]$_DFFE_PN0P_  (.D(_1173_),
    .Q(net814),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[93]$_DFFE_PN0P_  (.D(_1174_),
    .Q(net815),
    .RESET_B(net1274),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[94]$_DFFE_PN0P_  (.D(_1175_),
    .Q(net816),
    .RESET_B(net1274),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[95]$_DFFE_PN0P_  (.D(_1176_),
    .Q(net817),
    .RESET_B(net1275),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[96]$_DFFE_PN0P_  (.D(_1177_),
    .Q(net818),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[97]$_DFFE_PN0P_  (.D(_1178_),
    .Q(net819),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[98]$_DFFE_PN0P_  (.D(_1179_),
    .Q(net820),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[99]$_DFFE_PN0P_  (.D(_1180_),
    .Q(net821),
    .RESET_B(net1295),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_addr[9]$_DFFE_PN0P_  (.D(_1181_),
    .Q(net822),
    .RESET_B(net1278),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[0]$_DFFE_PN0P_  (.D(_1182_),
    .Q(net823),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[100]$_DFFE_PN0P_  (.D(_1183_),
    .Q(net824),
    .RESET_B(net1283),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[101]$_DFFE_PN0P_  (.D(_1184_),
    .Q(net825),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[102]$_DFFE_PN0P_  (.D(_1185_),
    .Q(net826),
    .RESET_B(net1283),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[103]$_DFFE_PN0P_  (.D(_1186_),
    .Q(net827),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[104]$_DFFE_PN0P_  (.D(_1187_),
    .Q(net828),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[105]$_DFFE_PN0P_  (.D(_1188_),
    .Q(net829),
    .RESET_B(net1284),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[106]$_DFFE_PN0P_  (.D(_1189_),
    .Q(net830),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[107]$_DFFE_PN0P_  (.D(_1190_),
    .Q(net831),
    .RESET_B(net1281),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[108]$_DFFE_PN0P_  (.D(_1191_),
    .Q(net832),
    .RESET_B(net1281),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[109]$_DFFE_PN0P_  (.D(_1192_),
    .Q(net833),
    .RESET_B(net1282),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[10]$_DFFE_PN0P_  (.D(_1193_),
    .Q(net834),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[110]$_DFFE_PN0P_  (.D(_1194_),
    .Q(net835),
    .RESET_B(net1282),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[111]$_DFFE_PN0P_  (.D(_1195_),
    .Q(net836),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[112]$_DFFE_PN0P_  (.D(_1196_),
    .Q(net837),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[113]$_DFFE_PN0P_  (.D(_1197_),
    .Q(net838),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[114]$_DFFE_PN0P_  (.D(_1198_),
    .Q(net839),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[115]$_DFFE_PN0P_  (.D(_1199_),
    .Q(net840),
    .RESET_B(net1281),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[116]$_DFFE_PN0P_  (.D(_1200_),
    .Q(net841),
    .RESET_B(net1282),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[117]$_DFFE_PN0P_  (.D(_1201_),
    .Q(net842),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[118]$_DFFE_PN0P_  (.D(_1202_),
    .Q(net843),
    .RESET_B(net1281),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[119]$_DFFE_PN0P_  (.D(_1203_),
    .Q(net844),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[11]$_DFFE_PN0P_  (.D(_1204_),
    .Q(net845),
    .RESET_B(net1278),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[120]$_DFFE_PN0P_  (.D(_1205_),
    .Q(net846),
    .RESET_B(net1281),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[121]$_DFFE_PN0P_  (.D(_1206_),
    .Q(net847),
    .RESET_B(net1281),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[122]$_DFFE_PN0P_  (.D(_1207_),
    .Q(net848),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[123]$_DFFE_PN0P_  (.D(_1208_),
    .Q(net849),
    .RESET_B(net1282),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[124]$_DFFE_PN0P_  (.D(_1209_),
    .Q(net850),
    .RESET_B(net1282),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[125]$_DFFE_PN0P_  (.D(_1210_),
    .Q(net851),
    .RESET_B(net1281),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[126]$_DFFE_PN0P_  (.D(_1211_),
    .Q(net852),
    .RESET_B(net1282),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[127]$_DFFE_PN0P_  (.D(_1212_),
    .Q(net853),
    .RESET_B(net1282),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[12]$_DFFE_PN0P_  (.D(_1213_),
    .Q(net854),
    .RESET_B(net1278),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[13]$_DFFE_PN0P_  (.D(_1214_),
    .Q(net855),
    .RESET_B(net1278),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[14]$_DFFE_PN0P_  (.D(_1215_),
    .Q(net856),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[15]$_DFFE_PN0P_  (.D(_1216_),
    .Q(net857),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[16]$_DFFE_PN0P_  (.D(_1217_),
    .Q(net858),
    .RESET_B(net1278),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[17]$_DFFE_PN0P_  (.D(_1218_),
    .Q(net859),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[18]$_DFFE_PN0P_  (.D(_1219_),
    .Q(net860),
    .RESET_B(net1277),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[19]$_DFFE_PN0P_  (.D(_1220_),
    .Q(net861),
    .RESET_B(net1277),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[1]$_DFFE_PN0P_  (.D(_1221_),
    .Q(net862),
    .RESET_B(net1277),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[20]$_DFFE_PN0P_  (.D(_1222_),
    .Q(net863),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[21]$_DFFE_PN0P_  (.D(_1223_),
    .Q(net864),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[22]$_DFFE_PN0P_  (.D(_1224_),
    .Q(net865),
    .RESET_B(net1277),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[23]$_DFFE_PN0P_  (.D(_1225_),
    .Q(net866),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[24]$_DFFE_PN0P_  (.D(_1226_),
    .Q(net867),
    .RESET_B(net1278),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[25]$_DFFE_PN0P_  (.D(_1227_),
    .Q(net868),
    .RESET_B(net1278),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[26]$_DFFE_PN0P_  (.D(_1228_),
    .Q(net869),
    .RESET_B(net1277),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[27]$_DFFE_PN0P_  (.D(_1229_),
    .Q(net870),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[28]$_DFFE_PN0P_  (.D(_1230_),
    .Q(net871),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[29]$_DFFE_PN0P_  (.D(_1231_),
    .Q(net872),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[2]$_DFFE_PN0P_  (.D(_1232_),
    .Q(net873),
    .RESET_B(net1278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[30]$_DFFE_PN0P_  (.D(_1233_),
    .Q(net874),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[31]$_DFFE_PN0P_  (.D(_1234_),
    .Q(net875),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[32]$_DFFE_PN0P_  (.D(_1235_),
    .Q(net876),
    .RESET_B(net1288),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[33]$_DFFE_PN0P_  (.D(_1236_),
    .Q(net877),
    .RESET_B(net1284),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[34]$_DFFE_PN0P_  (.D(_1237_),
    .Q(net878),
    .RESET_B(net1287),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[35]$_DFFE_PN0P_  (.D(_1238_),
    .Q(net879),
    .RESET_B(net1287),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[36]$_DFFE_PN0P_  (.D(_1239_),
    .Q(net880),
    .RESET_B(net1284),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[37]$_DFFE_PN0P_  (.D(_1240_),
    .Q(net881),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[38]$_DFFE_PN0P_  (.D(_1241_),
    .Q(net882),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[39]$_DFFE_PN0P_  (.D(_1242_),
    .Q(net883),
    .RESET_B(net1288),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[3]$_DFFE_PN0P_  (.D(_1243_),
    .Q(net884),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[40]$_DFFE_PN0P_  (.D(_1244_),
    .Q(net885),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[41]$_DFFE_PN0P_  (.D(_1245_),
    .Q(net886),
    .RESET_B(net1288),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[42]$_DFFE_PN0P_  (.D(_1246_),
    .Q(net887),
    .RESET_B(net1288),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[43]$_DFFE_PN0P_  (.D(_1247_),
    .Q(net888),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[44]$_DFFE_PN0P_  (.D(_1248_),
    .Q(net889),
    .RESET_B(net1284),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[45]$_DFFE_PN0P_  (.D(_1249_),
    .Q(net890),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[46]$_DFFE_PN0P_  (.D(_1250_),
    .Q(net891),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[47]$_DFFE_PN0P_  (.D(_1251_),
    .Q(net892),
    .RESET_B(net1284),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[48]$_DFFE_PN0P_  (.D(_1252_),
    .Q(net893),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[49]$_DFFE_PN0P_  (.D(_1253_),
    .Q(net894),
    .RESET_B(net1284),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[4]$_DFFE_PN0P_  (.D(_1254_),
    .Q(net895),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[50]$_DFFE_PN0P_  (.D(_1255_),
    .Q(net896),
    .RESET_B(net1284),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[51]$_DFFE_PN0P_  (.D(_1256_),
    .Q(net897),
    .RESET_B(net1284),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[52]$_DFFE_PN0P_  (.D(_1257_),
    .Q(net898),
    .RESET_B(net1288),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[53]$_DFFE_PN0P_  (.D(_1258_),
    .Q(net899),
    .RESET_B(net1286),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[54]$_DFFE_PN0P_  (.D(_1259_),
    .Q(net900),
    .RESET_B(net1284),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[55]$_DFFE_PN0P_  (.D(_1260_),
    .Q(net901),
    .RESET_B(net1287),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[56]$_DFFE_PN0P_  (.D(_1261_),
    .Q(net902),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[57]$_DFFE_PN0P_  (.D(_1262_),
    .Q(net903),
    .RESET_B(net1284),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[58]$_DFFE_PN0P_  (.D(_1263_),
    .Q(net904),
    .RESET_B(net1288),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[59]$_DFFE_PN0P_  (.D(_1264_),
    .Q(net905),
    .RESET_B(net1288),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[5]$_DFFE_PN0P_  (.D(_1265_),
    .Q(net906),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[60]$_DFFE_PN0P_  (.D(_1266_),
    .Q(net907),
    .RESET_B(net1288),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[61]$_DFFE_PN0P_  (.D(_1267_),
    .Q(net908),
    .RESET_B(net1288),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[62]$_DFFE_PN0P_  (.D(_1268_),
    .Q(net909),
    .RESET_B(net1288),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[63]$_DFFE_PN0P_  (.D(_1269_),
    .Q(net910),
    .RESET_B(net1288),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[64]$_DFFE_PN0P_  (.D(_1270_),
    .Q(net911),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[65]$_DFFE_PN0P_  (.D(_1271_),
    .Q(net912),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[66]$_DFFE_PN0P_  (.D(_1272_),
    .Q(net913),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[67]$_DFFE_PN0P_  (.D(_1273_),
    .Q(net914),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[68]$_DFFE_PN0P_  (.D(_1274_),
    .Q(net915),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[69]$_DFFE_PN0P_  (.D(_1275_),
    .Q(net916),
    .RESET_B(net1277),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[6]$_DFFE_PN0P_  (.D(_1276_),
    .Q(net917),
    .RESET_B(net1278),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[70]$_DFFE_PN0P_  (.D(_1277_),
    .Q(net918),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[71]$_DFFE_PN0P_  (.D(_1278_),
    .Q(net919),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[72]$_DFFE_PN0P_  (.D(_1279_),
    .Q(net920),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[73]$_DFFE_PN0P_  (.D(_1280_),
    .Q(net921),
    .RESET_B(net1295),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[74]$_DFFE_PN0P_  (.D(_1281_),
    .Q(net922),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[75]$_DFFE_PN0P_  (.D(_1282_),
    .Q(net923),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[76]$_DFFE_PN0P_  (.D(_1283_),
    .Q(net924),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[77]$_DFFE_PN0P_  (.D(_1284_),
    .Q(net925),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[78]$_DFFE_PN0P_  (.D(_1285_),
    .Q(net926),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[79]$_DFFE_PN0P_  (.D(_1286_),
    .Q(net927),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[7]$_DFFE_PN0P_  (.D(_1287_),
    .Q(net928),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[80]$_DFFE_PN0P_  (.D(_1288_),
    .Q(net929),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[81]$_DFFE_PN0P_  (.D(_1289_),
    .Q(net930),
    .RESET_B(net1276),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[82]$_DFFE_PN0P_  (.D(_1290_),
    .Q(net931),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[83]$_DFFE_PN0P_  (.D(_1291_),
    .Q(net932),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[84]$_DFFE_PN0P_  (.D(_1292_),
    .Q(net933),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[85]$_DFFE_PN0P_  (.D(_1293_),
    .Q(net934),
    .RESET_B(net1295),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[86]$_DFFE_PN0P_  (.D(_1294_),
    .Q(net935),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[87]$_DFFE_PN0P_  (.D(_1295_),
    .Q(net936),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[88]$_DFFE_PN0P_  (.D(_1296_),
    .Q(net937),
    .RESET_B(net1277),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[89]$_DFFE_PN0P_  (.D(_1297_),
    .Q(net938),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[8]$_DFFE_PN0P_  (.D(_1298_),
    .Q(net939),
    .RESET_B(net1278),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[90]$_DFFE_PN0P_  (.D(_1299_),
    .Q(net940),
    .RESET_B(net1277),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[91]$_DFFE_PN0P_  (.D(_1300_),
    .Q(net941),
    .RESET_B(net1277),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[92]$_DFFE_PN0P_  (.D(_1301_),
    .Q(net942),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[93]$_DFFE_PN0P_  (.D(_1302_),
    .Q(net943),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[94]$_DFFE_PN0P_  (.D(_1303_),
    .Q(net944),
    .RESET_B(net1277),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[95]$_DFFE_PN0P_  (.D(_1304_),
    .Q(net945),
    .RESET_B(net1277),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[96]$_DFFE_PN0P_  (.D(_1305_),
    .Q(net946),
    .RESET_B(net1283),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[97]$_DFFE_PN0P_  (.D(_1306_),
    .Q(net947),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[98]$_DFFE_PN0P_  (.D(_1307_),
    .Q(net948),
    .RESET_B(net1283),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[99]$_DFFE_PN0P_  (.D(_1308_),
    .Q(net949),
    .RESET_B(net1283),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wdata[9]$_DFFE_PN0P_  (.D(_1309_),
    .Q(net950),
    .RESET_B(net1278),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[0]$_DFFE_PN0P_  (.D(_1310_),
    .Q(net951),
    .RESET_B(net1278),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[1]$_DFFE_PN0P_  (.D(_1311_),
    .Q(net952),
    .RESET_B(net1292),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[2]$_DFFE_PN0P_  (.D(_1312_),
    .Q(net953),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_write[3]$_DFFE_PN0P_  (.D(_1313_),
    .Q(net954),
    .RESET_B(net1283),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wstrb[10]$_DFFE_PN0P_  (.D(_1314_),
    .Q(net957),
    .RESET_B(net1295),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wstrb[14]$_DFFE_PN0P_  (.D(_1315_),
    .Q(net961),
    .RESET_B(net1295),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wstrb[2]$_DFFE_PN0P_  (.D(_1316_),
    .Q(net964),
    .RESET_B(net1278),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfrtp_1 \dst_wstrb[6]$_DFFE_PN0P_  (.D(_1317_),
    .Q(net968),
    .RESET_B(net1288),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[0]$_DFFE_PN0P_  (.D(_1318_),
    .Q(net971),
    .RESET_B(net1278),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[100]$_DFFE_PN0P_  (.D(_1319_),
    .Q(net972),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[101]$_DFFE_PN0P_  (.D(_1320_),
    .Q(net973),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[102]$_DFFE_PN0P_  (.D(_1321_),
    .Q(net974),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[103]$_DFFE_PN0P_  (.D(_1322_),
    .Q(net975),
    .RESET_B(net1287),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[104]$_DFFE_PN0P_  (.D(_1323_),
    .Q(net976),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[105]$_DFFE_PN0P_  (.D(_1324_),
    .Q(net977),
    .RESET_B(net1286),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[106]$_DFFE_PN0P_  (.D(_1325_),
    .Q(net978),
    .RESET_B(net1286),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[107]$_DFFE_PN0P_  (.D(_1326_),
    .Q(net979),
    .RESET_B(net1284),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[108]$_DFFE_PN0P_  (.D(_1327_),
    .Q(net980),
    .RESET_B(net1284),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[109]$_DFFE_PN0P_  (.D(_1328_),
    .Q(net981),
    .RESET_B(net1284),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[10]$_DFFE_PN0P_  (.D(_1329_),
    .Q(net982),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[110]$_DFFE_PN0P_  (.D(_1330_),
    .Q(net983),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[111]$_DFFE_PN0P_  (.D(_1331_),
    .Q(net984),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[112]$_DFFE_PN0P_  (.D(_1332_),
    .Q(net985),
    .RESET_B(net1284),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[113]$_DFFE_PN0P_  (.D(_1333_),
    .Q(net986),
    .RESET_B(net1287),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[114]$_DFFE_PN0P_  (.D(_1334_),
    .Q(net987),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[115]$_DFFE_PN0P_  (.D(_1335_),
    .Q(net988),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[116]$_DFFE_PN0P_  (.D(_1336_),
    .Q(net989),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[117]$_DFFE_PN0P_  (.D(_1337_),
    .Q(net990),
    .RESET_B(net1286),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[118]$_DFFE_PN0P_  (.D(_1338_),
    .Q(net991),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[119]$_DFFE_PN0P_  (.D(_1339_),
    .Q(net992),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[11]$_DFFE_PN0P_  (.D(_1340_),
    .Q(net993),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[120]$_DFFE_PN0P_  (.D(_1341_),
    .Q(net994),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[121]$_DFFE_PN0P_  (.D(_1342_),
    .Q(net995),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[122]$_DFFE_PN0P_  (.D(_1343_),
    .Q(net996),
    .RESET_B(net1285),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[123]$_DFFE_PN0P_  (.D(_1344_),
    .Q(net997),
    .RESET_B(net1285),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[124]$_DFFE_PN0P_  (.D(_1345_),
    .Q(net998),
    .RESET_B(net1284),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[125]$_DFFE_PN0P_  (.D(_1346_),
    .Q(net999),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[126]$_DFFE_PN0P_  (.D(_1347_),
    .Q(net1000),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[127]$_DFFE_PN0P_  (.D(_1348_),
    .Q(net1001),
    .RESET_B(net1286),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[12]$_DFFE_PN0P_  (.D(_1349_),
    .Q(net1002),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[13]$_DFFE_PN0P_  (.D(_1350_),
    .Q(net1003),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[14]$_DFFE_PN0P_  (.D(_1351_),
    .Q(net1004),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[15]$_DFFE_PN0P_  (.D(_1352_),
    .Q(net1005),
    .RESET_B(net1279),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[16]$_DFFE_PN0P_  (.D(_1353_),
    .Q(net1006),
    .RESET_B(net1279),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[17]$_DFFE_PN0P_  (.D(_1354_),
    .Q(net1007),
    .RESET_B(net1279),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[18]$_DFFE_PN0P_  (.D(_1355_),
    .Q(net1008),
    .RESET_B(net1279),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[19]$_DFFE_PN0P_  (.D(_1356_),
    .Q(net1009),
    .RESET_B(net1278),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[1]$_DFFE_PN0P_  (.D(_1357_),
    .Q(net1010),
    .RESET_B(net1278),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[20]$_DFFE_PN0P_  (.D(_1358_),
    .Q(net1011),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[21]$_DFFE_PN0P_  (.D(_1359_),
    .Q(net1012),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[22]$_DFFE_PN0P_  (.D(_1360_),
    .Q(net1013),
    .RESET_B(net1279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[23]$_DFFE_PN0P_  (.D(_1361_),
    .Q(net1014),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[24]$_DFFE_PN0P_  (.D(_1362_),
    .Q(net1015),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[25]$_DFFE_PN0P_  (.D(_1363_),
    .Q(net1016),
    .RESET_B(net1291),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[26]$_DFFE_PN0P_  (.D(_1364_),
    .Q(net1017),
    .RESET_B(net1291),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[27]$_DFFE_PN0P_  (.D(_1365_),
    .Q(net1018),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[28]$_DFFE_PN0P_  (.D(_1366_),
    .Q(net1019),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[29]$_DFFE_PN0P_  (.D(_1367_),
    .Q(net1020),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[2]$_DFFE_PN0P_  (.D(_1368_),
    .Q(net1021),
    .RESET_B(net1279),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[30]$_DFFE_PN0P_  (.D(_1369_),
    .Q(net1022),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[31]$_DFFE_PN0P_  (.D(_1370_),
    .Q(net1023),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[32]$_DFFE_PN0P_  (.D(_1371_),
    .Q(net1024),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[33]$_DFFE_PN0P_  (.D(_1372_),
    .Q(net1025),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[34]$_DFFE_PN0P_  (.D(_1373_),
    .Q(net1026),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[35]$_DFFE_PN0P_  (.D(_1374_),
    .Q(net1027),
    .RESET_B(net1291),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[36]$_DFFE_PN0P_  (.D(_1375_),
    .Q(net1028),
    .RESET_B(net1291),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[37]$_DFFE_PN0P_  (.D(_1376_),
    .Q(net1029),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[38]$_DFFE_PN0P_  (.D(_1377_),
    .Q(net1030),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[39]$_DFFE_PN0P_  (.D(_1378_),
    .Q(net1031),
    .RESET_B(net1291),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[3]$_DFFE_PN0P_  (.D(_1379_),
    .Q(net1032),
    .RESET_B(net1279),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[40]$_DFFE_PN0P_  (.D(_1380_),
    .Q(net1033),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[41]$_DFFE_PN0P_  (.D(_1381_),
    .Q(net1034),
    .RESET_B(net1291),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[42]$_DFFE_PN0P_  (.D(_1382_),
    .Q(net1035),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[43]$_DFFE_PN0P_  (.D(_1383_),
    .Q(net1036),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[44]$_DFFE_PN0P_  (.D(_1384_),
    .Q(net1037),
    .RESET_B(net1292),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[45]$_DFFE_PN0P_  (.D(_1385_),
    .Q(net1038),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[46]$_DFFE_PN0P_  (.D(_1386_),
    .Q(net1039),
    .RESET_B(net1291),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[47]$_DFFE_PN0P_  (.D(_1387_),
    .Q(net1040),
    .RESET_B(net1291),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[48]$_DFFE_PN0P_  (.D(_1388_),
    .Q(net1041),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[49]$_DFFE_PN0P_  (.D(_1389_),
    .Q(net1042),
    .RESET_B(net1291),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[4]$_DFFE_PN0P_  (.D(_1390_),
    .Q(net1043),
    .RESET_B(net1279),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[50]$_DFFE_PN0P_  (.D(_1391_),
    .Q(net1044),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[51]$_DFFE_PN0P_  (.D(_1392_),
    .Q(net1045),
    .RESET_B(net1292),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[52]$_DFFE_PN0P_  (.D(_1393_),
    .Q(net1046),
    .RESET_B(net1292),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[53]$_DFFE_PN0P_  (.D(_1394_),
    .Q(net1047),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[54]$_DFFE_PN0P_  (.D(_1395_),
    .Q(net1048),
    .RESET_B(net1292),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[55]$_DFFE_PN0P_  (.D(_1396_),
    .Q(net1049),
    .RESET_B(net1291),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[56]$_DFFE_PN0P_  (.D(_1397_),
    .Q(net1050),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[57]$_DFFE_PN0P_  (.D(_1398_),
    .Q(net1051),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[58]$_DFFE_PN0P_  (.D(_1399_),
    .Q(net1052),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[59]$_DFFE_PN0P_  (.D(_1400_),
    .Q(net1053),
    .RESET_B(net1292),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[5]$_DFFE_PN0P_  (.D(_1401_),
    .Q(net1054),
    .RESET_B(net1279),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[60]$_DFFE_PN0P_  (.D(_1402_),
    .Q(net1055),
    .RESET_B(net1291),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[61]$_DFFE_PN0P_  (.D(_1403_),
    .Q(net1056),
    .RESET_B(net1291),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[62]$_DFFE_PN0P_  (.D(_1404_),
    .Q(net1057),
    .RESET_B(net1292),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[63]$_DFFE_PN0P_  (.D(_1405_),
    .Q(net1058),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[64]$_DFFE_PN0P_  (.D(_1406_),
    .Q(net1059),
    .RESET_B(net1281),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[65]$_DFFE_PN0P_  (.D(_1407_),
    .Q(net1060),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[66]$_DFFE_PN0P_  (.D(_1408_),
    .Q(net1061),
    .RESET_B(net1280),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[67]$_DFFE_PN0P_  (.D(_1409_),
    .Q(net1062),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[68]$_DFFE_PN0P_  (.D(_1410_),
    .Q(net1063),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[69]$_DFFE_PN0P_  (.D(_1411_),
    .Q(net1064),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[6]$_DFFE_PN0P_  (.D(_1412_),
    .Q(net1065),
    .RESET_B(net1279),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[70]$_DFFE_PN0P_  (.D(_1413_),
    .Q(net1066),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[71]$_DFFE_PN0P_  (.D(_1414_),
    .Q(net1067),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[72]$_DFFE_PN0P_  (.D(_1415_),
    .Q(net1068),
    .RESET_B(net1274),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[73]$_DFFE_PN0P_  (.D(_1416_),
    .Q(net1069),
    .RESET_B(net1282),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[74]$_DFFE_PN0P_  (.D(_1417_),
    .Q(net1070),
    .RESET_B(net1280),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[75]$_DFFE_PN0P_  (.D(_1418_),
    .Q(net1071),
    .RESET_B(net1281),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[76]$_DFFE_PN0P_  (.D(_1419_),
    .Q(net1072),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[77]$_DFFE_PN0P_  (.D(_1420_),
    .Q(net1073),
    .RESET_B(net1281),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[78]$_DFFE_PN0P_  (.D(_1421_),
    .Q(net1074),
    .RESET_B(net1280),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[79]$_DFFE_PN0P_  (.D(_1422_),
    .Q(net1075),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[7]$_DFFE_PN0P_  (.D(_1423_),
    .Q(net1076),
    .RESET_B(net1279),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[80]$_DFFE_PN0P_  (.D(_1424_),
    .Q(net1077),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[81]$_DFFE_PN0P_  (.D(_1425_),
    .Q(net1078),
    .RESET_B(net1280),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[82]$_DFFE_PN0P_  (.D(_1426_),
    .Q(net1079),
    .RESET_B(net1281),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[83]$_DFFE_PN0P_  (.D(_1427_),
    .Q(net1080),
    .RESET_B(net1281),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[84]$_DFFE_PN0P_  (.D(_1428_),
    .Q(net1081),
    .RESET_B(net1282),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[85]$_DFFE_PN0P_  (.D(_1429_),
    .Q(net1082),
    .RESET_B(net1282),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[86]$_DFFE_PN0P_  (.D(_1430_),
    .Q(net1083),
    .RESET_B(net1282),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[87]$_DFFE_PN0P_  (.D(_1431_),
    .Q(net1084),
    .RESET_B(net1281),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[88]$_DFFE_PN0P_  (.D(_1432_),
    .Q(net1085),
    .RESET_B(net1281),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[89]$_DFFE_PN0P_  (.D(_1433_),
    .Q(net1086),
    .RESET_B(net1282),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[8]$_DFFE_PN0P_  (.D(_1434_),
    .Q(net1087),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[90]$_DFFE_PN0P_  (.D(_1435_),
    .Q(net1088),
    .RESET_B(net1282),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[91]$_DFFE_PN0P_  (.D(_1436_),
    .Q(net1089),
    .RESET_B(net1281),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[92]$_DFFE_PN0P_  (.D(_1437_),
    .Q(net1090),
    .RESET_B(net1281),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[93]$_DFFE_PN0P_  (.D(_1438_),
    .Q(net1091),
    .RESET_B(net1281),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[94]$_DFFE_PN0P_  (.D(_1439_),
    .Q(net1092),
    .RESET_B(net1281),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[95]$_DFFE_PN0P_  (.D(_1440_),
    .Q(net1093),
    .RESET_B(net1282),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[96]$_DFFE_PN0P_  (.D(_1441_),
    .Q(net1094),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[97]$_DFFE_PN0P_  (.D(_1442_),
    .Q(net1095),
    .RESET_B(net1285),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[98]$_DFFE_PN0P_  (.D(_1443_),
    .Q(net1096),
    .RESET_B(net1284),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[99]$_DFFE_PN0P_  (.D(_1444_),
    .Q(net1097),
    .RESET_B(net1284),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_addr[9]$_DFFE_PN0P_  (.D(_1445_),
    .Q(net1098),
    .RESET_B(net1279),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_read[0]$_DFF_PN0_  (.D(net1252),
    .Q(net1099),
    .RESET_B(net1292),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_read[1]$_DFF_PN0_  (.D(net1269),
    .Q(net1100),
    .RESET_B(net1292),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_read[2]$_DFF_PN0_  (.D(net1254),
    .Q(net1101),
    .RESET_B(net1276),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_read[3]$_DFF_PN0_  (.D(net1253),
    .Q(net1102),
    .RESET_B(net1286),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_rready[0]$_DFFE_PN0P_  (.D(_1446_),
    .Q(net1103),
    .RESET_B(net1278),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_rready[1]$_DFFE_PN0P_  (.D(_1447_),
    .Q(net1104),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_rready[2]$_DFFE_PN0P_  (.D(_1448_),
    .Q(net1105),
    .RESET_B(net1276),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_rready[3]$_DFFE_PN0P_  (.D(_1449_),
    .Q(net1106),
    .RESET_B(net1283),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][0]$_DFF_PN0_  (.D(_0253_),
    .Q(net567),
    .RESET_B(net1279),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][10]$_DFF_PN0_  (.D(_0254_),
    .Q(net578),
    .RESET_B(net1279),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][11]$_DFF_PN0_  (.D(_0255_),
    .Q(net589),
    .RESET_B(net1277),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][12]$_DFF_PN0_  (.D(_0256_),
    .Q(net598),
    .RESET_B(net1277),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][13]$_DFF_PN0_  (.D(_0257_),
    .Q(net599),
    .RESET_B(net1277),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][14]$_DFF_PN0_  (.D(_0258_),
    .Q(net600),
    .RESET_B(net1277),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][15]$_DFF_PN0_  (.D(_0259_),
    .Q(net601),
    .RESET_B(net1277),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][16]$_DFF_PN0_  (.D(_0260_),
    .Q(net602),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][17]$_DFF_PN0_  (.D(_0261_),
    .Q(net603),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][18]$_DFF_PN0_  (.D(_0262_),
    .Q(net604),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][19]$_DFF_PN0_  (.D(_0263_),
    .Q(net605),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][1]$_DFF_PN0_  (.D(_0264_),
    .Q(net606),
    .RESET_B(net1279),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][20]$_DFF_PN0_  (.D(_0265_),
    .Q(net607),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][21]$_DFF_PN0_  (.D(_0266_),
    .Q(net608),
    .RESET_B(net1277),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][22]$_DFF_PN0_  (.D(_0267_),
    .Q(net609),
    .RESET_B(net1277),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][23]$_DFF_PN0_  (.D(_0268_),
    .Q(net610),
    .RESET_B(net1277),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][24]$_DFF_PN0_  (.D(_0269_),
    .Q(net611),
    .RESET_B(net1277),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][25]$_DFF_PN0_  (.D(_0270_),
    .Q(net612),
    .RESET_B(net1279),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][26]$_DFF_PN0_  (.D(_0271_),
    .Q(net613),
    .RESET_B(net1279),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][27]$_DFF_PN0_  (.D(_0272_),
    .Q(net614),
    .RESET_B(net1278),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][28]$_DFF_PN0_  (.D(_0273_),
    .Q(net615),
    .RESET_B(net1278),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][29]$_DFF_PN0_  (.D(_0274_),
    .Q(net616),
    .RESET_B(net1278),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][2]$_DFF_PN0_  (.D(_0275_),
    .Q(net617),
    .RESET_B(net1279),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][30]$_DFF_PN0_  (.D(_0276_),
    .Q(net618),
    .RESET_B(net1279),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][31]$_DFF_PN0_  (.D(_0277_),
    .Q(net619),
    .RESET_B(net1278),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][3]$_DFF_PN0_  (.D(_0278_),
    .Q(net628),
    .RESET_B(net1277),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][4]$_DFF_PN0_  (.D(_0279_),
    .Q(net639),
    .RESET_B(net1277),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][5]$_DFF_PN0_  (.D(_0280_),
    .Q(net650),
    .RESET_B(net1277),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][6]$_DFF_PN0_  (.D(_0281_),
    .Q(net661),
    .RESET_B(net1277),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][7]$_DFF_PN0_  (.D(_0282_),
    .Q(net672),
    .RESET_B(net1277),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][8]$_DFF_PN0_  (.D(_0283_),
    .Q(net683),
    .RESET_B(net1279),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[0][9]$_DFF_PN0_  (.D(_0284_),
    .Q(net694),
    .RESET_B(net1279),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][0]$_DFF_PN0_  (.D(_0285_),
    .Q(net620),
    .RESET_B(net1289),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][10]$_DFF_PN0_  (.D(_0286_),
    .Q(net631),
    .RESET_B(net1289),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][11]$_DFF_PN0_  (.D(_0287_),
    .Q(net632),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][12]$_DFF_PN0_  (.D(_0288_),
    .Q(net633),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][13]$_DFF_PN0_  (.D(_0289_),
    .Q(net634),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][14]$_DFF_PN0_  (.D(_0290_),
    .Q(net635),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][15]$_DFF_PN0_  (.D(_0291_),
    .Q(net636),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][16]$_DFF_PN0_  (.D(_0292_),
    .Q(net637),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][17]$_DFF_PN0_  (.D(_0293_),
    .Q(net638),
    .RESET_B(net1289),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][18]$_DFF_PN0_  (.D(_0294_),
    .Q(net640),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][19]$_DFF_PN0_  (.D(_0295_),
    .Q(net641),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][1]$_DFF_PN0_  (.D(_0296_),
    .Q(net621),
    .RESET_B(net1289),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][20]$_DFF_PN0_  (.D(_0297_),
    .Q(net642),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][21]$_DFF_PN0_  (.D(_0298_),
    .Q(net643),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][22]$_DFF_PN0_  (.D(_0299_),
    .Q(net644),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][23]$_DFF_PN0_  (.D(_0300_),
    .Q(net645),
    .RESET_B(net1290),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][24]$_DFF_PN0_  (.D(_0301_),
    .Q(net646),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][25]$_DFF_PN0_  (.D(_0302_),
    .Q(net647),
    .RESET_B(net1289),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][26]$_DFF_PN0_  (.D(_0303_),
    .Q(net648),
    .RESET_B(net1290),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][27]$_DFF_PN0_  (.D(_0304_),
    .Q(net649),
    .RESET_B(net1289),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][28]$_DFF_PN0_  (.D(_0305_),
    .Q(net651),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][29]$_DFF_PN0_  (.D(_0306_),
    .Q(net652),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][2]$_DFF_PN0_  (.D(_0307_),
    .Q(net622),
    .RESET_B(net1289),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][30]$_DFF_PN0_  (.D(_0308_),
    .Q(net653),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][31]$_DFF_PN0_  (.D(_0309_),
    .Q(net654),
    .RESET_B(net1290),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][3]$_DFF_PN0_  (.D(_0310_),
    .Q(net623),
    .RESET_B(net1289),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][4]$_DFF_PN0_  (.D(_0311_),
    .Q(net624),
    .RESET_B(net1284),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][5]$_DFF_PN0_  (.D(_0312_),
    .Q(net625),
    .RESET_B(net1284),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][6]$_DFF_PN0_  (.D(_0313_),
    .Q(net626),
    .RESET_B(net1290),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][7]$_DFF_PN0_  (.D(_0314_),
    .Q(net627),
    .RESET_B(net1290),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][8]$_DFF_PN0_  (.D(_0315_),
    .Q(net629),
    .RESET_B(net1290),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[1][9]$_DFF_PN0_  (.D(_0316_),
    .Q(net630),
    .RESET_B(net1290),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][0]$_DFF_PN0_  (.D(_0317_),
    .Q(net655),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][10]$_DFF_PN0_  (.D(_0318_),
    .Q(net666),
    .RESET_B(net1276),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][11]$_DFF_PN0_  (.D(_0319_),
    .Q(net667),
    .RESET_B(net1276),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][12]$_DFF_PN0_  (.D(_0320_),
    .Q(net668),
    .RESET_B(net1276),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][13]$_DFF_PN0_  (.D(_0321_),
    .Q(net669),
    .RESET_B(net1276),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][14]$_DFF_PN0_  (.D(_0322_),
    .Q(net670),
    .RESET_B(net1276),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][15]$_DFF_PN0_  (.D(_0323_),
    .Q(net671),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][16]$_DFF_PN0_  (.D(_0324_),
    .Q(net673),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][17]$_DFF_PN0_  (.D(_0325_),
    .Q(net674),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][18]$_DFF_PN0_  (.D(_0326_),
    .Q(net675),
    .RESET_B(net1276),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][19]$_DFF_PN0_  (.D(_0327_),
    .Q(net676),
    .RESET_B(net1276),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][1]$_DFF_PN0_  (.D(_0328_),
    .Q(net656),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][20]$_DFF_PN0_  (.D(_0329_),
    .Q(net677),
    .RESET_B(net1276),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][21]$_DFF_PN0_  (.D(_0330_),
    .Q(net678),
    .RESET_B(net1295),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][22]$_DFF_PN0_  (.D(_0331_),
    .Q(net679),
    .RESET_B(net1295),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][23]$_DFF_PN0_  (.D(_0332_),
    .Q(net680),
    .RESET_B(net1277),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][24]$_DFF_PN0_  (.D(_0333_),
    .Q(net681),
    .RESET_B(net1295),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][25]$_DFF_PN0_  (.D(_0334_),
    .Q(net682),
    .RESET_B(net1277),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][26]$_DFF_PN0_  (.D(_0335_),
    .Q(net684),
    .RESET_B(net1277),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][27]$_DFF_PN0_  (.D(_0336_),
    .Q(net685),
    .RESET_B(net1295),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][28]$_DFF_PN0_  (.D(_0337_),
    .Q(net686),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][29]$_DFF_PN0_  (.D(_0338_),
    .Q(net687),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][2]$_DFF_PN0_  (.D(_0339_),
    .Q(net657),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][30]$_DFF_PN0_  (.D(_0340_),
    .Q(net688),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][31]$_DFF_PN0_  (.D(_0341_),
    .Q(net689),
    .RESET_B(net1277),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][3]$_DFF_PN0_  (.D(_0342_),
    .Q(net658),
    .RESET_B(net1274),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][4]$_DFF_PN0_  (.D(_0343_),
    .Q(net659),
    .RESET_B(net1274),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][5]$_DFF_PN0_  (.D(_0344_),
    .Q(net660),
    .RESET_B(net1274),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][6]$_DFF_PN0_  (.D(_0345_),
    .Q(net662),
    .RESET_B(net1274),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][7]$_DFF_PN0_  (.D(_0346_),
    .Q(net663),
    .RESET_B(net1276),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][8]$_DFF_PN0_  (.D(_0347_),
    .Q(net664),
    .RESET_B(net1276),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[2][9]$_DFF_PN0_  (.D(_0348_),
    .Q(net665),
    .RESET_B(net1276),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][0]$_DFF_PN0_  (.D(_0349_),
    .Q(net690),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][10]$_DFF_PN0_  (.D(_0350_),
    .Q(net574),
    .RESET_B(net1283),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][11]$_DFF_PN0_  (.D(_0351_),
    .Q(net575),
    .RESET_B(net1283),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][12]$_DFF_PN0_  (.D(_0352_),
    .Q(net576),
    .RESET_B(net1283),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][13]$_DFF_PN0_  (.D(_0353_),
    .Q(net577),
    .RESET_B(net1283),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][14]$_DFF_PN0_  (.D(_0354_),
    .Q(net579),
    .RESET_B(net1283),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][15]$_DFF_PN0_  (.D(_0355_),
    .Q(net580),
    .RESET_B(net1283),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][16]$_DFF_PN0_  (.D(_0356_),
    .Q(net581),
    .RESET_B(net1283),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][17]$_DFF_PN0_  (.D(_0357_),
    .Q(net582),
    .RESET_B(net1283),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][18]$_DFF_PN0_  (.D(_0358_),
    .Q(net583),
    .RESET_B(net1283),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][19]$_DFF_PN0_  (.D(_0359_),
    .Q(net584),
    .RESET_B(net1283),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][1]$_DFF_PN0_  (.D(_0360_),
    .Q(net691),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][20]$_DFF_PN0_  (.D(_0361_),
    .Q(net585),
    .RESET_B(net1283),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][21]$_DFF_PN0_  (.D(_0362_),
    .Q(net586),
    .RESET_B(net1283),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][22]$_DFF_PN0_  (.D(_0363_),
    .Q(net587),
    .RESET_B(net1287),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][23]$_DFF_PN0_  (.D(_0364_),
    .Q(net588),
    .RESET_B(net1283),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][24]$_DFF_PN0_  (.D(_0365_),
    .Q(net590),
    .RESET_B(net1283),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][25]$_DFF_PN0_  (.D(_0366_),
    .Q(net591),
    .RESET_B(net1283),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][26]$_DFF_PN0_  (.D(_0367_),
    .Q(net592),
    .RESET_B(net1287),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][27]$_DFF_PN0_  (.D(_0368_),
    .Q(net593),
    .RESET_B(net1287),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][28]$_DFF_PN0_  (.D(_0369_),
    .Q(net594),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][29]$_DFF_PN0_  (.D(_0370_),
    .Q(net595),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][2]$_DFF_PN0_  (.D(_0371_),
    .Q(net692),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][30]$_DFF_PN0_  (.D(_0372_),
    .Q(net596),
    .RESET_B(net1283),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][31]$_DFF_PN0_  (.D(_0373_),
    .Q(net597),
    .RESET_B(net1287),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][3]$_DFF_PN0_  (.D(_0374_),
    .Q(net693),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][4]$_DFF_PN0_  (.D(_0375_),
    .Q(net568),
    .RESET_B(net1283),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][5]$_DFF_PN0_  (.D(_0376_),
    .Q(net569),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][6]$_DFF_PN0_  (.D(_0377_),
    .Q(net570),
    .RESET_B(net1283),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][7]$_DFF_PN0_  (.D(_0378_),
    .Q(net571),
    .RESET_B(net1283),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][8]$_DFF_PN0_  (.D(_0379_),
    .Q(net572),
    .RESET_B(net1283),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \transfer_count[3][9]$_DFF_PN0_  (.D(_0380_),
    .Q(net573),
    .RESET_B(net1283),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input222 (.A(channel_length[65]),
    .X(net222));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input223 (.A(channel_length[66]),
    .X(net223));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input224 (.A(channel_length[67]),
    .X(net224));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input225 (.A(channel_length[68]),
    .X(net225));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input226 (.A(channel_length[69]),
    .X(net226));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input227 (.A(channel_length[6]),
    .X(net227));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input228 (.A(channel_length[70]),
    .X(net228));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input229 (.A(channel_length[71]),
    .X(net229));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input230 (.A(channel_length[72]),
    .X(net230));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input231 (.A(channel_length[73]),
    .X(net231));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input232 (.A(channel_length[74]),
    .X(net232));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input233 (.A(channel_length[75]),
    .X(net233));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input234 (.A(channel_length[76]),
    .X(net234));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input235 (.A(channel_length[77]),
    .X(net235));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input236 (.A(channel_length[78]),
    .X(net236));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input237 (.A(channel_length[79]),
    .X(net237));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input238 (.A(channel_length[7]),
    .X(net238));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input239 (.A(channel_length[80]),
    .X(net239));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input240 (.A(channel_length[81]),
    .X(net240));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input241 (.A(channel_length[82]),
    .X(net241));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input242 (.A(channel_length[83]),
    .X(net242));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input243 (.A(channel_length[84]),
    .X(net243));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input244 (.A(channel_length[85]),
    .X(net244));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input245 (.A(channel_length[86]),
    .X(net245));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input246 (.A(channel_length[87]),
    .X(net246));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input247 (.A(channel_length[88]),
    .X(net247));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input248 (.A(channel_length[89]),
    .X(net248));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input249 (.A(channel_length[8]),
    .X(net249));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input250 (.A(channel_length[90]),
    .X(net250));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input251 (.A(channel_length[91]),
    .X(net251));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input252 (.A(channel_length[92]),
    .X(net252));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input253 (.A(channel_length[93]),
    .X(net253));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input254 (.A(channel_length[94]),
    .X(net254));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input255 (.A(channel_length[95]),
    .X(net255));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input256 (.A(channel_length[96]),
    .X(net256));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input257 (.A(channel_length[97]),
    .X(net257));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input258 (.A(channel_length[98]),
    .X(net258));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input259 (.A(channel_length[99]),
    .X(net259));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input260 (.A(channel_length[9]),
    .X(net260));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input261 (.A(channel_mode[0]),
    .X(net261));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input262 (.A(channel_mode[1]),
    .X(net262));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input263 (.A(channel_mode[2]),
    .X(net263));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input264 (.A(channel_mode[3]),
    .X(net264));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input265 (.A(channel_mode[4]),
    .X(net265));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input266 (.A(channel_mode[5]),
    .X(net266));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input267 (.A(channel_mode[6]),
    .X(net267));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input268 (.A(channel_mode[7]),
    .X(net268));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input269 (.A(net1593),
    .X(net269));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input270 (.A(net1571),
    .X(net270));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input271 (.A(channel_src_addr[101]),
    .X(net271));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input272 (.A(net1640),
    .X(net272));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input273 (.A(channel_src_addr[103]),
    .X(net273));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input274 (.A(net1599),
    .X(net274));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input275 (.A(net1488),
    .X(net275));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input276 (.A(net1423),
    .X(net276));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input277 (.A(net1518),
    .X(net277));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input278 (.A(net1566),
    .X(net278));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input279 (.A(net1437),
    .X(net279));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input280 (.A(net1533),
    .X(net280));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input281 (.A(net1591),
    .X(net281));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input282 (.A(net1392),
    .X(net282));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input283 (.A(net1430),
    .X(net283));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input284 (.A(net1462),
    .X(net284));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input285 (.A(net1641),
    .X(net285));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input286 (.A(net1551),
    .X(net286));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input287 (.A(net1532),
    .X(net287));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input288 (.A(net1477),
    .X(net288));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input289 (.A(net1486),
    .X(net289));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input290 (.A(channel_src_addr[119]),
    .X(net290));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input291 (.A(net1544),
    .X(net291));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input292 (.A(net1573),
    .X(net292));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input293 (.A(net1491),
    .X(net293));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input294 (.A(net1455),
    .X(net294));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input295 (.A(net1439),
    .X(net295));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input296 (.A(net1482),
    .X(net296));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input297 (.A(channel_src_addr[125]),
    .X(net297));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input298 (.A(channel_src_addr[126]),
    .X(net298));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input299 (.A(net1596),
    .X(net299));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input300 (.A(net1567),
    .X(net300));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input301 (.A(net1639),
    .X(net301));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input302 (.A(net1543),
    .X(net302));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input303 (.A(net1558),
    .X(net303));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input304 (.A(net1592),
    .X(net304));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input305 (.A(net1589),
    .X(net305));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input306 (.A(net1624),
    .X(net306));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input307 (.A(net1612),
    .X(net307));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input308 (.A(net1387),
    .X(net308));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input309 (.A(net1565),
    .X(net309));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input310 (.A(net1608),
    .X(net310));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input311 (.A(net1575),
    .X(net311));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input312 (.A(net1426),
    .X(net312));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input313 (.A(net1457),
    .X(net313));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input314 (.A(net1509),
    .X(net314));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input315 (.A(net1429),
    .X(net315));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input316 (.A(net1370),
    .X(net316));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input317 (.A(net1480),
    .X(net317));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input318 (.A(net1445),
    .X(net318));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input319 (.A(net1603),
    .X(net319));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input320 (.A(channel_src_addr[30]),
    .X(net320));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input321 (.A(net1534),
    .X(net321));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input322 (.A(net1303),
    .X(net322));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input323 (.A(net1305),
    .X(net323));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input324 (.A(net1522),
    .X(net324));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input325 (.A(channel_src_addr[35]),
    .X(net325));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input326 (.A(channel_src_addr[36]),
    .X(net326));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input327 (.A(channel_src_addr[37]),
    .X(net327));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input328 (.A(net1613),
    .X(net328));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input329 (.A(net1610),
    .X(net329));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input330 (.A(net1561),
    .X(net330));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input331 (.A(net1576),
    .X(net331));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input332 (.A(net1475),
    .X(net332));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input333 (.A(channel_src_addr[42]),
    .X(net333));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input334 (.A(net1379),
    .X(net334));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input335 (.A(net1456),
    .X(net335));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input336 (.A(net1422),
    .X(net336));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input337 (.A(channel_src_addr[46]),
    .X(net337));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input338 (.A(net1557),
    .X(net338));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input339 (.A(net1474),
    .X(net339));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input340 (.A(net1469),
    .X(net340));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input341 (.A(channel_src_addr[4]),
    .X(net341));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input342 (.A(net1619),
    .X(net342));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input343 (.A(net1452),
    .X(net343));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input344 (.A(net1420),
    .X(net344));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input345 (.A(net1421),
    .X(net345));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input346 (.A(net1633),
    .X(net346));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input347 (.A(net1583),
    .X(net347));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input348 (.A(net1481),
    .X(net348));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input349 (.A(net1564),
    .X(net349));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input350 (.A(net1537),
    .X(net350));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input351 (.A(net1443),
    .X(net351));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input352 (.A(net1617),
    .X(net352));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input353 (.A(net1520),
    .X(net353));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input354 (.A(net1466),
    .X(net354));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input355 (.A(net1440),
    .X(net355));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input356 (.A(net1435),
    .X(net356));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input357 (.A(net1326),
    .X(net357));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input358 (.A(net1296),
    .X(net358));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input359 (.A(net1331),
    .X(net359));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input360 (.A(net1463),
    .X(net360));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input361 (.A(net1465),
    .X(net361));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input362 (.A(net1504),
    .X(net362));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input363 (.A(net1584),
    .X(net363));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input364 (.A(channel_src_addr[70]),
    .X(net364));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input365 (.A(net1632),
    .X(net365));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input366 (.A(channel_src_addr[72]),
    .X(net366));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input367 (.A(net1442),
    .X(net367));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input368 (.A(net1316),
    .X(net368));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input369 (.A(net1327),
    .X(net369));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input370 (.A(net1626),
    .X(net370));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input371 (.A(net1367),
    .X(net371));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input372 (.A(net1476),
    .X(net372));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input373 (.A(net1400),
    .X(net373));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input374 (.A(net1642),
    .X(net374));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input375 (.A(net1340),
    .X(net375));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input376 (.A(channel_src_addr[81]),
    .X(net376));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input377 (.A(net1311),
    .X(net377));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input378 (.A(net1449),
    .X(net378));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input379 (.A(channel_src_addr[84]),
    .X(net379));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input380 (.A(net1602),
    .X(net380));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input381 (.A(net1346),
    .X(net381));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input382 (.A(net1394),
    .X(net382));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input383 (.A(net1306),
    .X(net383));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input384 (.A(net1451),
    .X(net384));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input385 (.A(channel_src_addr[8]),
    .X(net385));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input386 (.A(net1343),
    .X(net386));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input387 (.A(channel_src_addr[91]),
    .X(net387));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input388 (.A(net1308),
    .X(net388));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input389 (.A(net1471),
    .X(net389));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input390 (.A(net1307),
    .X(net390));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input391 (.A(net1318),
    .X(net391));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input392 (.A(net1304),
    .X(net392));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input393 (.A(net1330),
    .X(net393));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input394 (.A(net1629),
    .X(net394));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input395 (.A(net1595),
    .X(net395));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input396 (.A(net1552),
    .X(net396));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input397 (.A(net1600),
    .X(net397));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input398 (.A(net1598),
    .X(net398));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input399 (.A(net1637),
    .X(net399));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input400 (.A(channel_start[3]),
    .X(net400));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input401 (.A(dst_wready[0]),
    .X(net401));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input402 (.A(dst_wready[1]),
    .X(net402));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input403 (.A(dst_wready[2]),
    .X(net403));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input404 (.A(dst_wready[3]),
    .X(net404));
 sky130_fd_sc_hd__buf_8 input405 (.A(net1294),
    .X(net405));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input406 (.A(net1531),
    .X(net406));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input407 (.A(src_rdata[100]),
    .X(net407));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input408 (.A(net1448),
    .X(net408));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input409 (.A(src_rdata[102]),
    .X(net409));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input410 (.A(net1460),
    .X(net410));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input411 (.A(net1517),
    .X(net411));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input412 (.A(net1441),
    .X(net412));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input413 (.A(net1495),
    .X(net413));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input414 (.A(net1317),
    .X(net414));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input415 (.A(net1347),
    .X(net415));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input416 (.A(net1335),
    .X(net416));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input417 (.A(src_rdata[10]),
    .X(net417));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input418 (.A(net1320),
    .X(net418));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input419 (.A(net1339),
    .X(net419));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input420 (.A(net1321),
    .X(net420));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input421 (.A(net1315),
    .X(net421));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input422 (.A(net1337),
    .X(net422));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input423 (.A(net1333),
    .X(net423));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input424 (.A(net1319),
    .X(net424));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input425 (.A(net1332),
    .X(net425));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input426 (.A(net1323),
    .X(net426));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input427 (.A(net1511),
    .X(net427));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input428 (.A(net1502),
    .X(net428));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input429 (.A(net1322),
    .X(net429));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input430 (.A(net1324),
    .X(net430));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input431 (.A(net1329),
    .X(net431));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input432 (.A(net1354),
    .X(net432));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input433 (.A(net1341),
    .X(net433));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input434 (.A(net1403),
    .X(net434));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input435 (.A(net1334),
    .X(net435));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input436 (.A(src_rdata[127]),
    .X(net436));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input437 (.A(net1489),
    .X(net437));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input438 (.A(net1505),
    .X(net438));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input439 (.A(net1508),
    .X(net439));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input440 (.A(net1446),
    .X(net440));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input441 (.A(net1545),
    .X(net441));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input442 (.A(net1574),
    .X(net442));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input443 (.A(net1540),
    .X(net443));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input444 (.A(net1546),
    .X(net444));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input445 (.A(net1527),
    .X(net445));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input446 (.A(net1541),
    .X(net446));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input447 (.A(net1563),
    .X(net447));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input448 (.A(net1559),
    .X(net448));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input449 (.A(net1525),
    .X(net449));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input450 (.A(net1568),
    .X(net450));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input451 (.A(net1506),
    .X(net451));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input452 (.A(net1550),
    .X(net452));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input453 (.A(net1510),
    .X(net453));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input454 (.A(net1530),
    .X(net454));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input455 (.A(net1493),
    .X(net455));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input456 (.A(net1604),
    .X(net456));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input457 (.A(net1526),
    .X(net457));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input458 (.A(net1523),
    .X(net458));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input459 (.A(net1407),
    .X(net459));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input460 (.A(net1438),
    .X(net460));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input461 (.A(net1414),
    .X(net461));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input462 (.A(net1416),
    .X(net462));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input463 (.A(net1405),
    .X(net463));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input464 (.A(net1562),
    .X(net464));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input465 (.A(net1412),
    .X(net465));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input466 (.A(net1415),
    .X(net466));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input467 (.A(net1547),
    .X(net467));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input468 (.A(net1464),
    .X(net468));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input469 (.A(net1432),
    .X(net469));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input470 (.A(net1388),
    .X(net470));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input471 (.A(net1391),
    .X(net471));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input472 (.A(net1556),
    .X(net472));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input473 (.A(net1389),
    .X(net473));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input474 (.A(src_rdata[46]),
    .X(net474));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input475 (.A(src_rdata[47]),
    .X(net475));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input476 (.A(net1425),
    .X(net476));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input477 (.A(net1512),
    .X(net477));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input478 (.A(net1529),
    .X(net478));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input479 (.A(net1513),
    .X(net479));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input480 (.A(net1535),
    .X(net480));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input481 (.A(net1395),
    .X(net481));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input482 (.A(net1514),
    .X(net482));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input483 (.A(net1555),
    .X(net483));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input484 (.A(net1424),
    .X(net484));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input485 (.A(net1408),
    .X(net485));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input486 (.A(net1413),
    .X(net486));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input487 (.A(net1406),
    .X(net487));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input488 (.A(net1434),
    .X(net488));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input489 (.A(net1560),
    .X(net489));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input490 (.A(net1411),
    .X(net490));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input491 (.A(net1410),
    .X(net491));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input492 (.A(net1428),
    .X(net492));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input493 (.A(net1385),
    .X(net493));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input494 (.A(net1375),
    .X(net494));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input495 (.A(net1349),
    .X(net495));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input496 (.A(net1352),
    .X(net496));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input497 (.A(net1383),
    .X(net497));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input498 (.A(net1369),
    .X(net498));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input499 (.A(net1361),
    .X(net499));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input500 (.A(net1611),
    .X(net500));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input501 (.A(net1357),
    .X(net501));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input502 (.A(net1365),
    .X(net502));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input503 (.A(net1364),
    .X(net503));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input504 (.A(net1353),
    .X(net504));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input505 (.A(net1360),
    .X(net505));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input506 (.A(net1398),
    .X(net506));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input507 (.A(net1359),
    .X(net507));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input508 (.A(net1362),
    .X(net508));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input509 (.A(net1371),
    .X(net509));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input510 (.A(net1378),
    .X(net510));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input511 (.A(net1515),
    .X(net511));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input512 (.A(net1380),
    .X(net512));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input513 (.A(net1386),
    .X(net513));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input514 (.A(net1536),
    .X(net514));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input515 (.A(net1356),
    .X(net515));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input516 (.A(src_rdata[84]),
    .X(net516));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input517 (.A(net1487),
    .X(net517));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input518 (.A(net1390),
    .X(net518));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input519 (.A(net1454),
    .X(net519));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input520 (.A(net1397),
    .X(net520));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input521 (.A(src_rdata[89]),
    .X(net521));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input522 (.A(net1594),
    .X(net522));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input523 (.A(net1368),
    .X(net523));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input524 (.A(net1355),
    .X(net524));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input525 (.A(net1363),
    .X(net525));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input526 (.A(net1350),
    .X(net526));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input527 (.A(net1358),
    .X(net527));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input528 (.A(net1419),
    .X(net528));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input529 (.A(src_rdata[96]),
    .X(net529));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input530 (.A(net1447),
    .X(net530));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input531 (.A(net1478),
    .X(net531));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input532 (.A(src_rdata[99]),
    .X(net532));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input533 (.A(net1538),
    .X(net533));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input534 (.A(src_rvalid[0]),
    .X(net534));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input535 (.A(src_rvalid[1]),
    .X(net535));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input536 (.A(src_rvalid[2]),
    .X(net536));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input537 (.A(src_rvalid[3]),
    .X(net537));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output538 (.A(net538),
    .X(channel_busy[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output539 (.A(net539),
    .X(channel_busy[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output540 (.A(net540),
    .X(channel_busy[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output541 (.A(net541),
    .X(channel_busy[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output542 (.A(net542),
    .X(channel_done[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output543 (.A(net543),
    .X(channel_done[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output544 (.A(net544),
    .X(channel_done[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output545 (.A(net545),
    .X(channel_done[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output546 (.A(net546),
    .X(channel_error[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output547 (.A(net547),
    .X(channel_error[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output548 (.A(net548),
    .X(channel_error[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output549 (.A(net549),
    .X(channel_error[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output550 (.A(net550),
    .X(debug_active_channels[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output551 (.A(net551),
    .X(debug_active_channels[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output552 (.A(net552),
    .X(debug_active_channels[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output553 (.A(net553),
    .X(debug_active_channels[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output554 (.A(net554),
    .X(debug_channel_state[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output555 (.A(net555),
    .X(debug_channel_state[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output556 (.A(net556),
    .X(debug_channel_state[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output557 (.A(net557),
    .X(debug_channel_state[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output558 (.A(net558),
    .X(debug_channel_state[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output559 (.A(net1273),
    .X(debug_channel_state[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output560 (.A(net1272),
    .X(debug_channel_state[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output561 (.A(net1271),
    .X(debug_channel_state[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output562 (.A(net562),
    .X(debug_channel_state[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output563 (.A(net563),
    .X(debug_channel_state[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output564 (.A(net564),
    .X(debug_channel_state[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output565 (.A(net565),
    .X(debug_channel_state[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output566 (.A(net566),
    .X(debug_has_active_channels));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output567 (.A(net567),
    .X(debug_transfer_count[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output568 (.A(net568),
    .X(debug_transfer_count[100]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output569 (.A(net569),
    .X(debug_transfer_count[101]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output570 (.A(net570),
    .X(debug_transfer_count[102]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output571 (.A(net571),
    .X(debug_transfer_count[103]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output572 (.A(net572),
    .X(debug_transfer_count[104]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output573 (.A(net573),
    .X(debug_transfer_count[105]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output574 (.A(net574),
    .X(debug_transfer_count[106]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output575 (.A(net575),
    .X(debug_transfer_count[107]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output576 (.A(net576),
    .X(debug_transfer_count[108]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output577 (.A(net577),
    .X(debug_transfer_count[109]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output578 (.A(net578),
    .X(debug_transfer_count[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output579 (.A(net579),
    .X(debug_transfer_count[110]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output580 (.A(net580),
    .X(debug_transfer_count[111]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output581 (.A(net581),
    .X(debug_transfer_count[112]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output582 (.A(net582),
    .X(debug_transfer_count[113]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output583 (.A(net583),
    .X(debug_transfer_count[114]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output584 (.A(net584),
    .X(debug_transfer_count[115]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output585 (.A(net585),
    .X(debug_transfer_count[116]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output586 (.A(net586),
    .X(debug_transfer_count[117]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output587 (.A(net587),
    .X(debug_transfer_count[118]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output588 (.A(net588),
    .X(debug_transfer_count[119]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output589 (.A(net589),
    .X(debug_transfer_count[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output590 (.A(net590),
    .X(debug_transfer_count[120]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output591 (.A(net591),
    .X(debug_transfer_count[121]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output592 (.A(net592),
    .X(debug_transfer_count[122]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output593 (.A(net593),
    .X(debug_transfer_count[123]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output594 (.A(net594),
    .X(debug_transfer_count[124]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output595 (.A(net595),
    .X(debug_transfer_count[125]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output596 (.A(net596),
    .X(debug_transfer_count[126]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output597 (.A(net597),
    .X(debug_transfer_count[127]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output598 (.A(net598),
    .X(debug_transfer_count[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output599 (.A(net599),
    .X(debug_transfer_count[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output600 (.A(net600),
    .X(debug_transfer_count[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output601 (.A(net601),
    .X(debug_transfer_count[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output602 (.A(net602),
    .X(debug_transfer_count[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output603 (.A(net603),
    .X(debug_transfer_count[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output604 (.A(net604),
    .X(debug_transfer_count[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output605 (.A(net605),
    .X(debug_transfer_count[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output606 (.A(net606),
    .X(debug_transfer_count[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output607 (.A(net607),
    .X(debug_transfer_count[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output608 (.A(net608),
    .X(debug_transfer_count[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output609 (.A(net609),
    .X(debug_transfer_count[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output610 (.A(net610),
    .X(debug_transfer_count[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output611 (.A(net611),
    .X(debug_transfer_count[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output612 (.A(net612),
    .X(debug_transfer_count[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output613 (.A(net613),
    .X(debug_transfer_count[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output614 (.A(net614),
    .X(debug_transfer_count[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output615 (.A(net615),
    .X(debug_transfer_count[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output616 (.A(net616),
    .X(debug_transfer_count[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output617 (.A(net617),
    .X(debug_transfer_count[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output618 (.A(net618),
    .X(debug_transfer_count[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output619 (.A(net619),
    .X(debug_transfer_count[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output620 (.A(net620),
    .X(debug_transfer_count[32]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output621 (.A(net621),
    .X(debug_transfer_count[33]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output622 (.A(net622),
    .X(debug_transfer_count[34]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output623 (.A(net623),
    .X(debug_transfer_count[35]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output624 (.A(net624),
    .X(debug_transfer_count[36]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output625 (.A(net625),
    .X(debug_transfer_count[37]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output626 (.A(net626),
    .X(debug_transfer_count[38]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output627 (.A(net627),
    .X(debug_transfer_count[39]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output628 (.A(net628),
    .X(debug_transfer_count[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output629 (.A(net629),
    .X(debug_transfer_count[40]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output630 (.A(net630),
    .X(debug_transfer_count[41]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output631 (.A(net631),
    .X(debug_transfer_count[42]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output632 (.A(net632),
    .X(debug_transfer_count[43]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output633 (.A(net633),
    .X(debug_transfer_count[44]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output634 (.A(net634),
    .X(debug_transfer_count[45]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output635 (.A(net635),
    .X(debug_transfer_count[46]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output636 (.A(net636),
    .X(debug_transfer_count[47]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output637 (.A(net637),
    .X(debug_transfer_count[48]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output638 (.A(net638),
    .X(debug_transfer_count[49]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output639 (.A(net639),
    .X(debug_transfer_count[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output640 (.A(net640),
    .X(debug_transfer_count[50]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output641 (.A(net641),
    .X(debug_transfer_count[51]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output642 (.A(net642),
    .X(debug_transfer_count[52]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output643 (.A(net643),
    .X(debug_transfer_count[53]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output644 (.A(net644),
    .X(debug_transfer_count[54]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output645 (.A(net645),
    .X(debug_transfer_count[55]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output646 (.A(net646),
    .X(debug_transfer_count[56]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output647 (.A(net647),
    .X(debug_transfer_count[57]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output648 (.A(net648),
    .X(debug_transfer_count[58]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output649 (.A(net649),
    .X(debug_transfer_count[59]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output650 (.A(net650),
    .X(debug_transfer_count[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output651 (.A(net651),
    .X(debug_transfer_count[60]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output652 (.A(net652),
    .X(debug_transfer_count[61]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output653 (.A(net653),
    .X(debug_transfer_count[62]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output654 (.A(net654),
    .X(debug_transfer_count[63]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output655 (.A(net655),
    .X(debug_transfer_count[64]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output656 (.A(net656),
    .X(debug_transfer_count[65]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output657 (.A(net657),
    .X(debug_transfer_count[66]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output658 (.A(net658),
    .X(debug_transfer_count[67]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output659 (.A(net659),
    .X(debug_transfer_count[68]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output660 (.A(net660),
    .X(debug_transfer_count[69]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output661 (.A(net661),
    .X(debug_transfer_count[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output662 (.A(net662),
    .X(debug_transfer_count[70]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output663 (.A(net1270),
    .X(debug_transfer_count[71]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output664 (.A(net664),
    .X(debug_transfer_count[72]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output665 (.A(net665),
    .X(debug_transfer_count[73]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output666 (.A(net666),
    .X(debug_transfer_count[74]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output667 (.A(net667),
    .X(debug_transfer_count[75]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output668 (.A(net668),
    .X(debug_transfer_count[76]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output669 (.A(net669),
    .X(debug_transfer_count[77]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output670 (.A(net670),
    .X(debug_transfer_count[78]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output671 (.A(net671),
    .X(debug_transfer_count[79]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output672 (.A(net672),
    .X(debug_transfer_count[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output673 (.A(net673),
    .X(debug_transfer_count[80]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output674 (.A(net674),
    .X(debug_transfer_count[81]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output675 (.A(net675),
    .X(debug_transfer_count[82]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output676 (.A(net676),
    .X(debug_transfer_count[83]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output677 (.A(net677),
    .X(debug_transfer_count[84]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output678 (.A(net678),
    .X(debug_transfer_count[85]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output679 (.A(net679),
    .X(debug_transfer_count[86]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output680 (.A(net680),
    .X(debug_transfer_count[87]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output681 (.A(net681),
    .X(debug_transfer_count[88]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output682 (.A(net682),
    .X(debug_transfer_count[89]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output683 (.A(net683),
    .X(debug_transfer_count[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output684 (.A(net684),
    .X(debug_transfer_count[90]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output685 (.A(net685),
    .X(debug_transfer_count[91]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output686 (.A(net686),
    .X(debug_transfer_count[92]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output687 (.A(net687),
    .X(debug_transfer_count[93]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output688 (.A(net688),
    .X(debug_transfer_count[94]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output689 (.A(net689),
    .X(debug_transfer_count[95]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output690 (.A(net690),
    .X(debug_transfer_count[96]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output691 (.A(net691),
    .X(debug_transfer_count[97]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output692 (.A(net692),
    .X(debug_transfer_count[98]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output693 (.A(net693),
    .X(debug_transfer_count[99]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output694 (.A(net694),
    .X(debug_transfer_count[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output695 (.A(net695),
    .X(dst_addr[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output696 (.A(net696),
    .X(dst_addr[100]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output697 (.A(net697),
    .X(dst_addr[101]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output698 (.A(net698),
    .X(dst_addr[102]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output699 (.A(net699),
    .X(dst_addr[103]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output700 (.A(net700),
    .X(dst_addr[104]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output701 (.A(net701),
    .X(dst_addr[105]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output702 (.A(net702),
    .X(dst_addr[106]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output703 (.A(net703),
    .X(dst_addr[107]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output704 (.A(net704),
    .X(dst_addr[108]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output705 (.A(net705),
    .X(dst_addr[109]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output706 (.A(net706),
    .X(dst_addr[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output707 (.A(net707),
    .X(dst_addr[110]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output708 (.A(net708),
    .X(dst_addr[111]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output709 (.A(net709),
    .X(dst_addr[112]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output710 (.A(net710),
    .X(dst_addr[113]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output711 (.A(net711),
    .X(dst_addr[114]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output712 (.A(net712),
    .X(dst_addr[115]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output713 (.A(net713),
    .X(dst_addr[116]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output714 (.A(net714),
    .X(dst_addr[117]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output715 (.A(net715),
    .X(dst_addr[118]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output716 (.A(net716),
    .X(dst_addr[119]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output717 (.A(net717),
    .X(dst_addr[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output718 (.A(net718),
    .X(dst_addr[120]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output719 (.A(net719),
    .X(dst_addr[121]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output720 (.A(net720),
    .X(dst_addr[122]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output721 (.A(net721),
    .X(dst_addr[123]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output722 (.A(net722),
    .X(dst_addr[124]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output723 (.A(net723),
    .X(dst_addr[125]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output724 (.A(net724),
    .X(dst_addr[126]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output725 (.A(net725),
    .X(dst_addr[127]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output726 (.A(net726),
    .X(dst_addr[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output727 (.A(net727),
    .X(dst_addr[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output728 (.A(net728),
    .X(dst_addr[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output729 (.A(net729),
    .X(dst_addr[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output730 (.A(net730),
    .X(dst_addr[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output731 (.A(net731),
    .X(dst_addr[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output732 (.A(net732),
    .X(dst_addr[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output733 (.A(net733),
    .X(dst_addr[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output734 (.A(net734),
    .X(dst_addr[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output735 (.A(net735),
    .X(dst_addr[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output736 (.A(net736),
    .X(dst_addr[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output737 (.A(net737),
    .X(dst_addr[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output738 (.A(net738),
    .X(dst_addr[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output739 (.A(net739),
    .X(dst_addr[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output740 (.A(net740),
    .X(dst_addr[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output741 (.A(net741),
    .X(dst_addr[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output742 (.A(net742),
    .X(dst_addr[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output743 (.A(net743),
    .X(dst_addr[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output744 (.A(net744),
    .X(dst_addr[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output745 (.A(net745),
    .X(dst_addr[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output746 (.A(net746),
    .X(dst_addr[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output747 (.A(net747),
    .X(dst_addr[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output748 (.A(net748),
    .X(dst_addr[32]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output749 (.A(net749),
    .X(dst_addr[33]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output750 (.A(net750),
    .X(dst_addr[34]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output751 (.A(net751),
    .X(dst_addr[35]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output752 (.A(net752),
    .X(dst_addr[36]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output753 (.A(net753),
    .X(dst_addr[37]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output754 (.A(net754),
    .X(dst_addr[38]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output755 (.A(net755),
    .X(dst_addr[39]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output756 (.A(net756),
    .X(dst_addr[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output757 (.A(net757),
    .X(dst_addr[40]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output758 (.A(net758),
    .X(dst_addr[41]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output759 (.A(net759),
    .X(dst_addr[42]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output760 (.A(net760),
    .X(dst_addr[43]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output761 (.A(net761),
    .X(dst_addr[44]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output762 (.A(net762),
    .X(dst_addr[45]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output763 (.A(net763),
    .X(dst_addr[46]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output764 (.A(net764),
    .X(dst_addr[47]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output765 (.A(net765),
    .X(dst_addr[48]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output766 (.A(net766),
    .X(dst_addr[49]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output767 (.A(net767),
    .X(dst_addr[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output768 (.A(net768),
    .X(dst_addr[50]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output769 (.A(net769),
    .X(dst_addr[51]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output770 (.A(net770),
    .X(dst_addr[52]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output771 (.A(net771),
    .X(dst_addr[53]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output772 (.A(net772),
    .X(dst_addr[54]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output773 (.A(net773),
    .X(dst_addr[55]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output774 (.A(net774),
    .X(dst_addr[56]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output775 (.A(net775),
    .X(dst_addr[57]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output776 (.A(net776),
    .X(dst_addr[58]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output777 (.A(net777),
    .X(dst_addr[59]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output778 (.A(net778),
    .X(dst_addr[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output779 (.A(net779),
    .X(dst_addr[60]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output780 (.A(net780),
    .X(dst_addr[61]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output781 (.A(net781),
    .X(dst_addr[62]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output782 (.A(net782),
    .X(dst_addr[63]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output783 (.A(net783),
    .X(dst_addr[64]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output784 (.A(net784),
    .X(dst_addr[65]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output785 (.A(net785),
    .X(dst_addr[66]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output786 (.A(net786),
    .X(dst_addr[67]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output787 (.A(net787),
    .X(dst_addr[68]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output788 (.A(net788),
    .X(dst_addr[69]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output789 (.A(net789),
    .X(dst_addr[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output790 (.A(net790),
    .X(dst_addr[70]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output791 (.A(net791),
    .X(dst_addr[71]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output792 (.A(net792),
    .X(dst_addr[72]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output793 (.A(net793),
    .X(dst_addr[73]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output794 (.A(net794),
    .X(dst_addr[74]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output795 (.A(net795),
    .X(dst_addr[75]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output796 (.A(net796),
    .X(dst_addr[76]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output797 (.A(net797),
    .X(dst_addr[77]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output798 (.A(net798),
    .X(dst_addr[78]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output799 (.A(net799),
    .X(dst_addr[79]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output800 (.A(net800),
    .X(dst_addr[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output801 (.A(net801),
    .X(dst_addr[80]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output802 (.A(net802),
    .X(dst_addr[81]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output803 (.A(net803),
    .X(dst_addr[82]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output804 (.A(net804),
    .X(dst_addr[83]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output805 (.A(net805),
    .X(dst_addr[84]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output806 (.A(net806),
    .X(dst_addr[85]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output807 (.A(net807),
    .X(dst_addr[86]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output808 (.A(net808),
    .X(dst_addr[87]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output809 (.A(net809),
    .X(dst_addr[88]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output810 (.A(net810),
    .X(dst_addr[89]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output811 (.A(net811),
    .X(dst_addr[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output812 (.A(net812),
    .X(dst_addr[90]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output813 (.A(net813),
    .X(dst_addr[91]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output814 (.A(net814),
    .X(dst_addr[92]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output815 (.A(net815),
    .X(dst_addr[93]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output816 (.A(net816),
    .X(dst_addr[94]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output817 (.A(net817),
    .X(dst_addr[95]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output818 (.A(net818),
    .X(dst_addr[96]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output819 (.A(net819),
    .X(dst_addr[97]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output820 (.A(net820),
    .X(dst_addr[98]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output821 (.A(net821),
    .X(dst_addr[99]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output822 (.A(net822),
    .X(dst_addr[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output823 (.A(net823),
    .X(dst_wdata[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output824 (.A(net824),
    .X(dst_wdata[100]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output825 (.A(net825),
    .X(dst_wdata[101]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output826 (.A(net826),
    .X(dst_wdata[102]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output827 (.A(net827),
    .X(dst_wdata[103]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output828 (.A(net828),
    .X(dst_wdata[104]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output829 (.A(net829),
    .X(dst_wdata[105]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output830 (.A(net830),
    .X(dst_wdata[106]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output831 (.A(net831),
    .X(dst_wdata[107]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output832 (.A(net832),
    .X(dst_wdata[108]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output833 (.A(net833),
    .X(dst_wdata[109]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output834 (.A(net834),
    .X(dst_wdata[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output835 (.A(net835),
    .X(dst_wdata[110]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output836 (.A(net836),
    .X(dst_wdata[111]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output837 (.A(net837),
    .X(dst_wdata[112]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output838 (.A(net838),
    .X(dst_wdata[113]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output839 (.A(net839),
    .X(dst_wdata[114]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output840 (.A(net840),
    .X(dst_wdata[115]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output841 (.A(net841),
    .X(dst_wdata[116]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output842 (.A(net842),
    .X(dst_wdata[117]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output843 (.A(net843),
    .X(dst_wdata[118]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output844 (.A(net844),
    .X(dst_wdata[119]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output845 (.A(net845),
    .X(dst_wdata[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output846 (.A(net846),
    .X(dst_wdata[120]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output847 (.A(net847),
    .X(dst_wdata[121]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output848 (.A(net848),
    .X(dst_wdata[122]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output849 (.A(net849),
    .X(dst_wdata[123]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output850 (.A(net850),
    .X(dst_wdata[124]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output851 (.A(net851),
    .X(dst_wdata[125]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output852 (.A(net852),
    .X(dst_wdata[126]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output853 (.A(net853),
    .X(dst_wdata[127]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output854 (.A(net854),
    .X(dst_wdata[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output855 (.A(net855),
    .X(dst_wdata[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output856 (.A(net856),
    .X(dst_wdata[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output857 (.A(net857),
    .X(dst_wdata[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output858 (.A(net858),
    .X(dst_wdata[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output859 (.A(net859),
    .X(dst_wdata[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output860 (.A(net860),
    .X(dst_wdata[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output861 (.A(net861),
    .X(dst_wdata[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output862 (.A(net862),
    .X(dst_wdata[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output863 (.A(net863),
    .X(dst_wdata[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output864 (.A(net864),
    .X(dst_wdata[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output865 (.A(net865),
    .X(dst_wdata[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output866 (.A(net866),
    .X(dst_wdata[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output867 (.A(net867),
    .X(dst_wdata[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output868 (.A(net868),
    .X(dst_wdata[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output869 (.A(net869),
    .X(dst_wdata[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output870 (.A(net870),
    .X(dst_wdata[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output871 (.A(net871),
    .X(dst_wdata[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output872 (.A(net872),
    .X(dst_wdata[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output873 (.A(net873),
    .X(dst_wdata[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output874 (.A(net874),
    .X(dst_wdata[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output875 (.A(net875),
    .X(dst_wdata[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output876 (.A(net876),
    .X(dst_wdata[32]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output877 (.A(net877),
    .X(dst_wdata[33]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output878 (.A(net878),
    .X(dst_wdata[34]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output879 (.A(net879),
    .X(dst_wdata[35]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output880 (.A(net880),
    .X(dst_wdata[36]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output881 (.A(net881),
    .X(dst_wdata[37]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output882 (.A(net882),
    .X(dst_wdata[38]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output883 (.A(net883),
    .X(dst_wdata[39]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output884 (.A(net884),
    .X(dst_wdata[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output885 (.A(net885),
    .X(dst_wdata[40]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output886 (.A(net886),
    .X(dst_wdata[41]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output887 (.A(net887),
    .X(dst_wdata[42]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output888 (.A(net888),
    .X(dst_wdata[43]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output889 (.A(net889),
    .X(dst_wdata[44]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output890 (.A(net890),
    .X(dst_wdata[45]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output891 (.A(net891),
    .X(dst_wdata[46]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output892 (.A(net892),
    .X(dst_wdata[47]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output893 (.A(net893),
    .X(dst_wdata[48]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output894 (.A(net894),
    .X(dst_wdata[49]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output895 (.A(net895),
    .X(dst_wdata[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output896 (.A(net896),
    .X(dst_wdata[50]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output897 (.A(net897),
    .X(dst_wdata[51]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output898 (.A(net898),
    .X(dst_wdata[52]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output899 (.A(net899),
    .X(dst_wdata[53]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output900 (.A(net900),
    .X(dst_wdata[54]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output901 (.A(net901),
    .X(dst_wdata[55]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output902 (.A(net902),
    .X(dst_wdata[56]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output903 (.A(net903),
    .X(dst_wdata[57]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output904 (.A(net904),
    .X(dst_wdata[58]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output905 (.A(net905),
    .X(dst_wdata[59]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output906 (.A(net906),
    .X(dst_wdata[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output907 (.A(net907),
    .X(dst_wdata[60]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output908 (.A(net908),
    .X(dst_wdata[61]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output909 (.A(net909),
    .X(dst_wdata[62]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output910 (.A(net910),
    .X(dst_wdata[63]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output911 (.A(net911),
    .X(dst_wdata[64]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output912 (.A(net912),
    .X(dst_wdata[65]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output913 (.A(net913),
    .X(dst_wdata[66]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output914 (.A(net914),
    .X(dst_wdata[67]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output915 (.A(net915),
    .X(dst_wdata[68]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output916 (.A(net916),
    .X(dst_wdata[69]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output917 (.A(net917),
    .X(dst_wdata[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output918 (.A(net918),
    .X(dst_wdata[70]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output919 (.A(net919),
    .X(dst_wdata[71]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output920 (.A(net920),
    .X(dst_wdata[72]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output921 (.A(net921),
    .X(dst_wdata[73]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output922 (.A(net922),
    .X(dst_wdata[74]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output923 (.A(net923),
    .X(dst_wdata[75]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output924 (.A(net924),
    .X(dst_wdata[76]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output925 (.A(net925),
    .X(dst_wdata[77]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output926 (.A(net926),
    .X(dst_wdata[78]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output927 (.A(net927),
    .X(dst_wdata[79]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output928 (.A(net928),
    .X(dst_wdata[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output929 (.A(net929),
    .X(dst_wdata[80]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output930 (.A(net930),
    .X(dst_wdata[81]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output931 (.A(net931),
    .X(dst_wdata[82]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output932 (.A(net932),
    .X(dst_wdata[83]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output933 (.A(net933),
    .X(dst_wdata[84]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output934 (.A(net934),
    .X(dst_wdata[85]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output935 (.A(net935),
    .X(dst_wdata[86]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output936 (.A(net936),
    .X(dst_wdata[87]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output937 (.A(net937),
    .X(dst_wdata[88]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output938 (.A(net938),
    .X(dst_wdata[89]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output939 (.A(net939),
    .X(dst_wdata[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output940 (.A(net940),
    .X(dst_wdata[90]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output941 (.A(net941),
    .X(dst_wdata[91]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output942 (.A(net942),
    .X(dst_wdata[92]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output943 (.A(net943),
    .X(dst_wdata[93]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output944 (.A(net944),
    .X(dst_wdata[94]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output945 (.A(net945),
    .X(dst_wdata[95]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output946 (.A(net946),
    .X(dst_wdata[96]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output947 (.A(net947),
    .X(dst_wdata[97]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output948 (.A(net948),
    .X(dst_wdata[98]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output949 (.A(net949),
    .X(dst_wdata[99]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output950 (.A(net950),
    .X(dst_wdata[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output951 (.A(net951),
    .X(dst_write[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output952 (.A(net952),
    .X(dst_write[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output953 (.A(net953),
    .X(dst_write[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output954 (.A(net954),
    .X(dst_write[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output955 (.A(net964),
    .X(dst_wstrb[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output956 (.A(net957),
    .X(dst_wstrb[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output957 (.A(net957),
    .X(dst_wstrb[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output958 (.A(net961),
    .X(dst_wstrb[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output959 (.A(net961),
    .X(dst_wstrb[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output960 (.A(net961),
    .X(dst_wstrb[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output961 (.A(net961),
    .X(dst_wstrb[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output962 (.A(net964),
    .X(dst_wstrb[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output963 (.A(net964),
    .X(dst_wstrb[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output964 (.A(net964),
    .X(dst_wstrb[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output965 (.A(net968),
    .X(dst_wstrb[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output966 (.A(net968),
    .X(dst_wstrb[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output967 (.A(net968),
    .X(dst_wstrb[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output968 (.A(net968),
    .X(dst_wstrb[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output969 (.A(net957),
    .X(dst_wstrb[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output970 (.A(net957),
    .X(dst_wstrb[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output971 (.A(net971),
    .X(src_addr[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output972 (.A(net972),
    .X(src_addr[100]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output973 (.A(net973),
    .X(src_addr[101]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output974 (.A(net974),
    .X(src_addr[102]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output975 (.A(net975),
    .X(src_addr[103]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output976 (.A(net976),
    .X(src_addr[104]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output977 (.A(net977),
    .X(src_addr[105]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output978 (.A(net978),
    .X(src_addr[106]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output979 (.A(net979),
    .X(src_addr[107]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output980 (.A(net980),
    .X(src_addr[108]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output981 (.A(net981),
    .X(src_addr[109]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output982 (.A(net982),
    .X(src_addr[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output983 (.A(net983),
    .X(src_addr[110]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output984 (.A(net984),
    .X(src_addr[111]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output985 (.A(net985),
    .X(src_addr[112]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output986 (.A(net986),
    .X(src_addr[113]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output987 (.A(net987),
    .X(src_addr[114]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output988 (.A(net988),
    .X(src_addr[115]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output989 (.A(net989),
    .X(src_addr[116]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output990 (.A(net990),
    .X(src_addr[117]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output991 (.A(net991),
    .X(src_addr[118]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output992 (.A(net992),
    .X(src_addr[119]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output993 (.A(net993),
    .X(src_addr[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output994 (.A(net994),
    .X(src_addr[120]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output995 (.A(net995),
    .X(src_addr[121]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output996 (.A(net996),
    .X(src_addr[122]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output997 (.A(net997),
    .X(src_addr[123]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output998 (.A(net998),
    .X(src_addr[124]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output999 (.A(net999),
    .X(src_addr[125]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1000 (.A(net1000),
    .X(src_addr[126]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1001 (.A(net1001),
    .X(src_addr[127]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1002 (.A(net1002),
    .X(src_addr[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1003 (.A(net1003),
    .X(src_addr[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1004 (.A(net1004),
    .X(src_addr[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1005 (.A(net1005),
    .X(src_addr[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1006 (.A(net1006),
    .X(src_addr[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1007 (.A(net1007),
    .X(src_addr[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1008 (.A(net1008),
    .X(src_addr[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1009 (.A(net1009),
    .X(src_addr[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1010 (.A(net1010),
    .X(src_addr[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1011 (.A(net1011),
    .X(src_addr[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1012 (.A(net1012),
    .X(src_addr[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1013 (.A(net1013),
    .X(src_addr[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1014 (.A(net1014),
    .X(src_addr[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1015 (.A(net1015),
    .X(src_addr[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1016 (.A(net1016),
    .X(src_addr[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1017 (.A(net1017),
    .X(src_addr[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1018 (.A(net1018),
    .X(src_addr[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1019 (.A(net1019),
    .X(src_addr[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1020 (.A(net1020),
    .X(src_addr[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1021 (.A(net1021),
    .X(src_addr[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1022 (.A(net1022),
    .X(src_addr[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1023 (.A(net1023),
    .X(src_addr[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1024 (.A(net1024),
    .X(src_addr[32]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1025 (.A(net1025),
    .X(src_addr[33]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1026 (.A(net1026),
    .X(src_addr[34]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1027 (.A(net1027),
    .X(src_addr[35]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1028 (.A(net1028),
    .X(src_addr[36]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1029 (.A(net1029),
    .X(src_addr[37]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1030 (.A(net1030),
    .X(src_addr[38]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1031 (.A(net1031),
    .X(src_addr[39]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1032 (.A(net1032),
    .X(src_addr[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1033 (.A(net1033),
    .X(src_addr[40]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1034 (.A(net1034),
    .X(src_addr[41]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1035 (.A(net1035),
    .X(src_addr[42]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1036 (.A(net1036),
    .X(src_addr[43]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1037 (.A(net1037),
    .X(src_addr[44]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1038 (.A(net1038),
    .X(src_addr[45]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1039 (.A(net1039),
    .X(src_addr[46]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1040 (.A(net1040),
    .X(src_addr[47]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1041 (.A(net1041),
    .X(src_addr[48]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1042 (.A(net1042),
    .X(src_addr[49]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1043 (.A(net1043),
    .X(src_addr[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1044 (.A(net1044),
    .X(src_addr[50]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1045 (.A(net1045),
    .X(src_addr[51]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1046 (.A(net1046),
    .X(src_addr[52]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1047 (.A(net1047),
    .X(src_addr[53]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1048 (.A(net1048),
    .X(src_addr[54]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1049 (.A(net1049),
    .X(src_addr[55]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1050 (.A(net1050),
    .X(src_addr[56]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1051 (.A(net1051),
    .X(src_addr[57]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1052 (.A(net1052),
    .X(src_addr[58]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1053 (.A(net1053),
    .X(src_addr[59]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1054 (.A(net1054),
    .X(src_addr[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1055 (.A(net1055),
    .X(src_addr[60]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1056 (.A(net1056),
    .X(src_addr[61]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1057 (.A(net1057),
    .X(src_addr[62]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1058 (.A(net1058),
    .X(src_addr[63]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1059 (.A(net1059),
    .X(src_addr[64]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1060 (.A(net1060),
    .X(src_addr[65]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1061 (.A(net1061),
    .X(src_addr[66]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1062 (.A(net1062),
    .X(src_addr[67]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1063 (.A(net1063),
    .X(src_addr[68]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1064 (.A(net1064),
    .X(src_addr[69]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1065 (.A(net1065),
    .X(src_addr[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1066 (.A(net1066),
    .X(src_addr[70]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1067 (.A(net1067),
    .X(src_addr[71]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1068 (.A(net1068),
    .X(src_addr[72]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1069 (.A(net1069),
    .X(src_addr[73]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1070 (.A(net1070),
    .X(src_addr[74]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1071 (.A(net1071),
    .X(src_addr[75]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1072 (.A(net1072),
    .X(src_addr[76]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1073 (.A(net1073),
    .X(src_addr[77]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1074 (.A(net1074),
    .X(src_addr[78]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1075 (.A(net1075),
    .X(src_addr[79]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1076 (.A(net1076),
    .X(src_addr[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1077 (.A(net1077),
    .X(src_addr[80]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1078 (.A(net1078),
    .X(src_addr[81]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1079 (.A(net1079),
    .X(src_addr[82]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1080 (.A(net1080),
    .X(src_addr[83]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1081 (.A(net1081),
    .X(src_addr[84]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1082 (.A(net1082),
    .X(src_addr[85]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1083 (.A(net1083),
    .X(src_addr[86]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1084 (.A(net1084),
    .X(src_addr[87]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1085 (.A(net1085),
    .X(src_addr[88]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1086 (.A(net1086),
    .X(src_addr[89]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1087 (.A(net1087),
    .X(src_addr[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1088 (.A(net1088),
    .X(src_addr[90]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1089 (.A(net1089),
    .X(src_addr[91]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1090 (.A(net1090),
    .X(src_addr[92]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1091 (.A(net1091),
    .X(src_addr[93]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1092 (.A(net1092),
    .X(src_addr[94]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1093 (.A(net1093),
    .X(src_addr[95]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1094 (.A(net1094),
    .X(src_addr[96]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1095 (.A(net1095),
    .X(src_addr[97]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1096 (.A(net1096),
    .X(src_addr[98]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1097 (.A(net1097),
    .X(src_addr[99]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1098 (.A(net1098),
    .X(src_addr[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1099 (.A(net1099),
    .X(src_read[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1100 (.A(net1100),
    .X(src_read[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1101 (.A(net1101),
    .X(src_read[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1102 (.A(net1102),
    .X(src_read[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1103 (.A(net1103),
    .X(src_rready[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1104 (.A(net1104),
    .X(src_rready[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1105 (.A(net1105),
    .X(src_rready[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output1106 (.A(net1106),
    .X(src_rready[3]));
 sky130_fd_sc_hd__buf_12 place1283 (.A(net405),
    .X(net1283));
 sky130_fd_sc_hd__buf_4 place1239 (.A(_3049_),
    .X(net1239));
 sky130_fd_sc_hd__buf_4 place1237 (.A(_3307_),
    .X(net1237));
 sky130_fd_sc_hd__buf_4 place1238 (.A(_3292_),
    .X(net1238));
 sky130_fd_sc_hd__buf_4 place1259 (.A(net1258),
    .X(net1259));
 sky130_fd_sc_hd__buf_4 place1258 (.A(_3298_),
    .X(net1258));
 sky130_fd_sc_hd__buf_4 place1247 (.A(_1733_),
    .X(net1247));
 sky130_fd_sc_hd__buf_4 place1249 (.A(_1604_),
    .X(net1249));
 sky130_fd_sc_hd__buf_4 place1252 (.A(_1459_),
    .X(net1252));
 sky130_fd_sc_hd__buf_4 place1254 (.A(_1451_),
    .X(net1254));
 sky130_fd_sc_hd__buf_4 place1262 (.A(_3274_),
    .X(net1262));
 sky130_fd_sc_hd__buf_4 place1260 (.A(_3283_),
    .X(net1260));
 sky130_fd_sc_hd__buf_4 place1272 (.A(net560),
    .X(net1272));
 sky130_fd_sc_hd__buf_4 place1273 (.A(net559),
    .X(net1273));
 sky130_fd_sc_hd__buf_4 place1261 (.A(_3274_),
    .X(net1261));
 sky130_fd_sc_hd__buf_4 place1275 (.A(net405),
    .X(net1275));
 sky130_fd_sc_hd__buf_4 place1263 (.A(_1872_),
    .X(net1263));
 sky130_fd_sc_hd__buf_4 place1268 (.A(_1470_),
    .X(net1268));
 sky130_fd_sc_hd__buf_4 place1264 (.A(_1741_),
    .X(net1264));
 sky130_fd_sc_hd__buf_4 place1279 (.A(net1277),
    .X(net1279));
 sky130_fd_sc_hd__buf_4 place1265 (.A(_1736_),
    .X(net1265));
 sky130_fd_sc_hd__buf_4 place1267 (.A(_1474_),
    .X(net1267));
 sky130_fd_sc_hd__buf_12 place1278 (.A(net1277),
    .X(net1278));
 sky130_fd_sc_hd__buf_4 place1266 (.A(_1607_),
    .X(net1266));
 sky130_fd_sc_hd__buf_4 place1269 (.A(_1463_),
    .X(net1269));
 sky130_fd_sc_hd__buf_4 place1270 (.A(net663),
    .X(net1270));
 sky130_fd_sc_hd__buf_12 place1277 (.A(net405),
    .X(net1277));
 sky130_fd_sc_hd__buf_4 place1276 (.A(net405),
    .X(net1276));
 sky130_fd_sc_hd__buf_4 place1227 (.A(_3268_),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__buf_12 place1292 (.A(net1284),
    .X(net1292));
 sky130_fd_sc_hd__buf_12 place1291 (.A(net1284),
    .X(net1291));
 sky130_fd_sc_hd__buf_4 place1228 (.A(_2441_),
    .X(net1228));
 sky130_fd_sc_hd__buf_4 place1290 (.A(net1284),
    .X(net1290));
 sky130_fd_sc_hd__buf_4 place1289 (.A(net1284),
    .X(net1289));
 sky130_fd_sc_hd__buf_4 place1288 (.A(net1284),
    .X(net1288));
 sky130_fd_sc_hd__buf_4 place1287 (.A(net1284),
    .X(net1287));
 sky130_fd_sc_hd__buf_4 place1286 (.A(net1284),
    .X(net1286));
 sky130_fd_sc_hd__buf_4 place1229 (.A(_2444_),
    .X(net1229));
 sky130_fd_sc_hd__buf_4 place1285 (.A(net1284),
    .X(net1285));
 sky130_fd_sc_hd__buf_4 place1230 (.A(_2896_),
    .X(net1230));
 sky130_fd_sc_hd__buf_12 place1284 (.A(net405),
    .X(net1284));
 sky130_fd_sc_hd__buf_4 place1282 (.A(net1280),
    .X(net1282));
 sky130_fd_sc_hd__buf_4 place1231 (.A(_2783_),
    .X(net1231));
 sky130_fd_sc_hd__buf_4 place1281 (.A(net1280),
    .X(net1281));
 sky130_fd_sc_hd__buf_4 place1232 (.A(_2745_),
    .X(net1232));
 sky130_fd_sc_hd__buf_4 place1280 (.A(net405),
    .X(net1280));
 sky130_fd_sc_hd__buf_4 place1233 (.A(_2610_),
    .X(net1233));
 sky130_fd_sc_hd__buf_4 place1234 (.A(_2468_),
    .X(net1234));
 sky130_fd_sc_hd__buf_4 place1235 (.A(_3392_),
    .X(net1235));
 sky130_fd_sc_hd__buf_4 place1236 (.A(_3375_),
    .X(net1236));
 sky130_fd_sc_hd__buf_4 place1240 (.A(_3035_),
    .X(net1240));
 sky130_fd_sc_hd__buf_4 place1241 (.A(_2638_),
    .X(net1241));
 sky130_fd_sc_hd__buf_4 place1243 (.A(_1880_),
    .X(net1243));
 sky130_fd_sc_hd__buf_4 place1242 (.A(_2125_),
    .X(net1242));
 sky130_fd_sc_hd__buf_4 place1244 (.A(_1866_),
    .X(net1244));
 sky130_fd_sc_hd__buf_4 place1245 (.A(_1748_),
    .X(net1245));
 sky130_fd_sc_hd__buf_4 place1246 (.A(_1733_),
    .X(net1246));
 sky130_fd_sc_hd__buf_4 place1248 (.A(_1618_),
    .X(net1248));
 sky130_fd_sc_hd__buf_4 place1250 (.A(_1473_),
    .X(net1250));
 sky130_fd_sc_hd__buf_4 place1251 (.A(_1465_),
    .X(net1251));
 sky130_fd_sc_hd__buf_4 place1253 (.A(_1454_),
    .X(net1253));
 sky130_fd_sc_hd__buf_4 place1256 (.A(_3372_),
    .X(net1256));
 sky130_fd_sc_hd__buf_4 place1255 (.A(_3372_),
    .X(net1255));
 sky130_fd_sc_hd__buf_4 place1257 (.A(_3298_),
    .X(net1257));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__buf_4 place1293 (.A(net402),
    .X(net1293));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload3 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload8 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload9 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload14 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload15 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload16 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkinv_2 clkload17 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__bufinv_16 clkload18 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__inv_8 clkload19 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload20 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload21 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload22 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload23 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkinv_4 clkload26 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__inv_8 clkload27 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__inv_8 clkload28 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__inv_8 clkload29 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_4 clkload30 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__inv_6 clkload32 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload33 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_2 clkload34 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__bufinv_16 clkload35 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__bufinv_16 clkload37 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_2 clkload38 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinv_2 clkload39 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__bufinv_16 clkload40 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload41 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload42 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__bufinv_16 clkload43 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_2 clkload44 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__bufinv_16 clkload45 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinv_4 clkload46 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__inv_6 clkload47 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__inv_6 clkload48 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__bufinv_16 clkload49 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__bufinv_16 clkload50 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinv_2 clkload51 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload52 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload53 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload54 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload55 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload56 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload57 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload58 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload59 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload60 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__inv_6 clkload61 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload62 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload63 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload64 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload65 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkinv_2 clkload66 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkinv_2 clkload67 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload68 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload69 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload70 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload71 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload72 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload73 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload74 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload75 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_2 clkload76 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload77 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload78 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload79 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkinv_4 clkload80 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkinv_4 clkload81 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__inv_6 clkload82 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkinv_2 clkload83 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload84 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkinv_2 clkload85 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload86 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload87 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__bufinv_16 clkload88 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload89 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload90 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__inv_6 clkload91 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__bufinv_16 clkload92 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload93 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__bufinv_16 clkload94 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(rst_n),
    .X(net1294));
 sky130_fd_sc_hd__buf_16 hold1295 (.A(net405),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(channel_src_addr[65]),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(channel_dst_addr[64]),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(channel_dst_addr[65]),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(channel_dst_addr[33]),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(channel_dst_addr[81]),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(channel_dst_addr[68]),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(channel_dst_addr[32]),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(channel_src_addr[32]),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(channel_src_addr[96]),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(channel_src_addr[33]),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(channel_src_addr[88]),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(channel_src_addr[94]),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(channel_src_addr[92]),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(channel_dst_addr[82]),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(channel_dst_addr[72]),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(channel_src_addr[82]),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(channel_dst_addr[92]),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(channel_dst_addr[84]),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(channel_dst_addr[88]),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(src_rdata[113]),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(channel_src_addr[74]),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(src_rdata[107]),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(channel_src_addr[95]),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(src_rdata[116]),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(src_rdata[110]),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(src_rdata[112]),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(src_rdata[120]),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(src_rdata[118]),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(src_rdata[121]),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(channel_dst_addr[83]),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(channel_src_addr[64]),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(channel_src_addr[75]),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(channel_dst_addr[93]),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(src_rdata[122]),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(channel_src_addr[97]),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(channel_src_addr[66]),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(src_rdata[117]),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(src_rdata[115]),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(src_rdata[126]),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(src_rdata[109]),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(channel_dst_addr[66]),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(src_rdata[114]),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(channel_dst_addr[96]),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(src_rdata[111]),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(channel_src_addr[80]),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(src_rdata[124]),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(channel_dst_addr[35]),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(channel_src_addr[90]),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(channel_dst_addr[77]),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(channel_dst_addr[67]),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(channel_src_addr[86]),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(src_rdata[108]),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(channel_dst_addr[97]),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(src_rdata[65]),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(src_rdata[93]),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(channel_dst_addr[98]),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(src_rdata[66]),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(src_rdata[73]),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(src_rdata[123]),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(src_rdata[91]),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(src_rdata[83]),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(src_rdata[70]),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(src_rdata[94]),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(src_rdata[76]),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(src_rdata[74]),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(src_rdata[69]),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(src_rdata[77]),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(src_rdata[92]),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(src_rdata[72]),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(src_rdata[71]),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(channel_dst_addr[42]),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(channel_src_addr[77]),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(src_rdata[90]),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(src_rdata[68]),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(channel_src_addr[27]),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(src_rdata[78]),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(channel_dst_addr[114]),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(channel_dst_addr[99]),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(channel_dst_addr[0]),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(src_rdata[64]),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(channel_dst_addr[71]),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(channel_dst_addr[75]),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(src_rdata[79]),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(channel_src_addr[43]),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(src_rdata[80]),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(channel_dst_addr[79]),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(channel_dst_addr[86]),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(src_rdata[67]),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(channel_dst_addr[127]),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(src_rdata[63]),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(src_rdata[81]),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(channel_src_addr[1]),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(src_rdata[42]),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(src_rdata[45]),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(src_rdata[86]),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(src_rdata[43]),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(channel_src_addr[111]),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(channel_dst_addr[52]),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(channel_src_addr[87]),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(src_rdata[52]),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(channel_dst_addr[78]),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(src_rdata[88]),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(src_rdata[75]),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(channel_dst_addr[76]),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(channel_src_addr[79]),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(channel_dst_addr[50]),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(channel_dst_addr[58]),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(src_rdata[125]),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(channel_dst_addr[89]),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(src_rdata[36]),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(src_rdata[58]),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(src_rdata[32]),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(src_rdata[56]),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(channel_dst_addr[80]),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(src_rdata[61]),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(src_rdata[60]),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(src_rdata[38]),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(src_rdata[57]),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(src_rdata[34]),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(src_rdata[39]),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(src_rdata[35]),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(channel_dst_addr[105]),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(channel_dst_addr[125]),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(src_rdata[95]),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(channel_src_addr[52]),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(channel_src_addr[53]),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(channel_src_addr[45]),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(channel_src_addr[106]),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(src_rdata[55]),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(src_rdata[48]),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(channel_src_addr[23]),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(channel_dst_addr[70]),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(src_rdata[62]),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(channel_src_addr[26]),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(channel_src_addr[112]),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(channel_dst_addr[85]),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(src_rdata[41]),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(channel_dst_addr[56]),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(src_rdata[59]),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(channel_src_addr[63]),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(channel_dst_addr[44]),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(channel_src_addr[109]),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(src_rdata[33]),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(channel_src_addr[123]),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(channel_src_addr[62]),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(src_rdata[105]),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(channel_src_addr[73]),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(channel_src_addr[59]),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(channel_dst_addr[124]),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(channel_src_addr[29]),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(src_rdata[15]),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(src_rdata[97]),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(src_rdata[101]),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(channel_src_addr[83]),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(channel_dst_addr[51]),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(channel_src_addr[89]),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(channel_src_addr[51]),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(channel_dst_addr[102]),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(src_rdata[87]),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(channel_src_addr[122]),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(channel_src_addr[44]),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(channel_src_addr[24]),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(channel_dst_addr[63]),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(channel_dst_addr[39]),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(src_rdata[103]),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(channel_dst_addr[49]),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(channel_src_addr[113]),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(channel_src_addr[67]),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(src_rdata[40]),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(channel_src_addr[68]),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(channel_src_addr[61]),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(channel_dst_addr[1]),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(channel_dst_addr[123]),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(channel_src_addr[49]),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(channel_dst_addr[46]),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(channel_src_addr[93]),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(channel_dst_addr[106]),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(channel_dst_addr[40]),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(channel_src_addr[48]),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(channel_src_addr[41]),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(channel_src_addr[78]),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(channel_src_addr[117]),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(src_rdata[98]),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(channel_dst_addr[59]),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(channel_src_addr[28]),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(channel_src_addr[56]),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(channel_src_addr[124]),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(channel_dst_addr[113]),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(channel_dst_addr[74]),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(channel_dst_addr[109]),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(channel_src_addr[118]),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(src_rdata[85]),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(channel_src_addr[105]),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(src_rdata[12]),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(channel_dst_addr[54]),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(channel_src_addr[121]),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(channel_dst_addr[111]),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(src_rdata[29]),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(channel_dst_addr[69]),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(src_rdata[106]),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(channel_dst_addr[126]),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(channel_dst_addr[100]),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(channel_dst_addr[108]),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(channel_dst_addr[115]),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(channel_dst_addr[60]),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(channel_dst_addr[101]),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(src_rdata[11]),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(channel_dst_addr[73]),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(channel_src_addr[69]),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(src_rdata[13]),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(src_rdata[25]),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(channel_dst_addr[104]),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(src_rdata[14]),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(channel_src_addr[25]),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(src_rdata[27]),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(src_rdata[119]),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(src_rdata[49]),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(src_rdata[50]),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(src_rdata[53]),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(src_rdata[7]),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(channel_dst_addr[87]),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(src_rdata[104]),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(channel_src_addr[107]),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(channel_dst_addr[3]),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(channel_src_addr[60]),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(channel_dst_addr[90]),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(channel_src_addr[34]),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(src_rdata[31]),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(channel_dst_addr[7]),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(src_rdata[23]),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(src_rdata[30]),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(src_rdata[1]),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(channel_dst_addr[110]),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(src_rdata[4]),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(src_rdata[28]),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(src_rdata[0]),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(channel_src_addr[116]),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(channel_src_addr[10]),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(channel_src_addr[31]),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(src_rdata[51]),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(src_rdata[82]),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(channel_src_addr[58]),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(src_rdata[9]),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(channel_dst_addr[21]),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(src_rdata[18]),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(src_rdata[20]),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(channel_dst_addr[117]),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(channel_src_addr[14]),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(channel_src_addr[11]),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(src_rdata[16]),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(src_rdata[19]),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(src_rdata[3]),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(channel_dst_addr[91]),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(channel_dst_addr[61]),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(src_rdata[26]),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(channel_src_addr[115]),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(channel_src_addr[9]),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(channel_dst_addr[23]),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(channel_dst_addr[95]),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(src_rdata[54]),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(src_rdata[44]),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(channel_src_addr[47]),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(channel_src_addr[15]),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(src_rdata[22]),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(src_rdata[5]),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(channel_src_addr[3]),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(src_rdata[37]),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(src_rdata[21]),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(channel_src_addr[57]),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(channel_src_addr[20]),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(channel_src_addr[108]),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(channel_src_addr[12]),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(src_rdata[24]),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(channel_dst_addr[25]),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(channel_dst_addr[45]),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(channel_src_addr[100]),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(channel_dst_addr[118]),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(channel_src_addr[120]),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(src_rdata[17]),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(channel_src_addr[22]),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(channel_src_addr[40]),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(channel_dst_addr[27]),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(channel_dst_addr[26]),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(channel_dst_addr[20]),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(channel_dst_addr[119]),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(channel_dst_addr[38]),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(channel_dst_addr[34]),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(channel_src_addr[55]),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(channel_src_addr[6]),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(channel_dst_addr[29]),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(channel_dst_addr[121]),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(channel_dst_addr[53]),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(channel_dst_addr[9]),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(channel_src_addr[17]),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(channel_dst_addr[103]),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(channel_src_addr[110]),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(channel_src_addr[16]),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(channel_src_addr[0]),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(src_rdata[8]),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(channel_src_addr[99]),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(channel_src_addr[127]),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(channel_dst_addr[14]),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(channel_start[1]),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(channel_src_addr[104]),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(channel_start[0]),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(channel_dst_addr[94]),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(channel_src_addr[85]),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(channel_src_addr[2]),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(src_rdata[2]),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(channel_dst_addr[112]),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(channel_dst_addr[2]),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(channel_dst_addr[48]),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(channel_src_addr[21]),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(channel_dst_addr[62]),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(channel_src_addr[39]),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(src_rdata[6]),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(channel_src_addr[19]),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(channel_src_addr[38]),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(channel_dst_addr[55]),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(channel_dst_addr[30]),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(channel_dst_addr[5]),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(channel_src_addr[5]),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(channel_dst_addr[116]),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(channel_src_addr[50]),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(channel_dst_addr[57]),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(channel_dst_addr[28]),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(channel_dst_addr[120]),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(channel_dst_addr[24]),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(channel_src_addr[18]),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(channel_dst_addr[6]),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(channel_src_addr[76]),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(channel_dst_addr[12]),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(channel_dst_addr[36]),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(channel_src_addr[98]),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(channel_dst_addr[18]),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(channel_dst_addr[122]),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(channel_src_addr[71]),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(channel_src_addr[54]),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(channel_dst_addr[107]),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(channel_dst_addr[47]),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(channel_dst_addr[41]),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(channel_start[2]),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(channel_dst_addr[11]),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(channel_src_addr[13]),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(channel_src_addr[102]),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(channel_src_addr[114]),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(channel_src_addr[7]),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(channel_dst_addr[37]),
    .X(net1643));
endmodule
