module spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \debug_miso_samples[0] ;
 wire \debug_miso_samples[1] ;
 wire \debug_miso_samples[2] ;
 wire \debug_miso_samples[3] ;
 wire \debug_miso_samples[4] ;
 wire \debug_miso_samples[5] ;
 wire \debug_miso_samples[6] ;
 wire \debug_miso_samples[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \tx_shift[0] ;
 wire \tx_shift[1] ;
 wire \tx_shift[2] ;
 wire \tx_shift[3] ;
 wire \tx_shift[4] ;
 wire \tx_shift[5] ;
 wire \tx_shift[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 BUF_X4 _230_ (.A(\bit_count[2] ),
    .Z(_037_));
 INV_X1 _231_ (.A(\bit_count[3] ),
    .ZN(_038_));
 BUF_X4 _232_ (.A(_225_),
    .Z(_039_));
 NAND3_X4 _233_ (.A1(_037_),
    .A2(_038_),
    .A3(_039_),
    .ZN(_211_));
 INV_X1 _234_ (.A(_211_),
    .ZN(_216_));
 INV_X1 _235_ (.A(net1),
    .ZN(_040_));
 CLKBUF_X3 _236_ (.A(_040_),
    .Z(_041_));
 CLKBUF_X2 _237_ (.A(tx_valid),
    .Z(_042_));
 BUF_X4 _238_ (.A(\state[0] ),
    .Z(_043_));
 NAND2_X1 _239_ (.A1(_042_),
    .A2(_043_),
    .ZN(_044_));
 BUF_X4 _240_ (.A(\state[2] ),
    .Z(_045_));
 CLKBUF_X3 _241_ (.A(_045_),
    .Z(_046_));
 OAI21_X1 _242_ (.A(_046_),
    .B1(_211_),
    .B2(net20),
    .ZN(_047_));
 AOI21_X1 _243_ (.A(_041_),
    .B1(_044_),
    .B2(_047_),
    .ZN(_002_));
 INV_X1 _244_ (.A(_042_),
    .ZN(_048_));
 NAND2_X1 _245_ (.A1(_048_),
    .A2(_043_),
    .ZN(_049_));
 BUF_X4 _246_ (.A(\state[1] ),
    .Z(_050_));
 NOR2_X1 _247_ (.A1(_050_),
    .A2(_041_),
    .ZN(_051_));
 NAND2_X1 _248_ (.A1(_049_),
    .A2(_051_),
    .ZN(_001_));
 INV_X2 _249_ (.A(_045_),
    .ZN(_052_));
 NOR4_X1 _250_ (.A1(_041_),
    .A2(net20),
    .A3(_052_),
    .A4(_211_),
    .ZN(_000_));
 BUF_X1 _251_ (.A(\bit_count[0] ),
    .Z(_053_));
 NAND3_X1 _252_ (.A1(_037_),
    .A2(\bit_count[1] ),
    .A3(_053_),
    .ZN(_227_));
 OR2_X1 _253_ (.A1(\bit_count[3] ),
    .A2(_227_),
    .ZN(_219_));
 NAND3_X1 _254_ (.A1(_037_),
    .A2(_038_),
    .A3(_039_),
    .ZN(_222_));
 BUF_X2 _255_ (.A(net1),
    .Z(_054_));
 BUF_X2 _256_ (.A(_004_),
    .Z(_055_));
 NAND2_X1 _257_ (.A1(_045_),
    .A2(_055_),
    .ZN(_056_));
 AOI21_X2 _258_ (.A(_056_),
    .B1(_043_),
    .B2(_048_),
    .ZN(_057_));
 MUX2_X1 _259_ (.A(_043_),
    .B(_055_),
    .S(_045_),
    .Z(_058_));
 INV_X2 _260_ (.A(\state[0] ),
    .ZN(_059_));
 OAI21_X2 _261_ (.A(_058_),
    .B1(_059_),
    .B2(_042_),
    .ZN(_060_));
 MUX2_X1 _262_ (.A(_057_),
    .B(_060_),
    .S(_053_),
    .Z(_061_));
 AND2_X1 _263_ (.A1(_054_),
    .A2(_061_),
    .ZN(_005_));
 CLKBUF_X3 _264_ (.A(_041_),
    .Z(_062_));
 BUF_X2 _265_ (.A(_226_),
    .Z(_063_));
 AOI22_X1 _266_ (.A1(\bit_count[1] ),
    .A2(_060_),
    .B1(_057_),
    .B2(_063_),
    .ZN(_064_));
 NOR2_X1 _267_ (.A1(_062_),
    .A2(_064_),
    .ZN(_006_));
 AND2_X2 _268_ (.A1(_045_),
    .A2(_055_),
    .ZN(_065_));
 INV_X1 _269_ (.A(_039_),
    .ZN(_066_));
 AOI211_X4 _270_ (.A(_037_),
    .B(_066_),
    .C1(_048_),
    .C2(_043_),
    .ZN(_067_));
 AND2_X1 _271_ (.A1(_037_),
    .A2(_066_),
    .ZN(_068_));
 OAI21_X1 _272_ (.A(_065_),
    .B1(_067_),
    .B2(_068_),
    .ZN(_069_));
 NAND2_X1 _273_ (.A1(_037_),
    .A2(_060_),
    .ZN(_070_));
 AOI21_X1 _274_ (.A(_041_),
    .B1(_069_),
    .B2(_070_),
    .ZN(_007_));
 BUF_X2 _275_ (.A(_229_),
    .Z(_071_));
 AOI22_X1 _276_ (.A1(\bit_count[3] ),
    .A2(_060_),
    .B1(_057_),
    .B2(_071_),
    .ZN(_072_));
 NOR2_X1 _277_ (.A1(_062_),
    .A2(_072_),
    .ZN(_008_));
 AOI21_X4 _278_ (.A(_040_),
    .B1(_052_),
    .B2(_043_),
    .ZN(_073_));
 NAND2_X1 _279_ (.A1(_053_),
    .A2(_065_),
    .ZN(_074_));
 NAND3_X1 _280_ (.A1(\debug_miso_samples[0] ),
    .A2(_073_),
    .A3(_074_),
    .ZN(_075_));
 CLKBUF_X2 _281_ (.A(_213_),
    .Z(_076_));
 INV_X1 _282_ (.A(_076_),
    .ZN(_077_));
 INV_X1 _283_ (.A(_071_),
    .ZN(_078_));
 XOR2_X2 _284_ (.A(_037_),
    .B(_039_),
    .Z(_079_));
 NOR4_X2 _285_ (.A1(_077_),
    .A2(_063_),
    .A3(_078_),
    .A4(_079_),
    .ZN(_080_));
 NAND4_X4 _286_ (.A1(net1),
    .A2(_045_),
    .A3(_055_),
    .A4(net2),
    .ZN(_081_));
 NOR4_X2 _287_ (.A1(_217_),
    .A2(_214_),
    .A3(_003_),
    .A4(_081_),
    .ZN(_082_));
 INV_X1 _288_ (.A(_220_),
    .ZN(_083_));
 AND2_X1 _289_ (.A1(_076_),
    .A2(_221_),
    .ZN(_084_));
 NOR2_X1 _290_ (.A1(_223_),
    .A2(_228_),
    .ZN(_085_));
 AND4_X2 _291_ (.A1(_224_),
    .A2(_083_),
    .A3(_084_),
    .A4(_085_),
    .ZN(_086_));
 AND2_X1 _292_ (.A1(_220_),
    .A2(_223_),
    .ZN(_087_));
 NOR2_X2 _293_ (.A1(_221_),
    .A2(_224_),
    .ZN(_088_));
 AND4_X2 _294_ (.A1(_077_),
    .A2(_228_),
    .A3(_087_),
    .A4(_088_),
    .ZN(_089_));
 OAI211_X2 _295_ (.A(_080_),
    .B(_082_),
    .C1(_086_),
    .C2(_089_),
    .ZN(_090_));
 AND3_X1 _296_ (.A1(net1),
    .A2(_045_),
    .A3(_055_),
    .ZN(_091_));
 NAND2_X1 _297_ (.A1(\debug_miso_samples[0] ),
    .A2(_091_),
    .ZN(_092_));
 INV_X1 _298_ (.A(_063_),
    .ZN(_093_));
 XNOR2_X2 _299_ (.A(_037_),
    .B(_039_),
    .ZN(_094_));
 NAND4_X1 _300_ (.A1(_076_),
    .A2(_093_),
    .A3(_071_),
    .A4(_094_),
    .ZN(_095_));
 NOR2_X4 _301_ (.A1(_217_),
    .A2(_214_),
    .ZN(_096_));
 INV_X1 _302_ (.A(_096_),
    .ZN(_097_));
 NAND4_X1 _303_ (.A1(_224_),
    .A2(_083_),
    .A3(_084_),
    .A4(_085_),
    .ZN(_098_));
 NAND4_X4 _304_ (.A1(_077_),
    .A2(_228_),
    .A3(_087_),
    .A4(_088_),
    .ZN(_099_));
 AOI211_X2 _305_ (.A(_095_),
    .B(_097_),
    .C1(_098_),
    .C2(_099_),
    .ZN(_100_));
 OAI211_X2 _306_ (.A(_075_),
    .B(_090_),
    .C1(_092_),
    .C2(_100_),
    .ZN(_009_));
 INV_X1 _307_ (.A(\debug_miso_samples[1] ),
    .ZN(_101_));
 AOI21_X2 _308_ (.A(_065_),
    .B1(_052_),
    .B2(_043_),
    .ZN(_102_));
 NOR2_X1 _309_ (.A1(\bit_count[3] ),
    .A2(_053_),
    .ZN(_103_));
 NAND4_X1 _310_ (.A1(_063_),
    .A2(_078_),
    .A3(_079_),
    .A4(_103_),
    .ZN(_104_));
 AOI21_X1 _311_ (.A(_102_),
    .B1(_104_),
    .B2(_065_),
    .ZN(_105_));
 NOR2_X1 _312_ (.A1(_076_),
    .A2(_053_),
    .ZN(_106_));
 AND4_X1 _313_ (.A1(net2),
    .A2(_091_),
    .A3(_096_),
    .A4(_106_),
    .ZN(_107_));
 OAI21_X2 _314_ (.A(_107_),
    .B1(_089_),
    .B2(_086_),
    .ZN(_108_));
 NAND2_X1 _315_ (.A1(_063_),
    .A2(_078_),
    .ZN(_109_));
 OAI33_X1 _316_ (.A1(_041_),
    .A2(_101_),
    .A3(_105_),
    .B1(_108_),
    .B2(_094_),
    .B3(_109_),
    .ZN(_010_));
 NAND2_X1 _317_ (.A1(\debug_miso_samples[2] ),
    .A2(_073_),
    .ZN(_110_));
 NOR2_X1 _318_ (.A1(_076_),
    .A2(_003_),
    .ZN(_111_));
 NAND4_X1 _319_ (.A1(_063_),
    .A2(_078_),
    .A3(_096_),
    .A4(_111_),
    .ZN(_112_));
 NOR4_X1 _320_ (.A1(_102_),
    .A2(_099_),
    .A3(_094_),
    .A4(_112_),
    .ZN(_113_));
 OR2_X1 _321_ (.A1(_076_),
    .A2(_003_),
    .ZN(_114_));
 NOR4_X2 _322_ (.A1(_093_),
    .A2(_071_),
    .A3(_081_),
    .A4(_114_),
    .ZN(_115_));
 OAI211_X2 _323_ (.A(_096_),
    .B(_115_),
    .C1(_086_),
    .C2(_089_),
    .ZN(_116_));
 OAI22_X1 _324_ (.A1(_110_),
    .A2(_113_),
    .B1(_116_),
    .B2(_094_),
    .ZN(_011_));
 NOR2_X2 _325_ (.A1(_063_),
    .A2(_071_),
    .ZN(_117_));
 NAND2_X1 _326_ (.A1(_079_),
    .A2(_117_),
    .ZN(_118_));
 NAND2_X1 _327_ (.A1(_065_),
    .A2(_103_),
    .ZN(_119_));
 NOR2_X1 _328_ (.A1(_118_),
    .A2(_119_),
    .ZN(_120_));
 NAND2_X1 _329_ (.A1(\debug_miso_samples[3] ),
    .A2(_073_),
    .ZN(_121_));
 OAI22_X1 _330_ (.A1(_108_),
    .A2(_118_),
    .B1(_120_),
    .B2(_121_),
    .ZN(_012_));
 NAND2_X1 _331_ (.A1(_054_),
    .A2(\debug_miso_samples[4] ),
    .ZN(_122_));
 NOR2_X1 _332_ (.A1(_056_),
    .A2(_122_),
    .ZN(_123_));
 NAND4_X1 _333_ (.A1(_079_),
    .A2(_096_),
    .A3(_111_),
    .A4(_117_),
    .ZN(_124_));
 OAI21_X1 _334_ (.A(_123_),
    .B1(_124_),
    .B2(_099_),
    .ZN(_125_));
 OR2_X1 _335_ (.A1(_099_),
    .A2(_124_),
    .ZN(_126_));
 OAI221_X1 _336_ (.A(_125_),
    .B1(_126_),
    .B2(_081_),
    .C1(_058_),
    .C2(_122_),
    .ZN(_013_));
 NOR3_X1 _337_ (.A1(_079_),
    .A2(_109_),
    .A3(_119_),
    .ZN(_127_));
 INV_X1 _338_ (.A(_073_),
    .ZN(_128_));
 INV_X1 _339_ (.A(\debug_miso_samples[5] ),
    .ZN(_129_));
 OAI33_X1 _340_ (.A1(_079_),
    .A2(_109_),
    .A3(_108_),
    .B1(_127_),
    .B2(_128_),
    .B3(_129_),
    .ZN(_014_));
 NAND2_X1 _341_ (.A1(\debug_miso_samples[6] ),
    .A2(_073_),
    .ZN(_130_));
 NOR4_X1 _342_ (.A1(_102_),
    .A2(_099_),
    .A3(_079_),
    .A4(_112_),
    .ZN(_131_));
 OAI22_X1 _343_ (.A1(_079_),
    .A2(_116_),
    .B1(_130_),
    .B2(_131_),
    .ZN(_015_));
 NAND4_X1 _344_ (.A1(_058_),
    .A2(_094_),
    .A3(_103_),
    .A4(_117_),
    .ZN(_132_));
 NAND2_X1 _345_ (.A1(\debug_miso_samples[7] ),
    .A2(_132_),
    .ZN(_133_));
 AND4_X1 _346_ (.A1(net2),
    .A2(_094_),
    .A3(_106_),
    .A4(_117_),
    .ZN(_134_));
 OAI211_X2 _347_ (.A(_096_),
    .B(_134_),
    .C1(_086_),
    .C2(_089_),
    .ZN(_135_));
 OAI21_X1 _348_ (.A(\debug_miso_samples[7] ),
    .B1(_046_),
    .B2(_059_),
    .ZN(_136_));
 AOI221_X1 _349_ (.A(_041_),
    .B1(_133_),
    .B2(_135_),
    .C1(_136_),
    .C2(_056_),
    .ZN(_016_));
 MUX2_X1 _350_ (.A(net11),
    .B(\debug_miso_samples[0] ),
    .S(_050_),
    .Z(_137_));
 AND2_X1 _351_ (.A1(_054_),
    .A2(_137_),
    .ZN(_017_));
 MUX2_X1 _352_ (.A(net12),
    .B(\debug_miso_samples[1] ),
    .S(_050_),
    .Z(_138_));
 AND2_X1 _353_ (.A1(_054_),
    .A2(_138_),
    .ZN(_018_));
 MUX2_X1 _354_ (.A(net13),
    .B(\debug_miso_samples[2] ),
    .S(_050_),
    .Z(_139_));
 AND2_X1 _355_ (.A1(_054_),
    .A2(_139_),
    .ZN(_019_));
 MUX2_X1 _356_ (.A(net14),
    .B(\debug_miso_samples[3] ),
    .S(_050_),
    .Z(_140_));
 AND2_X1 _357_ (.A1(_054_),
    .A2(_140_),
    .ZN(_020_));
 MUX2_X1 _358_ (.A(net15),
    .B(\debug_miso_samples[4] ),
    .S(_050_),
    .Z(_141_));
 AND2_X1 _359_ (.A1(_054_),
    .A2(_141_),
    .ZN(_021_));
 MUX2_X1 _360_ (.A(net16),
    .B(\debug_miso_samples[5] ),
    .S(_050_),
    .Z(_142_));
 AND2_X1 _361_ (.A1(_054_),
    .A2(_142_),
    .ZN(_022_));
 MUX2_X1 _362_ (.A(net17),
    .B(\debug_miso_samples[6] ),
    .S(_050_),
    .Z(_143_));
 AND2_X1 _363_ (.A1(_054_),
    .A2(_143_),
    .ZN(_023_));
 MUX2_X1 _364_ (.A(net18),
    .B(\debug_miso_samples[7] ),
    .S(\state[1] ),
    .Z(_144_));
 AND2_X1 _365_ (.A1(_054_),
    .A2(_144_),
    .ZN(_024_));
 AOI21_X1 _366_ (.A(_050_),
    .B1(_059_),
    .B2(net19),
    .ZN(_145_));
 NOR2_X1 _367_ (.A1(_062_),
    .A2(_145_),
    .ZN(_025_));
 AOI21_X1 _368_ (.A(_065_),
    .B1(_052_),
    .B2(net20),
    .ZN(_146_));
 NOR4_X1 _369_ (.A1(_050_),
    .A2(_043_),
    .A3(_041_),
    .A4(_146_),
    .ZN(_026_));
 NAND2_X1 _370_ (.A1(_059_),
    .A2(net21),
    .ZN(_147_));
 NAND3_X1 _371_ (.A1(_049_),
    .A2(_051_),
    .A3(_147_),
    .ZN(_027_));
 OAI21_X1 _372_ (.A(net20),
    .B1(_055_),
    .B2(_212_),
    .ZN(_148_));
 NAND2_X2 _373_ (.A1(_046_),
    .A2(_148_),
    .ZN(_149_));
 MUX2_X2 _374_ (.A(_046_),
    .B(_042_),
    .S(_043_),
    .Z(_150_));
 AOI21_X1 _375_ (.A(net22),
    .B1(_149_),
    .B2(_150_),
    .ZN(_151_));
 AND2_X1 _376_ (.A1(_045_),
    .A2(_148_),
    .ZN(_152_));
 BUF_X2 _377_ (.A(_152_),
    .Z(_153_));
 MUX2_X2 _378_ (.A(_048_),
    .B(_052_),
    .S(_059_),
    .Z(_154_));
 MUX2_X1 _379_ (.A(net10),
    .B(\tx_shift[6] ),
    .S(_046_),
    .Z(_155_));
 NOR3_X1 _380_ (.A1(_153_),
    .A2(_154_),
    .A3(_155_),
    .ZN(_156_));
 NOR3_X1 _381_ (.A1(_062_),
    .A2(_151_),
    .A3(_156_),
    .ZN(_028_));
 AOI21_X1 _382_ (.A(_041_),
    .B1(net23),
    .B2(_059_),
    .ZN(_157_));
 NAND2_X1 _383_ (.A1(_049_),
    .A2(_157_),
    .ZN(_029_));
 OAI21_X1 _384_ (.A(\tx_shift[0] ),
    .B1(_153_),
    .B2(_154_),
    .ZN(_158_));
 NAND4_X1 _385_ (.A1(_042_),
    .A2(_043_),
    .A3(_052_),
    .A4(net3),
    .ZN(_159_));
 AOI21_X1 _386_ (.A(_041_),
    .B1(_158_),
    .B2(_159_),
    .ZN(_030_));
 AOI21_X1 _387_ (.A(\tx_shift[1] ),
    .B1(_149_),
    .B2(_150_),
    .ZN(_160_));
 MUX2_X1 _388_ (.A(net4),
    .B(\tx_shift[0] ),
    .S(_046_),
    .Z(_161_));
 NOR3_X1 _389_ (.A1(_153_),
    .A2(_154_),
    .A3(_161_),
    .ZN(_162_));
 NOR3_X1 _390_ (.A1(_062_),
    .A2(_160_),
    .A3(_162_),
    .ZN(_031_));
 AOI21_X1 _391_ (.A(\tx_shift[2] ),
    .B1(_149_),
    .B2(_150_),
    .ZN(_163_));
 MUX2_X1 _392_ (.A(net5),
    .B(\tx_shift[1] ),
    .S(_046_),
    .Z(_164_));
 NOR3_X1 _393_ (.A1(_153_),
    .A2(_154_),
    .A3(_164_),
    .ZN(_165_));
 NOR3_X1 _394_ (.A1(_062_),
    .A2(_163_),
    .A3(_165_),
    .ZN(_032_));
 AOI21_X1 _395_ (.A(\tx_shift[3] ),
    .B1(_149_),
    .B2(_150_),
    .ZN(_166_));
 MUX2_X1 _396_ (.A(net6),
    .B(\tx_shift[2] ),
    .S(_046_),
    .Z(_167_));
 NOR3_X1 _397_ (.A1(_153_),
    .A2(_154_),
    .A3(_167_),
    .ZN(_168_));
 NOR3_X1 _398_ (.A1(_062_),
    .A2(_166_),
    .A3(_168_),
    .ZN(_033_));
 AOI21_X1 _399_ (.A(\tx_shift[4] ),
    .B1(_149_),
    .B2(_150_),
    .ZN(_169_));
 MUX2_X1 _400_ (.A(net7),
    .B(\tx_shift[3] ),
    .S(_046_),
    .Z(_170_));
 NOR3_X1 _401_ (.A1(_153_),
    .A2(_154_),
    .A3(_170_),
    .ZN(_171_));
 NOR3_X1 _402_ (.A1(_062_),
    .A2(_169_),
    .A3(_171_),
    .ZN(_034_));
 AOI21_X1 _403_ (.A(\tx_shift[5] ),
    .B1(_149_),
    .B2(_150_),
    .ZN(_172_));
 MUX2_X1 _404_ (.A(net8),
    .B(\tx_shift[4] ),
    .S(_046_),
    .Z(_173_));
 NOR3_X1 _405_ (.A1(_153_),
    .A2(_154_),
    .A3(_173_),
    .ZN(_174_));
 NOR3_X1 _406_ (.A1(_062_),
    .A2(_172_),
    .A3(_174_),
    .ZN(_035_));
 AOI21_X1 _407_ (.A(\tx_shift[6] ),
    .B1(_149_),
    .B2(_150_),
    .ZN(_175_));
 MUX2_X1 _408_ (.A(net9),
    .B(\tx_shift[5] ),
    .S(_045_),
    .Z(_176_));
 NOR3_X1 _409_ (.A1(_153_),
    .A2(_154_),
    .A3(_176_),
    .ZN(_177_));
 NOR3_X1 _410_ (.A1(_062_),
    .A2(_175_),
    .A3(_177_),
    .ZN(_036_));
 HA_X1 _411_ (.A(_210_),
    .B(_211_),
    .CO(_212_),
    .S(_213_));
 HA_X1 _412_ (.A(\bit_count[3] ),
    .B(_211_),
    .CO(_214_),
    .S(_215_));
 HA_X1 _413_ (.A(\bit_count[3] ),
    .B(_216_),
    .CO(_217_),
    .S(_218_));
 HA_X1 _414_ (.A(_210_),
    .B(_219_),
    .CO(_220_),
    .S(_221_));
 HA_X1 _415_ (.A(_210_),
    .B(_222_),
    .CO(_223_),
    .S(_224_));
 HA_X1 _416_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_225_),
    .S(_226_));
 HA_X1 _417_ (.A(_210_),
    .B(_227_),
    .CO(_228_),
    .S(_229_));
 DFF_X1 \bit_count[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[0] ),
    .QN(_003_));
 DFF_X1 \bit_count[1]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_count[1] ),
    .QN(_206_));
 DFF_X1 \bit_count[2]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_count[2] ),
    .QN(_205_));
 DFF_X2 \bit_count[3]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_count[3] ),
    .QN(_210_));
 DFF_X1 \debug_miso_samples[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\debug_miso_samples[0] ),
    .QN(_204_));
 DFF_X1 \debug_miso_samples[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[1] ),
    .QN(_203_));
 DFF_X1 \debug_miso_samples[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[2] ),
    .QN(_202_));
 DFF_X1 \debug_miso_samples[3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[3] ),
    .QN(_201_));
 DFF_X1 \debug_miso_samples[4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[4] ),
    .QN(_200_));
 DFF_X1 \debug_miso_samples[5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[5] ),
    .QN(_199_));
 DFF_X1 \debug_miso_samples[6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\debug_miso_samples[6] ),
    .QN(_198_));
 DFF_X1 \debug_miso_samples[7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\debug_miso_samples[7] ),
    .QN(_197_));
 DFF_X1 \rx_data[0]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net11),
    .QN(_196_));
 DFF_X1 \rx_data[1]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net12),
    .QN(_195_));
 DFF_X1 \rx_data[2]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net13),
    .QN(_194_));
 DFF_X1 \rx_data[3]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net14),
    .QN(_193_));
 DFF_X1 \rx_data[4]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_192_));
 DFF_X1 \rx_data[5]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net16),
    .QN(_191_));
 DFF_X1 \rx_data[6]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_190_));
 DFF_X1 \rx_data[7]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net18),
    .QN(_189_));
 DFF_X1 \rx_valid$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net19),
    .QN(_188_));
 DFF_X2 \spi_clk$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net20),
    .QN(_004_));
 DFF_X1 \spi_cs_n$_SDFFE_PN1P_  (.D(_027_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net21),
    .QN(_187_));
 DFF_X1 \spi_mosi$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net22),
    .QN(_207_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[0] ),
    .QN(_208_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[1] ),
    .QN(_209_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[2] ),
    .QN(_186_));
 DFF_X1 \tx_ready$_SDFFE_PN1P_  (.D(_029_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net23),
    .QN(_185_));
 DFF_X1 \tx_shift[0]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[0] ),
    .QN(_184_));
 DFF_X1 \tx_shift[1]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[1] ),
    .QN(_183_));
 DFF_X1 \tx_shift[2]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[2] ),
    .QN(_182_));
 DFF_X1 \tx_shift[3]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[3] ),
    .QN(_181_));
 DFF_X1 \tx_shift[4]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[4] ),
    .QN(_180_));
 DFF_X1 \tx_shift[5]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[5] ),
    .QN(_179_));
 DFF_X1 \tx_shift[6]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[6] ),
    .QN(_178_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_55 ();
 CLKBUF_X2 input1 (.A(rst_n),
    .Z(net1));
 CLKBUF_X2 input2 (.A(spi_miso),
    .Z(net2));
 BUF_X1 input3 (.A(tx_data[0]),
    .Z(net3));
 BUF_X1 input4 (.A(tx_data[1]),
    .Z(net4));
 BUF_X1 input5 (.A(tx_data[2]),
    .Z(net5));
 BUF_X1 input6 (.A(tx_data[3]),
    .Z(net6));
 BUF_X1 input7 (.A(tx_data[4]),
    .Z(net7));
 BUF_X1 input8 (.A(tx_data[5]),
    .Z(net8));
 BUF_X1 input9 (.A(tx_data[6]),
    .Z(net9));
 BUF_X1 input10 (.A(tx_data[7]),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(rx_data[0]));
 BUF_X1 output12 (.A(net12),
    .Z(rx_data[1]));
 BUF_X1 output13 (.A(net13),
    .Z(rx_data[2]));
 BUF_X1 output14 (.A(net14),
    .Z(rx_data[3]));
 BUF_X1 output15 (.A(net15),
    .Z(rx_data[4]));
 BUF_X1 output16 (.A(net16),
    .Z(rx_data[5]));
 BUF_X1 output17 (.A(net17),
    .Z(rx_data[6]));
 BUF_X1 output18 (.A(net18),
    .Z(rx_data[7]));
 BUF_X1 output19 (.A(net19),
    .Z(rx_valid));
 BUF_X1 output20 (.A(net20),
    .Z(spi_clk));
 BUF_X1 output21 (.A(net21),
    .Z(spi_cs_n));
 BUF_X1 output22 (.A(net22),
    .Z(spi_mosi));
 BUF_X1 output23 (.A(net23),
    .Z(tx_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X1 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_2__leaf_clk));
 INV_X1 clkload2 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X2 FILLER_0_33 ();
 FILLCELL_X1 FILLER_0_35 ();
 FILLCELL_X32 FILLER_0_39 ();
 FILLCELL_X8 FILLER_0_71 ();
 FILLCELL_X1 FILLER_0_79 ();
 FILLCELL_X8 FILLER_0_83 ();
 FILLCELL_X4 FILLER_0_91 ();
 FILLCELL_X2 FILLER_0_95 ();
 FILLCELL_X4 FILLER_0_100 ();
 FILLCELL_X2 FILLER_0_104 ();
 FILLCELL_X1 FILLER_0_106 ();
 FILLCELL_X2 FILLER_0_110 ();
 FILLCELL_X16 FILLER_0_116 ();
 FILLCELL_X1 FILLER_0_132 ();
 FILLCELL_X8 FILLER_0_136 ();
 FILLCELL_X2 FILLER_0_144 ();
 FILLCELL_X8 FILLER_0_149 ();
 FILLCELL_X4 FILLER_0_157 ();
 FILLCELL_X2 FILLER_0_161 ();
 FILLCELL_X2 FILLER_0_169 ();
 FILLCELL_X32 FILLER_0_174 ();
 FILLCELL_X2 FILLER_0_206 ();
 FILLCELL_X1 FILLER_0_208 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X4 FILLER_1_33 ();
 FILLCELL_X2 FILLER_1_37 ();
 FILLCELL_X1 FILLER_1_39 ();
 FILLCELL_X4 FILLER_1_60 ();
 FILLCELL_X2 FILLER_1_64 ();
 FILLCELL_X1 FILLER_1_66 ();
 FILLCELL_X2 FILLER_1_84 ();
 FILLCELL_X8 FILLER_1_89 ();
 FILLCELL_X4 FILLER_1_97 ();
 FILLCELL_X2 FILLER_1_101 ();
 FILLCELL_X1 FILLER_1_103 ();
 FILLCELL_X4 FILLER_1_111 ();
 FILLCELL_X2 FILLER_1_115 ();
 FILLCELL_X4 FILLER_1_141 ();
 FILLCELL_X2 FILLER_1_145 ();
 FILLCELL_X1 FILLER_1_147 ();
 FILLCELL_X2 FILLER_1_165 ();
 FILLCELL_X2 FILLER_1_174 ();
 FILLCELL_X1 FILLER_1_176 ();
 FILLCELL_X1 FILLER_1_181 ();
 FILLCELL_X4 FILLER_1_203 ();
 FILLCELL_X2 FILLER_1_207 ();
 FILLCELL_X16 FILLER_2_1 ();
 FILLCELL_X2 FILLER_2_17 ();
 FILLCELL_X4 FILLER_2_43 ();
 FILLCELL_X16 FILLER_2_54 ();
 FILLCELL_X4 FILLER_2_70 ();
 FILLCELL_X2 FILLER_2_74 ();
 FILLCELL_X4 FILLER_2_83 ();
 FILLCELL_X1 FILLER_2_87 ();
 FILLCELL_X1 FILLER_2_105 ();
 FILLCELL_X2 FILLER_2_110 ();
 FILLCELL_X2 FILLER_2_116 ();
 FILLCELL_X4 FILLER_2_122 ();
 FILLCELL_X2 FILLER_2_126 ();
 FILLCELL_X1 FILLER_2_128 ();
 FILLCELL_X8 FILLER_2_133 ();
 FILLCELL_X4 FILLER_2_141 ();
 FILLCELL_X2 FILLER_2_145 ();
 FILLCELL_X4 FILLER_2_155 ();
 FILLCELL_X8 FILLER_2_163 ();
 FILLCELL_X1 FILLER_2_171 ();
 FILLCELL_X2 FILLER_2_179 ();
 FILLCELL_X1 FILLER_2_181 ();
 FILLCELL_X16 FILLER_2_186 ();
 FILLCELL_X4 FILLER_2_202 ();
 FILLCELL_X2 FILLER_2_206 ();
 FILLCELL_X1 FILLER_2_208 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X2 FILLER_3_49 ();
 FILLCELL_X32 FILLER_3_54 ();
 FILLCELL_X8 FILLER_3_86 ();
 FILLCELL_X2 FILLER_3_94 ();
 FILLCELL_X1 FILLER_3_96 ();
 FILLCELL_X2 FILLER_3_101 ();
 FILLCELL_X32 FILLER_3_108 ();
 FILLCELL_X32 FILLER_3_140 ();
 FILLCELL_X32 FILLER_3_172 ();
 FILLCELL_X4 FILLER_3_204 ();
 FILLCELL_X1 FILLER_3_208 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_33 ();
 FILLCELL_X8 FILLER_4_44 ();
 FILLCELL_X2 FILLER_4_52 ();
 FILLCELL_X32 FILLER_4_57 ();
 FILLCELL_X8 FILLER_4_89 ();
 FILLCELL_X16 FILLER_4_120 ();
 FILLCELL_X8 FILLER_4_136 ();
 FILLCELL_X4 FILLER_4_144 ();
 FILLCELL_X1 FILLER_4_148 ();
 FILLCELL_X4 FILLER_4_173 ();
 FILLCELL_X1 FILLER_4_177 ();
 FILLCELL_X16 FILLER_4_182 ();
 FILLCELL_X8 FILLER_4_198 ();
 FILLCELL_X2 FILLER_4_206 ();
 FILLCELL_X1 FILLER_4_208 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X1 FILLER_5_50 ();
 FILLCELL_X4 FILLER_5_61 ();
 FILLCELL_X2 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_67 ();
 FILLCELL_X8 FILLER_5_87 ();
 FILLCELL_X4 FILLER_5_95 ();
 FILLCELL_X2 FILLER_5_99 ();
 FILLCELL_X32 FILLER_5_103 ();
 FILLCELL_X8 FILLER_5_135 ();
 FILLCELL_X4 FILLER_5_143 ();
 FILLCELL_X2 FILLER_5_147 ();
 FILLCELL_X8 FILLER_5_168 ();
 FILLCELL_X4 FILLER_5_176 ();
 FILLCELL_X2 FILLER_5_188 ();
 FILLCELL_X2 FILLER_5_207 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X4 FILLER_6_73 ();
 FILLCELL_X4 FILLER_6_86 ();
 FILLCELL_X1 FILLER_6_90 ();
 FILLCELL_X16 FILLER_6_95 ();
 FILLCELL_X8 FILLER_6_111 ();
 FILLCELL_X1 FILLER_6_119 ();
 FILLCELL_X16 FILLER_6_124 ();
 FILLCELL_X8 FILLER_6_140 ();
 FILLCELL_X4 FILLER_6_148 ();
 FILLCELL_X2 FILLER_6_152 ();
 FILLCELL_X16 FILLER_6_158 ();
 FILLCELL_X4 FILLER_6_174 ();
 FILLCELL_X2 FILLER_6_178 ();
 FILLCELL_X1 FILLER_6_180 ();
 FILLCELL_X16 FILLER_6_185 ();
 FILLCELL_X8 FILLER_6_201 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_61 ();
 FILLCELL_X8 FILLER_7_93 ();
 FILLCELL_X1 FILLER_7_101 ();
 FILLCELL_X8 FILLER_7_107 ();
 FILLCELL_X4 FILLER_7_122 ();
 FILLCELL_X1 FILLER_7_126 ();
 FILLCELL_X16 FILLER_7_132 ();
 FILLCELL_X8 FILLER_7_148 ();
 FILLCELL_X4 FILLER_7_160 ();
 FILLCELL_X1 FILLER_7_164 ();
 FILLCELL_X4 FILLER_7_169 ();
 FILLCELL_X2 FILLER_7_173 ();
 FILLCELL_X1 FILLER_7_186 ();
 FILLCELL_X16 FILLER_7_190 ();
 FILLCELL_X2 FILLER_7_206 ();
 FILLCELL_X1 FILLER_7_208 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_33 ();
 FILLCELL_X1 FILLER_8_41 ();
 FILLCELL_X4 FILLER_8_49 ();
 FILLCELL_X16 FILLER_8_68 ();
 FILLCELL_X2 FILLER_8_84 ();
 FILLCELL_X1 FILLER_8_86 ();
 FILLCELL_X8 FILLER_8_94 ();
 FILLCELL_X2 FILLER_8_109 ();
 FILLCELL_X1 FILLER_8_111 ();
 FILLCELL_X8 FILLER_8_115 ();
 FILLCELL_X4 FILLER_8_152 ();
 FILLCELL_X8 FILLER_8_173 ();
 FILLCELL_X1 FILLER_8_181 ();
 FILLCELL_X4 FILLER_8_186 ();
 FILLCELL_X1 FILLER_8_190 ();
 FILLCELL_X8 FILLER_8_194 ();
 FILLCELL_X4 FILLER_8_202 ();
 FILLCELL_X2 FILLER_8_206 ();
 FILLCELL_X1 FILLER_8_208 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X2 FILLER_9_57 ();
 FILLCELL_X1 FILLER_9_59 ();
 FILLCELL_X8 FILLER_9_64 ();
 FILLCELL_X1 FILLER_9_72 ();
 FILLCELL_X8 FILLER_9_83 ();
 FILLCELL_X4 FILLER_9_106 ();
 FILLCELL_X2 FILLER_9_110 ();
 FILLCELL_X1 FILLER_9_112 ();
 FILLCELL_X32 FILLER_9_117 ();
 FILLCELL_X16 FILLER_9_149 ();
 FILLCELL_X8 FILLER_9_165 ();
 FILLCELL_X2 FILLER_9_173 ();
 FILLCELL_X16 FILLER_9_192 ();
 FILLCELL_X1 FILLER_9_208 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_17 ();
 FILLCELL_X1 FILLER_10_25 ();
 FILLCELL_X8 FILLER_10_45 ();
 FILLCELL_X2 FILLER_10_53 ();
 FILLCELL_X1 FILLER_10_55 ();
 FILLCELL_X16 FILLER_10_58 ();
 FILLCELL_X1 FILLER_10_74 ();
 FILLCELL_X8 FILLER_10_79 ();
 FILLCELL_X4 FILLER_10_87 ();
 FILLCELL_X2 FILLER_10_91 ();
 FILLCELL_X1 FILLER_10_93 ();
 FILLCELL_X32 FILLER_10_99 ();
 FILLCELL_X8 FILLER_10_131 ();
 FILLCELL_X4 FILLER_10_139 ();
 FILLCELL_X2 FILLER_10_143 ();
 FILLCELL_X1 FILLER_10_145 ();
 FILLCELL_X32 FILLER_10_151 ();
 FILLCELL_X16 FILLER_10_183 ();
 FILLCELL_X8 FILLER_10_199 ();
 FILLCELL_X2 FILLER_10_207 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_33 ();
 FILLCELL_X2 FILLER_11_40 ();
 FILLCELL_X1 FILLER_11_42 ();
 FILLCELL_X8 FILLER_11_46 ();
 FILLCELL_X2 FILLER_11_54 ();
 FILLCELL_X2 FILLER_11_69 ();
 FILLCELL_X1 FILLER_11_73 ();
 FILLCELL_X8 FILLER_11_84 ();
 FILLCELL_X4 FILLER_11_92 ();
 FILLCELL_X16 FILLER_11_101 ();
 FILLCELL_X4 FILLER_11_117 ();
 FILLCELL_X1 FILLER_11_121 ();
 FILLCELL_X2 FILLER_11_126 ();
 FILLCELL_X1 FILLER_11_128 ();
 FILLCELL_X8 FILLER_11_146 ();
 FILLCELL_X2 FILLER_11_154 ();
 FILLCELL_X1 FILLER_11_156 ();
 FILLCELL_X2 FILLER_11_164 ();
 FILLCELL_X1 FILLER_11_166 ();
 FILLCELL_X2 FILLER_11_195 ();
 FILLCELL_X8 FILLER_11_200 ();
 FILLCELL_X1 FILLER_11_208 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_43 ();
 FILLCELL_X4 FILLER_12_51 ();
 FILLCELL_X2 FILLER_12_55 ();
 FILLCELL_X1 FILLER_12_59 ();
 FILLCELL_X2 FILLER_12_67 ();
 FILLCELL_X1 FILLER_12_69 ();
 FILLCELL_X8 FILLER_12_80 ();
 FILLCELL_X1 FILLER_12_88 ();
 FILLCELL_X2 FILLER_12_92 ();
 FILLCELL_X1 FILLER_12_94 ();
 FILLCELL_X2 FILLER_12_97 ();
 FILLCELL_X1 FILLER_12_99 ();
 FILLCELL_X2 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_148 ();
 FILLCELL_X16 FILLER_12_180 ();
 FILLCELL_X8 FILLER_12_196 ();
 FILLCELL_X4 FILLER_12_204 ();
 FILLCELL_X1 FILLER_12_208 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_17 ();
 FILLCELL_X2 FILLER_13_21 ();
 FILLCELL_X2 FILLER_13_27 ();
 FILLCELL_X1 FILLER_13_29 ();
 FILLCELL_X8 FILLER_13_46 ();
 FILLCELL_X1 FILLER_13_54 ();
 FILLCELL_X16 FILLER_13_59 ();
 FILLCELL_X4 FILLER_13_75 ();
 FILLCELL_X1 FILLER_13_88 ();
 FILLCELL_X32 FILLER_13_112 ();
 FILLCELL_X32 FILLER_13_144 ();
 FILLCELL_X32 FILLER_13_176 ();
 FILLCELL_X1 FILLER_13_208 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X8 FILLER_14_17 ();
 FILLCELL_X4 FILLER_14_25 ();
 FILLCELL_X1 FILLER_14_32 ();
 FILLCELL_X8 FILLER_14_50 ();
 FILLCELL_X8 FILLER_14_68 ();
 FILLCELL_X2 FILLER_14_76 ();
 FILLCELL_X16 FILLER_14_87 ();
 FILLCELL_X8 FILLER_14_103 ();
 FILLCELL_X1 FILLER_14_111 ();
 FILLCELL_X16 FILLER_14_117 ();
 FILLCELL_X32 FILLER_14_136 ();
 FILLCELL_X32 FILLER_14_168 ();
 FILLCELL_X8 FILLER_14_200 ();
 FILLCELL_X1 FILLER_14_208 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_25 ();
 FILLCELL_X1 FILLER_15_40 ();
 FILLCELL_X8 FILLER_15_48 ();
 FILLCELL_X4 FILLER_15_56 ();
 FILLCELL_X2 FILLER_15_60 ();
 FILLCELL_X4 FILLER_15_71 ();
 FILLCELL_X2 FILLER_15_75 ();
 FILLCELL_X1 FILLER_15_77 ();
 FILLCELL_X16 FILLER_15_85 ();
 FILLCELL_X4 FILLER_15_101 ();
 FILLCELL_X2 FILLER_15_105 ();
 FILLCELL_X4 FILLER_15_112 ();
 FILLCELL_X1 FILLER_15_116 ();
 FILLCELL_X4 FILLER_15_122 ();
 FILLCELL_X2 FILLER_15_126 ();
 FILLCELL_X2 FILLER_15_142 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X2 FILLER_15_162 ();
 FILLCELL_X4 FILLER_15_167 ();
 FILLCELL_X8 FILLER_15_182 ();
 FILLCELL_X2 FILLER_15_207 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X8 FILLER_16_17 ();
 FILLCELL_X1 FILLER_16_25 ();
 FILLCELL_X4 FILLER_16_30 ();
 FILLCELL_X2 FILLER_16_34 ();
 FILLCELL_X32 FILLER_16_40 ();
 FILLCELL_X2 FILLER_16_72 ();
 FILLCELL_X1 FILLER_16_74 ();
 FILLCELL_X4 FILLER_16_78 ();
 FILLCELL_X1 FILLER_16_82 ();
 FILLCELL_X32 FILLER_16_99 ();
 FILLCELL_X32 FILLER_16_131 ();
 FILLCELL_X32 FILLER_16_163 ();
 FILLCELL_X8 FILLER_16_195 ();
 FILLCELL_X2 FILLER_16_203 ();
 FILLCELL_X1 FILLER_16_205 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_33 ();
 FILLCELL_X1 FILLER_17_37 ();
 FILLCELL_X16 FILLER_17_42 ();
 FILLCELL_X8 FILLER_17_58 ();
 FILLCELL_X2 FILLER_17_66 ();
 FILLCELL_X1 FILLER_17_68 ();
 FILLCELL_X2 FILLER_17_72 ();
 FILLCELL_X8 FILLER_17_82 ();
 FILLCELL_X16 FILLER_17_102 ();
 FILLCELL_X32 FILLER_17_121 ();
 FILLCELL_X16 FILLER_17_153 ();
 FILLCELL_X8 FILLER_17_169 ();
 FILLCELL_X4 FILLER_17_177 ();
 FILLCELL_X16 FILLER_17_185 ();
 FILLCELL_X8 FILLER_17_201 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_33 ();
 FILLCELL_X1 FILLER_18_35 ();
 FILLCELL_X1 FILLER_18_46 ();
 FILLCELL_X1 FILLER_18_51 ();
 FILLCELL_X1 FILLER_18_72 ();
 FILLCELL_X8 FILLER_18_82 ();
 FILLCELL_X2 FILLER_18_90 ();
 FILLCELL_X2 FILLER_18_94 ();
 FILLCELL_X2 FILLER_18_105 ();
 FILLCELL_X1 FILLER_18_112 ();
 FILLCELL_X16 FILLER_18_151 ();
 FILLCELL_X8 FILLER_18_167 ();
 FILLCELL_X1 FILLER_18_199 ();
 FILLCELL_X4 FILLER_18_203 ();
 FILLCELL_X2 FILLER_18_207 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_33 ();
 FILLCELL_X2 FILLER_19_37 ();
 FILLCELL_X2 FILLER_19_58 ();
 FILLCELL_X4 FILLER_19_67 ();
 FILLCELL_X2 FILLER_19_71 ();
 FILLCELL_X1 FILLER_19_73 ();
 FILLCELL_X2 FILLER_19_83 ();
 FILLCELL_X1 FILLER_19_85 ();
 FILLCELL_X32 FILLER_19_102 ();
 FILLCELL_X4 FILLER_19_134 ();
 FILLCELL_X1 FILLER_19_138 ();
 FILLCELL_X4 FILLER_19_142 ();
 FILLCELL_X32 FILLER_19_153 ();
 FILLCELL_X16 FILLER_19_185 ();
 FILLCELL_X8 FILLER_19_201 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_33 ();
 FILLCELL_X2 FILLER_20_41 ();
 FILLCELL_X1 FILLER_20_43 ();
 FILLCELL_X16 FILLER_20_58 ();
 FILLCELL_X8 FILLER_20_74 ();
 FILLCELL_X16 FILLER_20_84 ();
 FILLCELL_X4 FILLER_20_100 ();
 FILLCELL_X16 FILLER_20_112 ();
 FILLCELL_X8 FILLER_20_128 ();
 FILLCELL_X1 FILLER_20_136 ();
 FILLCELL_X2 FILLER_20_141 ();
 FILLCELL_X32 FILLER_20_151 ();
 FILLCELL_X16 FILLER_20_183 ();
 FILLCELL_X8 FILLER_20_199 ();
 FILLCELL_X2 FILLER_20_207 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X16 FILLER_21_33 ();
 FILLCELL_X4 FILLER_21_49 ();
 FILLCELL_X4 FILLER_21_70 ();
 FILLCELL_X2 FILLER_21_74 ();
 FILLCELL_X16 FILLER_21_85 ();
 FILLCELL_X8 FILLER_21_101 ();
 FILLCELL_X1 FILLER_21_114 ();
 FILLCELL_X8 FILLER_21_120 ();
 FILLCELL_X4 FILLER_21_128 ();
 FILLCELL_X2 FILLER_21_132 ();
 FILLCELL_X1 FILLER_21_134 ();
 FILLCELL_X1 FILLER_21_137 ();
 FILLCELL_X1 FILLER_21_148 ();
 FILLCELL_X8 FILLER_21_151 ();
 FILLCELL_X4 FILLER_21_176 ();
 FILLCELL_X2 FILLER_21_180 ();
 FILLCELL_X16 FILLER_21_186 ();
 FILLCELL_X4 FILLER_21_202 ();
 FILLCELL_X2 FILLER_21_206 ();
 FILLCELL_X1 FILLER_21_208 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_65 ();
 FILLCELL_X2 FILLER_22_77 ();
 FILLCELL_X1 FILLER_22_79 ();
 FILLCELL_X16 FILLER_22_83 ();
 FILLCELL_X4 FILLER_22_99 ();
 FILLCELL_X4 FILLER_22_111 ();
 FILLCELL_X2 FILLER_22_115 ();
 FILLCELL_X8 FILLER_22_122 ();
 FILLCELL_X2 FILLER_22_130 ();
 FILLCELL_X1 FILLER_22_135 ();
 FILLCELL_X16 FILLER_22_153 ();
 FILLCELL_X4 FILLER_22_169 ();
 FILLCELL_X2 FILLER_22_173 ();
 FILLCELL_X1 FILLER_22_175 ();
 FILLCELL_X4 FILLER_22_200 ();
 FILLCELL_X2 FILLER_22_207 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_82 ();
 FILLCELL_X8 FILLER_23_115 ();
 FILLCELL_X1 FILLER_23_123 ();
 FILLCELL_X32 FILLER_23_141 ();
 FILLCELL_X32 FILLER_23_173 ();
 FILLCELL_X4 FILLER_23_205 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X16 FILLER_24_129 ();
 FILLCELL_X4 FILLER_24_145 ();
 FILLCELL_X2 FILLER_24_149 ();
 FILLCELL_X1 FILLER_24_151 ();
 FILLCELL_X32 FILLER_24_159 ();
 FILLCELL_X16 FILLER_24_191 ();
 FILLCELL_X2 FILLER_24_207 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_33 ();
 FILLCELL_X4 FILLER_25_41 ();
 FILLCELL_X2 FILLER_25_45 ();
 FILLCELL_X4 FILLER_25_51 ();
 FILLCELL_X8 FILLER_25_62 ();
 FILLCELL_X32 FILLER_25_87 ();
 FILLCELL_X32 FILLER_25_119 ();
 FILLCELL_X4 FILLER_25_151 ();
 FILLCELL_X2 FILLER_25_155 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_193 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X8 FILLER_26_33 ();
 FILLCELL_X1 FILLER_26_41 ();
 FILLCELL_X16 FILLER_26_59 ();
 FILLCELL_X8 FILLER_26_75 ();
 FILLCELL_X1 FILLER_26_83 ();
 FILLCELL_X1 FILLER_26_101 ();
 FILLCELL_X4 FILLER_26_113 ();
 FILLCELL_X2 FILLER_26_134 ();
 FILLCELL_X4 FILLER_26_147 ();
 FILLCELL_X2 FILLER_26_151 ();
 FILLCELL_X32 FILLER_26_170 ();
 FILLCELL_X4 FILLER_26_202 ();
 FILLCELL_X2 FILLER_26_206 ();
 FILLCELL_X1 FILLER_26_208 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X16 FILLER_27_33 ();
 FILLCELL_X4 FILLER_27_49 ();
 FILLCELL_X2 FILLER_27_53 ();
 FILLCELL_X1 FILLER_27_55 ();
 FILLCELL_X32 FILLER_27_59 ();
 FILLCELL_X2 FILLER_27_91 ();
 FILLCELL_X32 FILLER_27_96 ();
 FILLCELL_X8 FILLER_27_128 ();
 FILLCELL_X16 FILLER_27_139 ();
 FILLCELL_X8 FILLER_27_155 ();
 FILLCELL_X2 FILLER_27_163 ();
 FILLCELL_X32 FILLER_27_168 ();
 FILLCELL_X8 FILLER_27_200 ();
 FILLCELL_X1 FILLER_27_208 ();
endmodule
