module ahb_lite_master (hbusreq,
    hclk,
    hgrant,
    hready,
    hreset,
    hwrite,
    start_trans,
    trans_done,
    trans_write,
    haddr,
    hburst,
    hrdata,
    hresp,
    hsize,
    htrans,
    hwdata,
    read_data,
    trans_addr,
    trans_burst,
    trans_resp,
    trans_size,
    write_data);
 output hbusreq;
 input hclk;
 input hgrant;
 input hready;
 input hreset;
 output hwrite;
 input start_trans;
 output trans_done;
 input trans_write;
 output [31:0] haddr;
 output [2:0] hburst;
 input [31:0] hrdata;
 input [1:0] hresp;
 output [2:0] hsize;
 output [1:0] htrans;
 output [31:0] hwdata;
 output [31:0] read_data;
 input [31:0] trans_addr;
 input [2:0] trans_burst;
 output [1:0] trans_resp;
 input [2:0] trans_size;
 input [31:0] write_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire \burst_count[0] ;
 wire \burst_count[1] ;
 wire \burst_count[2] ;
 wire \burst_count[3] ;
 wire \burst_count[4] ;
 wire \burst_count[5] ;
 wire \burst_count[6] ;
 wire \burst_count[7] ;
 wire \burst_total[0] ;
 wire \burst_total[2] ;
 wire \burst_total[3] ;
 wire \burst_total[4] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;

 sky130_fd_sc_hd__nor3_1 _482_ (.A(\burst_total[3] ),
    .B(\burst_total[2] ),
    .C(\burst_total[0] ),
    .Y(_440_));
 sky130_fd_sc_hd__inv_1 _483_ (.A(\burst_total[4] ),
    .Y(_439_));
 sky130_fd_sc_hd__xnor2_1 _484_ (.A(\burst_total[3] ),
    .B(_450_),
    .Y(_445_));
 sky130_fd_sc_hd__or3b_1 _485_ (.A(net148),
    .B(net149),
    .C_N(net147),
    .X(_426_));
 sky130_fd_sc_hd__inv_1 _486_ (.A(_426_),
    .Y(_459_));
 sky130_fd_sc_hd__nor3b_1 _487_ (.A(net147),
    .B(net149),
    .C_N(net148),
    .Y(_462_));
 sky130_fd_sc_hd__and3b_1 _488_ (.A_N(net149),
    .B(net147),
    .C(net148),
    .X(_465_));
 sky130_fd_sc_hd__nor3b_1 _489_ (.A(net148),
    .B(net147),
    .C_N(net149),
    .Y(_468_));
 sky130_fd_sc_hd__nand2_1 _490_ (.A(net147),
    .B(net149),
    .Y(_121_));
 sky130_fd_sc_hd__nor2_1 _491_ (.A(net148),
    .B(_121_),
    .Y(_471_));
 sky130_fd_sc_hd__and3b_1 _492_ (.A_N(net147),
    .B(net149),
    .C(net148),
    .X(_474_));
 sky130_fd_sc_hd__and3_1 _493_ (.A(net148),
    .B(net147),
    .C(net149),
    .X(_477_));
 sky130_fd_sc_hd__buf_6 _494_ (.A(\state[2] ),
    .X(_122_));
 sky130_fd_sc_hd__clkbuf_4 _495_ (.A(\state[1] ),
    .X(_123_));
 sky130_fd_sc_hd__nand2b_1 _496_ (.A_N(net35),
    .B(\state[1] ),
    .Y(_124_));
 sky130_fd_sc_hd__buf_6 _497_ (.A(\state[0] ),
    .X(_125_));
 sky130_fd_sc_hd__o211ai_1 _498_ (.A1(_123_),
    .A2(net2),
    .B1(_124_),
    .C1(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2b_1 _499_ (.A(_123_),
    .B_N(net39),
    .Y(_127_));
 sky130_fd_sc_hd__a211o_1 _500_ (.A1(_123_),
    .A2(net35),
    .B1(_127_),
    .C1(_125_),
    .X(_128_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(_126_),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nand4b_4 _502_ (.A_N(_122_),
    .B(_125_),
    .C(_123_),
    .D(net35),
    .Y(_130_));
 sky130_fd_sc_hd__nand2_1 _503_ (.A(_432_),
    .B(_435_),
    .Y(_131_));
 sky130_fd_sc_hd__nand2_1 _504_ (.A(_438_),
    .B(_444_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2_1 _505_ (.A(_131_),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__inv_1 _506_ (.A(_446_),
    .Y(_134_));
 sky130_fd_sc_hd__o21ai_0 _507_ (.A1(_453_),
    .A2(_452_),
    .B1(_447_),
    .Y(_135_));
 sky130_fd_sc_hd__o21ai_0 _508_ (.A1(\burst_total[0] ),
    .A2(\burst_count[0] ),
    .B1(_455_),
    .Y(_136_));
 sky130_fd_sc_hd__nor3_1 _509_ (.A(_446_),
    .B(_452_),
    .C(_454_),
    .Y(_137_));
 sky130_fd_sc_hd__a22oi_2 _510_ (.A1(_134_),
    .A2(_135_),
    .B1(_136_),
    .B2(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__a21oi_1 _511_ (.A1(_443_),
    .A2(_438_),
    .B1(_437_),
    .Y(_139_));
 sky130_fd_sc_hd__a21oi_1 _512_ (.A1(_432_),
    .A2(_434_),
    .B1(_431_),
    .Y(_140_));
 sky130_fd_sc_hd__o21ai_2 _513_ (.A1(_131_),
    .A2(_139_),
    .B1(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__a21oi_1 _514_ (.A1(_133_),
    .A2(_138_),
    .B1(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__nor3_2 _515_ (.A(_441_),
    .B(_130_),
    .C(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__o21bai_1 _516_ (.A1(_122_),
    .A2(_129_),
    .B1_N(_143_),
    .Y(_422_));
 sky130_fd_sc_hd__xnor2_1 _517_ (.A(_122_),
    .B(_123_),
    .Y(_144_));
 sky130_fd_sc_hd__nand3b_1 _518_ (.A_N(_123_),
    .B(net2),
    .C(_125_),
    .Y(_145_));
 sky130_fd_sc_hd__a21o_1 _519_ (.A1(_124_),
    .A2(_145_),
    .B1(_122_),
    .X(_146_));
 sky130_fd_sc_hd__o21ai_0 _520_ (.A1(_125_),
    .A2(_144_),
    .B1(_146_),
    .Y(_423_));
 sky130_fd_sc_hd__inv_1 _521_ (.A(_130_),
    .Y(_424_));
 sky130_fd_sc_hd__inv_1 _522_ (.A(net122),
    .Y(_425_));
 sky130_fd_sc_hd__inv_1 _523_ (.A(_457_),
    .Y(_427_));
 sky130_fd_sc_hd__inv_1 _524_ (.A(\burst_total[0] ),
    .Y(_448_));
 sky130_fd_sc_hd__nor2_1 _525_ (.A(\burst_total[3] ),
    .B(\burst_total[4] ),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _526_ (.A(_450_),
    .B(_147_),
    .Y(_430_));
 sky130_fd_sc_hd__nand2_1 _527_ (.A(_439_),
    .B(_440_),
    .Y(_433_));
 sky130_fd_sc_hd__nand2_1 _528_ (.A(_439_),
    .B(_440_),
    .Y(_436_));
 sky130_fd_sc_hd__inv_1 _529_ (.A(\burst_total[2] ),
    .Y(_449_));
 sky130_fd_sc_hd__nor3_1 _530_ (.A(net148),
    .B(net147),
    .C(net149),
    .Y(_456_));
 sky130_fd_sc_hd__nor2_1 _531_ (.A(_441_),
    .B(_142_),
    .Y(_148_));
 sky130_fd_sc_hd__nor3b_4 _532_ (.A(_122_),
    .B(_125_),
    .C_N(\state[1] ),
    .Y(_149_));
 sky130_fd_sc_hd__nand2_1 _533_ (.A(net35),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__a211oi_2 _534_ (.A1(_133_),
    .A2(_138_),
    .B1(_141_),
    .C1(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__nor2_2 _535_ (.A(_122_),
    .B(_125_),
    .Y(_152_));
 sky130_fd_sc_hd__nand2_2 _536_ (.A(_127_),
    .B(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__nand3_1 _537_ (.A(net35),
    .B(_441_),
    .C(_149_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _538_ (.A(_153_),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__nor2_2 _539_ (.A(_151_),
    .B(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _540_ (.A(\burst_count[0] ),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__o31ai_1 _541_ (.A1(\burst_count[0] ),
    .A2(_148_),
    .A3(_150_),
    .B1(_157_),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _542_ (.A(_481_),
    .B(_149_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2_1 _543_ (.A(\burst_count[1] ),
    .B(_156_),
    .Y(_159_));
 sky130_fd_sc_hd__o21ai_0 _544_ (.A1(_156_),
    .A2(_158_),
    .B1(_159_),
    .Y(_001_));
 sky130_fd_sc_hd__and2_0 _545_ (.A(_127_),
    .B(_152_),
    .X(_160_));
 sky130_fd_sc_hd__buf_4 _546_ (.A(_160_),
    .X(_161_));
 sky130_fd_sc_hd__o21ai_0 _547_ (.A1(_151_),
    .A2(_155_),
    .B1(_480_),
    .Y(_162_));
 sky130_fd_sc_hd__xor2_1 _548_ (.A(\burst_count[2] ),
    .B(_162_),
    .X(_163_));
 sky130_fd_sc_hd__nor2_1 _549_ (.A(_161_),
    .B(_163_),
    .Y(_002_));
 sky130_fd_sc_hd__o2111ai_1 _550_ (.A1(_151_),
    .A2(_155_),
    .B1(\burst_count[2] ),
    .C1(\burst_count[0] ),
    .D1(\burst_count[1] ),
    .Y(_164_));
 sky130_fd_sc_hd__xor2_1 _551_ (.A(\burst_count[3] ),
    .B(_164_),
    .X(_165_));
 sky130_fd_sc_hd__nor2_1 _552_ (.A(_161_),
    .B(_165_),
    .Y(_003_));
 sky130_fd_sc_hd__nand3_1 _553_ (.A(\burst_count[2] ),
    .B(_480_),
    .C(\burst_count[3] ),
    .Y(_166_));
 sky130_fd_sc_hd__o21ai_0 _554_ (.A1(_156_),
    .A2(_166_),
    .B1(\burst_count[4] ),
    .Y(_167_));
 sky130_fd_sc_hd__or3_1 _555_ (.A(\burst_count[4] ),
    .B(_156_),
    .C(_166_),
    .X(_168_));
 sky130_fd_sc_hd__a21oi_1 _556_ (.A1(_167_),
    .A2(_168_),
    .B1(_161_),
    .Y(_004_));
 sky130_fd_sc_hd__and4_1 _557_ (.A(\burst_count[4] ),
    .B(\burst_count[2] ),
    .C(\burst_count[0] ),
    .D(\burst_count[1] ),
    .X(_169_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(\burst_count[3] ),
    .B(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__o21ai_0 _559_ (.A1(_156_),
    .A2(_170_),
    .B1(\burst_count[5] ),
    .Y(_171_));
 sky130_fd_sc_hd__or3_1 _560_ (.A(\burst_count[5] ),
    .B(_156_),
    .C(_170_),
    .X(_172_));
 sky130_fd_sc_hd__a21oi_1 _561_ (.A1(_171_),
    .A2(_172_),
    .B1(_161_),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _562_ (.A(\burst_count[6] ),
    .B(_153_),
    .Y(_173_));
 sky130_fd_sc_hd__nand2b_1 _563_ (.A_N(\burst_count[6] ),
    .B(_153_),
    .Y(_174_));
 sky130_fd_sc_hd__o211ai_1 _564_ (.A1(_151_),
    .A2(_155_),
    .B1(\burst_count[5] ),
    .C1(\burst_count[3] ),
    .Y(_175_));
 sky130_fd_sc_hd__nand3_1 _565_ (.A(\burst_count[4] ),
    .B(\burst_count[2] ),
    .C(_480_),
    .Y(_176_));
 sky130_fd_sc_hd__nor2_1 _566_ (.A(_175_),
    .B(_176_),
    .Y(_177_));
 sky130_fd_sc_hd__mux2i_1 _567_ (.A0(_173_),
    .A1(_174_),
    .S(_177_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _568_ (.A(\burst_count[6] ),
    .B(_169_),
    .Y(_178_));
 sky130_fd_sc_hd__o21ai_0 _569_ (.A1(_175_),
    .A2(_178_),
    .B1(\burst_count[7] ),
    .Y(_179_));
 sky130_fd_sc_hd__or3_1 _570_ (.A(\burst_count[7] ),
    .B(_175_),
    .C(_178_),
    .X(_180_));
 sky130_fd_sc_hd__a21oi_1 _571_ (.A1(_179_),
    .A2(_180_),
    .B1(_161_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_1 _572_ (.A(net72),
    .B(net73),
    .Y(_181_));
 sky130_fd_sc_hd__nand3b_1 _573_ (.A_N(net74),
    .B(_161_),
    .C(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__o21ai_0 _574_ (.A1(_448_),
    .A2(_161_),
    .B1(_182_),
    .Y(_008_));
 sky130_fd_sc_hd__or3_1 _575_ (.A(net74),
    .B(_153_),
    .C(_181_),
    .X(_183_));
 sky130_fd_sc_hd__o21ai_0 _576_ (.A1(_449_),
    .A2(_161_),
    .B1(_183_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _577_ (.A(\burst_total[3] ),
    .B(_153_),
    .Y(_184_));
 sky130_fd_sc_hd__nand3b_1 _578_ (.A_N(net73),
    .B(_161_),
    .C(net74),
    .Y(_185_));
 sky130_fd_sc_hd__nand2_1 _579_ (.A(_184_),
    .B(_185_),
    .Y(_010_));
 sky130_fd_sc_hd__nand3_1 _580_ (.A(net74),
    .B(net73),
    .C(_160_),
    .Y(_186_));
 sky130_fd_sc_hd__o21ai_0 _581_ (.A1(_439_),
    .A2(_161_),
    .B1(_186_),
    .Y(_011_));
 sky130_fd_sc_hd__nor3b_2 _582_ (.A(_122_),
    .B(\state[1] ),
    .C_N(_125_),
    .Y(_187_));
 sky130_fd_sc_hd__o21a_1 _583_ (.A1(\state[1] ),
    .A2(net2),
    .B1(_187_),
    .X(_188_));
 sky130_fd_sc_hd__clkbuf_4 _584_ (.A(_188_),
    .X(_189_));
 sky130_fd_sc_hd__mux2_1 _585_ (.A0(net143),
    .A1(net72),
    .S(_189_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _586_ (.A0(net144),
    .A1(net73),
    .S(_189_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _587_ (.A0(net145),
    .A1(net74),
    .S(_189_),
    .X(_014_));
 sky130_fd_sc_hd__nand2_2 _588_ (.A(_123_),
    .B(_152_),
    .Y(_190_));
 sky130_fd_sc_hd__buf_4 _589_ (.A(_190_),
    .X(_191_));
 sky130_fd_sc_hd__a21oi_1 _590_ (.A1(net39),
    .A2(_191_),
    .B1(_187_),
    .Y(_192_));
 sky130_fd_sc_hd__inv_1 _591_ (.A(net146),
    .Y(_193_));
 sky130_fd_sc_hd__or3_1 _592_ (.A(net145),
    .B(net144),
    .C(net143),
    .X(_194_));
 sky130_fd_sc_hd__nand2_1 _593_ (.A(_149_),
    .B(_194_),
    .Y(_195_));
 sky130_fd_sc_hd__nand2b_1 _594_ (.A_N(_125_),
    .B(net35),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_1 _595_ (.A1(_123_),
    .A2(_196_),
    .B1(_122_),
    .Y(_197_));
 sky130_fd_sc_hd__o21ai_2 _596_ (.A1(_148_),
    .A2(_195_),
    .B1(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__mux2i_1 _597_ (.A0(_192_),
    .A1(_193_),
    .S(_198_),
    .Y(_015_));
 sky130_fd_sc_hd__mux2_1 _598_ (.A0(net147),
    .A1(net75),
    .S(_189_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _599_ (.A0(net148),
    .A1(net76),
    .S(_189_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _600_ (.A0(net149),
    .A1(net77),
    .S(_189_),
    .X(_018_));
 sky130_fd_sc_hd__nor2_1 _601_ (.A(_122_),
    .B(\state[1] ),
    .Y(_199_));
 sky130_fd_sc_hd__a22o_1 _602_ (.A1(_124_),
    .A2(_152_),
    .B1(_199_),
    .B2(net2),
    .X(_200_));
 sky130_fd_sc_hd__nor2b_1 _603_ (.A(net2),
    .B_N(_187_),
    .Y(_201_));
 sky130_fd_sc_hd__o22a_1 _604_ (.A1(net150),
    .A2(_200_),
    .B1(_198_),
    .B2(_201_),
    .X(_019_));
 sky130_fd_sc_hd__o22a_1 _605_ (.A1(net151),
    .A2(_200_),
    .B1(_198_),
    .B2(_187_),
    .X(_020_));
 sky130_fd_sc_hd__nand3_4 _606_ (.A(net35),
    .B(net184),
    .C(_149_),
    .Y(_202_));
 sky130_fd_sc_hd__clkbuf_4 _607_ (.A(_202_),
    .X(_203_));
 sky130_fd_sc_hd__mux2_1 _608_ (.A0(net79),
    .A1(net152),
    .S(_203_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _609_ (.A0(net80),
    .A1(net153),
    .S(_203_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _610_ (.A0(net81),
    .A1(net154),
    .S(_203_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _611_ (.A0(net82),
    .A1(net155),
    .S(_203_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _612_ (.A0(net83),
    .A1(net156),
    .S(_203_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _613_ (.A0(net84),
    .A1(net157),
    .S(_203_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _614_ (.A0(net85),
    .A1(net158),
    .S(_203_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _615_ (.A0(net86),
    .A1(net159),
    .S(_203_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _616_ (.A0(net87),
    .A1(net160),
    .S(_203_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _617_ (.A0(net88),
    .A1(net161),
    .S(_203_),
    .X(_030_));
 sky130_fd_sc_hd__buf_4 _618_ (.A(_202_),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _619_ (.A0(net89),
    .A1(net162),
    .S(_204_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _620_ (.A0(net90),
    .A1(net163),
    .S(_204_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _621_ (.A0(net91),
    .A1(net164),
    .S(_204_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _622_ (.A0(net92),
    .A1(net165),
    .S(_204_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _623_ (.A0(net93),
    .A1(net166),
    .S(_204_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _624_ (.A0(net94),
    .A1(net167),
    .S(_204_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _625_ (.A0(net95),
    .A1(net168),
    .S(_204_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _626_ (.A0(net96),
    .A1(net169),
    .S(_204_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _627_ (.A0(net97),
    .A1(net170),
    .S(_204_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _628_ (.A0(net98),
    .A1(net171),
    .S(_204_),
    .X(_040_));
 sky130_fd_sc_hd__clkbuf_4 _629_ (.A(_202_),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _630_ (.A0(net99),
    .A1(net172),
    .S(_205_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _631_ (.A0(net100),
    .A1(net173),
    .S(_205_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _632_ (.A0(net101),
    .A1(net174),
    .S(_205_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _633_ (.A0(net102),
    .A1(net175),
    .S(_205_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _634_ (.A0(net103),
    .A1(net176),
    .S(_205_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _635_ (.A0(net104),
    .A1(net177),
    .S(_205_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _636_ (.A0(net105),
    .A1(net178),
    .S(_205_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _637_ (.A0(net106),
    .A1(net179),
    .S(_205_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _638_ (.A0(net107),
    .A1(net180),
    .S(_205_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _639_ (.A0(net108),
    .A1(net181),
    .S(_205_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _640_ (.A0(net109),
    .A1(net182),
    .S(_202_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _641_ (.A0(net110),
    .A1(net183),
    .S(_202_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _642_ (.A0(net184),
    .A1(net78),
    .S(_189_),
    .X(_053_));
 sky130_fd_sc_hd__nand4_1 _643_ (.A(_123_),
    .B(net35),
    .C(_152_),
    .D(_194_),
    .Y(_206_));
 sky130_fd_sc_hd__a211oi_2 _644_ (.A1(_133_),
    .A2(_138_),
    .B1(_141_),
    .C1(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__a41o_1 _645_ (.A1(_441_),
    .A2(_149_),
    .A3(_200_),
    .A4(_194_),
    .B1(_189_),
    .X(_208_));
 sky130_fd_sc_hd__or2_0 _646_ (.A(_207_),
    .B(_208_),
    .X(_209_));
 sky130_fd_sc_hd__buf_6 _647_ (.A(_209_),
    .X(_210_));
 sky130_fd_sc_hd__buf_6 _648_ (.A(_210_),
    .X(_211_));
 sky130_fd_sc_hd__nor2_1 _649_ (.A(net111),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__clkbuf_4 _650_ (.A(_190_),
    .X(_213_));
 sky130_fd_sc_hd__nor2_1 _651_ (.A(net145),
    .B(net144),
    .Y(_214_));
 sky130_fd_sc_hd__nor2_1 _652_ (.A(net143),
    .B(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__nor2_1 _653_ (.A(_190_),
    .B(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__clkbuf_4 _654_ (.A(_216_),
    .X(_217_));
 sky130_fd_sc_hd__nor2_4 _655_ (.A(_207_),
    .B(_208_),
    .Y(_218_));
 sky130_fd_sc_hd__clkbuf_4 _656_ (.A(_218_),
    .X(_219_));
 sky130_fd_sc_hd__a221oi_1 _657_ (.A1(net40),
    .A2(_213_),
    .B1(_217_),
    .B2(_458_),
    .C1(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__nor2_1 _658_ (.A(_212_),
    .B(_220_),
    .Y(_054_));
 sky130_fd_sc_hd__buf_2 _659_ (.A(_218_),
    .X(_221_));
 sky130_fd_sc_hd__nand2b_1 _660_ (.A_N(_428_),
    .B(_464_),
    .Y(_222_));
 sky130_fd_sc_hd__nor2_1 _661_ (.A(_463_),
    .B(_466_),
    .Y(_223_));
 sky130_fd_sc_hd__o211ai_1 _662_ (.A1(_467_),
    .A2(_466_),
    .B1(_473_),
    .C1(_470_),
    .Y(_224_));
 sky130_fd_sc_hd__a21o_1 _663_ (.A1(_222_),
    .A2(_223_),
    .B1(_224_),
    .X(_225_));
 sky130_fd_sc_hd__clkbuf_2 _664_ (.A(_479_),
    .X(_226_));
 sky130_fd_sc_hd__a21oi_1 _665_ (.A1(_226_),
    .A2(_475_),
    .B1(_478_),
    .Y(_227_));
 sky130_fd_sc_hd__a21oi_1 _666_ (.A1(_473_),
    .A2(_469_),
    .B1(_472_),
    .Y(_228_));
 sky130_fd_sc_hd__and2_0 _667_ (.A(_227_),
    .B(_228_),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_2 _668_ (.A(_476_),
    .X(_230_));
 sky130_fd_sc_hd__o21a_1 _669_ (.A1(_230_),
    .A2(_475_),
    .B1(_226_),
    .X(_231_));
 sky130_fd_sc_hd__and2_0 _670_ (.A(net141),
    .B(net142),
    .X(_232_));
 sky130_fd_sc_hd__buf_4 _671_ (.A(_232_),
    .X(_233_));
 sky130_fd_sc_hd__o21ai_1 _672_ (.A1(_478_),
    .A2(_231_),
    .B1(_233_),
    .Y(_234_));
 sky130_fd_sc_hd__a21oi_2 _673_ (.A1(_225_),
    .A2(_229_),
    .B1(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__o21ai_2 _674_ (.A1(net143),
    .A2(_214_),
    .B1(_149_),
    .Y(_236_));
 sky130_fd_sc_hd__clkbuf_4 _675_ (.A(_236_),
    .X(_237_));
 sky130_fd_sc_hd__nor2_1 _676_ (.A(net112),
    .B(_237_),
    .Y(_238_));
 sky130_fd_sc_hd__a22oi_1 _677_ (.A1(net41),
    .A2(_213_),
    .B1(_235_),
    .B2(_238_),
    .Y(_239_));
 sky130_fd_sc_hd__buf_2 _678_ (.A(_236_),
    .X(_240_));
 sky130_fd_sc_hd__nor2_1 _679_ (.A(_240_),
    .B(_235_),
    .Y(_241_));
 sky130_fd_sc_hd__o21ai_0 _680_ (.A1(_221_),
    .A2(_241_),
    .B1(net112),
    .Y(_242_));
 sky130_fd_sc_hd__o21ai_0 _681_ (.A1(_221_),
    .A2(_239_),
    .B1(_242_),
    .Y(_055_));
 sky130_fd_sc_hd__clkbuf_4 _682_ (.A(_236_),
    .X(_243_));
 sky130_fd_sc_hd__o211ai_1 _683_ (.A1(_464_),
    .A2(_463_),
    .B1(_470_),
    .C1(_467_),
    .Y(_244_));
 sky130_fd_sc_hd__a211oi_1 _684_ (.A1(_457_),
    .A2(_461_),
    .B1(_460_),
    .C1(_463_),
    .Y(_245_));
 sky130_fd_sc_hd__a21oi_1 _685_ (.A1(_470_),
    .A2(_466_),
    .B1(_469_),
    .Y(_246_));
 sky130_fd_sc_hd__o21ai_2 _686_ (.A1(_244_),
    .A2(_245_),
    .B1(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__nand3_1 _687_ (.A(_230_),
    .B(_226_),
    .C(_472_),
    .Y(_248_));
 sky130_fd_sc_hd__nand2_1 _688_ (.A(_227_),
    .B(_248_),
    .Y(_249_));
 sky130_fd_sc_hd__a41oi_2 _689_ (.A1(_473_),
    .A2(_230_),
    .A3(_226_),
    .A4(_247_),
    .B1(_249_),
    .Y(_250_));
 sky130_fd_sc_hd__clkbuf_4 _690_ (.A(_250_),
    .X(_251_));
 sky130_fd_sc_hd__nand2_1 _691_ (.A(net112),
    .B(_233_),
    .Y(_252_));
 sky130_fd_sc_hd__nor4_1 _692_ (.A(net113),
    .B(_243_),
    .C(_251_),
    .D(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__a21oi_1 _693_ (.A1(net42),
    .A2(_191_),
    .B1(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__a41o_2 _694_ (.A1(_473_),
    .A2(_230_),
    .A3(_226_),
    .A4(_247_),
    .B1(_249_),
    .X(_255_));
 sky130_fd_sc_hd__buf_2 _695_ (.A(_236_),
    .X(_256_));
 sky130_fd_sc_hd__a31oi_1 _696_ (.A1(net112),
    .A2(_233_),
    .A3(_255_),
    .B1(_256_),
    .Y(_257_));
 sky130_fd_sc_hd__o21ai_0 _697_ (.A1(_219_),
    .A2(_257_),
    .B1(net113),
    .Y(_258_));
 sky130_fd_sc_hd__o21ai_0 _698_ (.A1(_221_),
    .A2(_254_),
    .B1(_258_),
    .Y(_056_));
 sky130_fd_sc_hd__inv_1 _699_ (.A(net114),
    .Y(_259_));
 sky130_fd_sc_hd__nand2_1 _700_ (.A(_230_),
    .B(_226_),
    .Y(_260_));
 sky130_fd_sc_hd__a21o_1 _701_ (.A1(_225_),
    .A2(_228_),
    .B1(_260_),
    .X(_261_));
 sky130_fd_sc_hd__nand2_1 _702_ (.A(net112),
    .B(net113),
    .Y(_262_));
 sky130_fd_sc_hd__nand2_2 _703_ (.A(net141),
    .B(net142),
    .Y(_263_));
 sky130_fd_sc_hd__a211o_1 _704_ (.A1(_227_),
    .A2(_261_),
    .B1(_262_),
    .C1(_263_),
    .X(_264_));
 sky130_fd_sc_hd__a21oi_1 _705_ (.A1(_217_),
    .A2(_264_),
    .B1(_218_),
    .Y(_265_));
 sky130_fd_sc_hd__clkbuf_4 _706_ (.A(_190_),
    .X(_266_));
 sky130_fd_sc_hd__nand2_1 _707_ (.A(net43),
    .B(_266_),
    .Y(_267_));
 sky130_fd_sc_hd__o31a_1 _708_ (.A1(net114),
    .A2(_243_),
    .A3(_264_),
    .B1(_267_),
    .X(_268_));
 sky130_fd_sc_hd__clkbuf_4 _709_ (.A(_218_),
    .X(_269_));
 sky130_fd_sc_hd__o22ai_1 _710_ (.A1(_259_),
    .A2(_265_),
    .B1(_268_),
    .B2(_269_),
    .Y(_057_));
 sky130_fd_sc_hd__buf_2 _711_ (.A(_209_),
    .X(_270_));
 sky130_fd_sc_hd__and3_1 _712_ (.A(net112),
    .B(net113),
    .C(net114),
    .X(_271_));
 sky130_fd_sc_hd__nand2_2 _713_ (.A(_233_),
    .B(_271_),
    .Y(_272_));
 sky130_fd_sc_hd__nand2_1 _714_ (.A(net44),
    .B(_266_),
    .Y(_273_));
 sky130_fd_sc_hd__o41ai_1 _715_ (.A1(net115),
    .A2(_236_),
    .A3(_251_),
    .A4(_272_),
    .B1(_273_),
    .Y(_274_));
 sky130_fd_sc_hd__o21ai_0 _716_ (.A1(_251_),
    .A2(_272_),
    .B1(_217_),
    .Y(_275_));
 sky130_fd_sc_hd__nand2_1 _717_ (.A(_210_),
    .B(_275_),
    .Y(_276_));
 sky130_fd_sc_hd__a22o_1 _718_ (.A1(_270_),
    .A2(_274_),
    .B1(_276_),
    .B2(net115),
    .X(_058_));
 sky130_fd_sc_hd__nand2_1 _719_ (.A(net115),
    .B(_271_),
    .Y(_277_));
 sky130_fd_sc_hd__nor3_1 _720_ (.A(net116),
    .B(_243_),
    .C(_277_),
    .Y(_278_));
 sky130_fd_sc_hd__a22oi_1 _721_ (.A1(net45),
    .A2(_213_),
    .B1(_235_),
    .B2(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__a31oi_1 _722_ (.A1(net115),
    .A2(_235_),
    .A3(_271_),
    .B1(_256_),
    .Y(_280_));
 sky130_fd_sc_hd__o21ai_0 _723_ (.A1(_219_),
    .A2(_280_),
    .B1(net116),
    .Y(_281_));
 sky130_fd_sc_hd__o21ai_0 _724_ (.A1(_221_),
    .A2(_279_),
    .B1(_281_),
    .Y(_059_));
 sky130_fd_sc_hd__nand2_1 _725_ (.A(net116),
    .B(_233_),
    .Y(_282_));
 sky130_fd_sc_hd__nor2_1 _726_ (.A(_277_),
    .B(_282_),
    .Y(_283_));
 sky130_fd_sc_hd__nor4b_1 _727_ (.A(net117),
    .B(_243_),
    .C(_251_),
    .D_N(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__a21oi_1 _728_ (.A1(net46),
    .A2(_191_),
    .B1(_284_),
    .Y(_285_));
 sky130_fd_sc_hd__a21oi_1 _729_ (.A1(_255_),
    .A2(_283_),
    .B1(_240_),
    .Y(_286_));
 sky130_fd_sc_hd__o21ai_0 _730_ (.A1(_219_),
    .A2(_286_),
    .B1(net117),
    .Y(_287_));
 sky130_fd_sc_hd__o21ai_0 _731_ (.A1(_221_),
    .A2(_285_),
    .B1(_287_),
    .Y(_060_));
 sky130_fd_sc_hd__and2_0 _732_ (.A(_225_),
    .B(_229_),
    .X(_288_));
 sky130_fd_sc_hd__buf_2 _733_ (.A(_288_),
    .X(_289_));
 sky130_fd_sc_hd__nand3_1 _734_ (.A(net112),
    .B(net113),
    .C(net114),
    .Y(_290_));
 sky130_fd_sc_hd__nand3_2 _735_ (.A(net115),
    .B(net116),
    .C(net117),
    .Y(_291_));
 sky130_fd_sc_hd__nor2_1 _736_ (.A(_290_),
    .B(_291_),
    .Y(_292_));
 sky130_fd_sc_hd__nand2b_1 _737_ (.A_N(_234_),
    .B(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__buf_2 _738_ (.A(_293_),
    .X(_294_));
 sky130_fd_sc_hd__or3_1 _739_ (.A(_236_),
    .B(_289_),
    .C(_294_),
    .X(_295_));
 sky130_fd_sc_hd__nand2_1 _740_ (.A(net47),
    .B(_266_),
    .Y(_296_));
 sky130_fd_sc_hd__o21ai_0 _741_ (.A1(net118),
    .A2(_295_),
    .B1(_296_),
    .Y(_297_));
 sky130_fd_sc_hd__o21ai_0 _742_ (.A1(_289_),
    .A2(_294_),
    .B1(_216_),
    .Y(_298_));
 sky130_fd_sc_hd__a21boi_0 _743_ (.A1(_210_),
    .A2(_298_),
    .B1_N(net118),
    .Y(_299_));
 sky130_fd_sc_hd__a21o_1 _744_ (.A1(_211_),
    .A2(_297_),
    .B1(_299_),
    .X(_061_));
 sky130_fd_sc_hd__nor3_1 _745_ (.A(_251_),
    .B(_272_),
    .C(_291_),
    .Y(_300_));
 sky130_fd_sc_hd__nor3b_1 _746_ (.A(net119),
    .B(_243_),
    .C_N(net118),
    .Y(_301_));
 sky130_fd_sc_hd__a22oi_1 _747_ (.A1(net48),
    .A2(_213_),
    .B1(_300_),
    .B2(_301_),
    .Y(_302_));
 sky130_fd_sc_hd__a41oi_1 _748_ (.A1(net118),
    .A2(_233_),
    .A3(_255_),
    .A4(_292_),
    .B1(_256_),
    .Y(_303_));
 sky130_fd_sc_hd__o21ai_0 _749_ (.A1(_219_),
    .A2(_303_),
    .B1(net119),
    .Y(_304_));
 sky130_fd_sc_hd__o21ai_0 _750_ (.A1(_221_),
    .A2(_302_),
    .B1(_304_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2_1 _751_ (.A(net118),
    .B(net119),
    .Y(_305_));
 sky130_fd_sc_hd__nand2_1 _752_ (.A(net49),
    .B(_266_),
    .Y(_306_));
 sky130_fd_sc_hd__o31ai_1 _753_ (.A1(net120),
    .A2(_295_),
    .A3(_305_),
    .B1(_306_),
    .Y(_307_));
 sky130_fd_sc_hd__nor3_1 _754_ (.A(_289_),
    .B(_294_),
    .C(_305_),
    .Y(_308_));
 sky130_fd_sc_hd__o21ai_0 _755_ (.A1(_256_),
    .A2(_308_),
    .B1(_210_),
    .Y(_309_));
 sky130_fd_sc_hd__a22o_1 _756_ (.A1(_270_),
    .A2(_307_),
    .B1(_309_),
    .B2(net120),
    .X(_063_));
 sky130_fd_sc_hd__or2_1 _757_ (.A(_290_),
    .B(_291_),
    .X(_310_));
 sky130_fd_sc_hd__nand3_1 _758_ (.A(net118),
    .B(net119),
    .C(net120),
    .Y(_311_));
 sky130_fd_sc_hd__nor4_1 _759_ (.A(_263_),
    .B(_251_),
    .C(_310_),
    .D(_311_),
    .Y(_312_));
 sky130_fd_sc_hd__o21ai_0 _760_ (.A1(_240_),
    .A2(_312_),
    .B1(_270_),
    .Y(_313_));
 sky130_fd_sc_hd__nor2_1 _761_ (.A(net121),
    .B(_256_),
    .Y(_314_));
 sky130_fd_sc_hd__a22oi_1 _762_ (.A1(net50),
    .A2(_191_),
    .B1(_312_),
    .B2(_314_),
    .Y(_315_));
 sky130_fd_sc_hd__o2bb2ai_1 _763_ (.A1_N(net121),
    .A2_N(_313_),
    .B1(_315_),
    .B2(_269_),
    .Y(_064_));
 sky130_fd_sc_hd__a221oi_1 _764_ (.A1(net51),
    .A2(_266_),
    .B1(_217_),
    .B2(_429_),
    .C1(_218_),
    .Y(_316_));
 sky130_fd_sc_hd__a21oi_1 _765_ (.A1(_425_),
    .A2(_269_),
    .B1(_316_),
    .Y(_065_));
 sky130_fd_sc_hd__nand4_2 _766_ (.A(net118),
    .B(net119),
    .C(net120),
    .D(net121),
    .Y(_317_));
 sky130_fd_sc_hd__nor3_1 _767_ (.A(_289_),
    .B(_294_),
    .C(_317_),
    .Y(_318_));
 sky130_fd_sc_hd__o21ai_0 _768_ (.A1(_237_),
    .A2(_318_),
    .B1(_210_),
    .Y(_319_));
 sky130_fd_sc_hd__inv_1 _769_ (.A(net123),
    .Y(_320_));
 sky130_fd_sc_hd__a32o_1 _770_ (.A1(_320_),
    .A2(_216_),
    .A3(_318_),
    .B1(net52),
    .B2(_266_),
    .X(_321_));
 sky130_fd_sc_hd__a22o_1 _771_ (.A1(net123),
    .A2(_319_),
    .B1(_321_),
    .B2(_211_),
    .X(_066_));
 sky130_fd_sc_hd__nor3_1 _772_ (.A(_243_),
    .B(_251_),
    .C(_272_),
    .Y(_322_));
 sky130_fd_sc_hd__nor2_1 _773_ (.A(_320_),
    .B(_317_),
    .Y(_323_));
 sky130_fd_sc_hd__nor2_1 _774_ (.A(net124),
    .B(_291_),
    .Y(_324_));
 sky130_fd_sc_hd__a32oi_1 _775_ (.A1(_322_),
    .A2(_323_),
    .A3(_324_),
    .B1(_191_),
    .B2(net53),
    .Y(_325_));
 sky130_fd_sc_hd__a41oi_1 _776_ (.A1(_233_),
    .A2(_255_),
    .A3(_292_),
    .A4(_323_),
    .B1(_256_),
    .Y(_326_));
 sky130_fd_sc_hd__o21ai_0 _777_ (.A1(_219_),
    .A2(_326_),
    .B1(net124),
    .Y(_327_));
 sky130_fd_sc_hd__o21ai_0 _778_ (.A1(_221_),
    .A2(_325_),
    .B1(_327_),
    .Y(_067_));
 sky130_fd_sc_hd__nand2_1 _779_ (.A(net124),
    .B(_323_),
    .Y(_328_));
 sky130_fd_sc_hd__nor3_1 _780_ (.A(_289_),
    .B(_294_),
    .C(_328_),
    .Y(_329_));
 sky130_fd_sc_hd__o21ai_0 _781_ (.A1(_237_),
    .A2(_329_),
    .B1(_210_),
    .Y(_330_));
 sky130_fd_sc_hd__nand2_1 _782_ (.A(net54),
    .B(_266_),
    .Y(_331_));
 sky130_fd_sc_hd__o31ai_1 _783_ (.A1(net125),
    .A2(_295_),
    .A3(_328_),
    .B1(_331_),
    .Y(_332_));
 sky130_fd_sc_hd__a22o_1 _784_ (.A1(net125),
    .A2(_330_),
    .B1(_332_),
    .B2(_211_),
    .X(_068_));
 sky130_fd_sc_hd__nand3_1 _785_ (.A(net123),
    .B(net124),
    .C(net125),
    .Y(_333_));
 sky130_fd_sc_hd__or2_1 _786_ (.A(_317_),
    .B(_333_),
    .X(_334_));
 sky130_fd_sc_hd__nor4_1 _787_ (.A(_263_),
    .B(_251_),
    .C(_310_),
    .D(_334_),
    .Y(_335_));
 sky130_fd_sc_hd__o21ai_0 _788_ (.A1(_240_),
    .A2(_335_),
    .B1(_270_),
    .Y(_336_));
 sky130_fd_sc_hd__nor2_1 _789_ (.A(net126),
    .B(_256_),
    .Y(_337_));
 sky130_fd_sc_hd__a22oi_1 _790_ (.A1(net55),
    .A2(_191_),
    .B1(_335_),
    .B2(_337_),
    .Y(_338_));
 sky130_fd_sc_hd__o2bb2ai_1 _791_ (.A1_N(net126),
    .A2_N(_336_),
    .B1(_338_),
    .B2(_269_),
    .Y(_069_));
 sky130_fd_sc_hd__nor4b_1 _792_ (.A(_289_),
    .B(_294_),
    .C(_334_),
    .D_N(net126),
    .Y(_339_));
 sky130_fd_sc_hd__o21ai_0 _793_ (.A1(_240_),
    .A2(_339_),
    .B1(_270_),
    .Y(_340_));
 sky130_fd_sc_hd__nor2_1 _794_ (.A(net127),
    .B(_256_),
    .Y(_341_));
 sky130_fd_sc_hd__a22oi_1 _795_ (.A1(net56),
    .A2(_191_),
    .B1(_339_),
    .B2(_341_),
    .Y(_342_));
 sky130_fd_sc_hd__o2bb2ai_1 _796_ (.A1_N(net127),
    .A2_N(_340_),
    .B1(_342_),
    .B2(_269_),
    .Y(_070_));
 sky130_fd_sc_hd__nor2_1 _797_ (.A(_317_),
    .B(_333_),
    .Y(_343_));
 sky130_fd_sc_hd__nand3_1 _798_ (.A(net126),
    .B(net127),
    .C(_343_),
    .Y(_344_));
 sky130_fd_sc_hd__nor4_1 _799_ (.A(_250_),
    .B(_272_),
    .C(_291_),
    .D(_344_),
    .Y(_345_));
 sky130_fd_sc_hd__o21ai_0 _800_ (.A1(_237_),
    .A2(_345_),
    .B1(_210_),
    .Y(_346_));
 sky130_fd_sc_hd__nor2_1 _801_ (.A(net128),
    .B(_243_),
    .Y(_347_));
 sky130_fd_sc_hd__a22o_1 _802_ (.A1(net57),
    .A2(_266_),
    .B1(_345_),
    .B2(_347_),
    .X(_348_));
 sky130_fd_sc_hd__a22o_1 _803_ (.A1(net128),
    .A2(_346_),
    .B1(_348_),
    .B2(_211_),
    .X(_071_));
 sky130_fd_sc_hd__nand3_1 _804_ (.A(net126),
    .B(net127),
    .C(net128),
    .Y(_349_));
 sky130_fd_sc_hd__nor4_1 _805_ (.A(_289_),
    .B(_294_),
    .C(_334_),
    .D(_349_),
    .Y(_350_));
 sky130_fd_sc_hd__o21ai_0 _806_ (.A1(_240_),
    .A2(_350_),
    .B1(_270_),
    .Y(_351_));
 sky130_fd_sc_hd__nor2_1 _807_ (.A(net129),
    .B(_256_),
    .Y(_352_));
 sky130_fd_sc_hd__a22oi_1 _808_ (.A1(net58),
    .A2(_191_),
    .B1(_350_),
    .B2(_352_),
    .Y(_353_));
 sky130_fd_sc_hd__o2bb2ai_1 _809_ (.A1_N(net129),
    .A2_N(_351_),
    .B1(_353_),
    .B2(_269_),
    .Y(_072_));
 sky130_fd_sc_hd__nand4_1 _810_ (.A(net126),
    .B(net127),
    .C(net128),
    .D(net129),
    .Y(_354_));
 sky130_fd_sc_hd__nor3_1 _811_ (.A(net130),
    .B(_243_),
    .C(_354_),
    .Y(_355_));
 sky130_fd_sc_hd__a22oi_1 _812_ (.A1(net59),
    .A2(_266_),
    .B1(_335_),
    .B2(_355_),
    .Y(_356_));
 sky130_fd_sc_hd__nor4_1 _813_ (.A(_263_),
    .B(_310_),
    .C(_334_),
    .D(_354_),
    .Y(_357_));
 sky130_fd_sc_hd__a21oi_1 _814_ (.A1(_255_),
    .A2(_357_),
    .B1(_240_),
    .Y(_358_));
 sky130_fd_sc_hd__o21ai_0 _815_ (.A1(_219_),
    .A2(_358_),
    .B1(net130),
    .Y(_359_));
 sky130_fd_sc_hd__o21ai_0 _816_ (.A1(_221_),
    .A2(_356_),
    .B1(_359_),
    .Y(_073_));
 sky130_fd_sc_hd__and4_1 _817_ (.A(net126),
    .B(net127),
    .C(net128),
    .D(net129),
    .X(_360_));
 sky130_fd_sc_hd__nand2_1 _818_ (.A(net130),
    .B(_360_),
    .Y(_361_));
 sky130_fd_sc_hd__nor4_1 _819_ (.A(_289_),
    .B(_294_),
    .C(_334_),
    .D(_361_),
    .Y(_362_));
 sky130_fd_sc_hd__o21ai_0 _820_ (.A1(_237_),
    .A2(_362_),
    .B1(_210_),
    .Y(_363_));
 sky130_fd_sc_hd__nor2_1 _821_ (.A(net131),
    .B(_243_),
    .Y(_364_));
 sky130_fd_sc_hd__a22o_1 _822_ (.A1(net60),
    .A2(_190_),
    .B1(_362_),
    .B2(_364_),
    .X(_365_));
 sky130_fd_sc_hd__a22o_1 _823_ (.A1(net131),
    .A2(_363_),
    .B1(_365_),
    .B2(_270_),
    .X(_074_));
 sky130_fd_sc_hd__and3_1 _824_ (.A(net130),
    .B(net131),
    .C(_360_),
    .X(_366_));
 sky130_fd_sc_hd__nand2_1 _825_ (.A(_343_),
    .B(_366_),
    .Y(_367_));
 sky130_fd_sc_hd__nor4_1 _826_ (.A(_251_),
    .B(_272_),
    .C(_291_),
    .D(_367_),
    .Y(_368_));
 sky130_fd_sc_hd__o21ai_0 _827_ (.A1(_240_),
    .A2(_368_),
    .B1(_270_),
    .Y(_369_));
 sky130_fd_sc_hd__nor3_1 _828_ (.A(net132),
    .B(_237_),
    .C(_367_),
    .Y(_370_));
 sky130_fd_sc_hd__and2b_1 _829_ (.A_N(_149_),
    .B(net61),
    .X(_371_));
 sky130_fd_sc_hd__a21oi_1 _830_ (.A1(_300_),
    .A2(_370_),
    .B1(_371_),
    .Y(_372_));
 sky130_fd_sc_hd__o2bb2ai_1 _831_ (.A1_N(net132),
    .A2_N(_369_),
    .B1(_269_),
    .B2(_372_),
    .Y(_075_));
 sky130_fd_sc_hd__nand2b_1 _832_ (.A_N(_464_),
    .B(_428_),
    .Y(_373_));
 sky130_fd_sc_hd__a32oi_1 _833_ (.A1(_217_),
    .A2(_222_),
    .A3(_373_),
    .B1(_191_),
    .B2(net62),
    .Y(_374_));
 sky130_fd_sc_hd__nand2_1 _834_ (.A(net133),
    .B(_269_),
    .Y(_375_));
 sky130_fd_sc_hd__o21ai_0 _835_ (.A1(_221_),
    .A2(_374_),
    .B1(_375_),
    .Y(_076_));
 sky130_fd_sc_hd__nor4b_1 _836_ (.A(_289_),
    .B(_294_),
    .C(_367_),
    .D_N(net132),
    .Y(_376_));
 sky130_fd_sc_hd__o21ai_0 _837_ (.A1(_237_),
    .A2(_376_),
    .B1(_210_),
    .Y(_377_));
 sky130_fd_sc_hd__nor2_1 _838_ (.A(net134),
    .B(_243_),
    .Y(_378_));
 sky130_fd_sc_hd__a22o_1 _839_ (.A1(net63),
    .A2(_190_),
    .B1(_376_),
    .B2(_378_),
    .X(_379_));
 sky130_fd_sc_hd__a22o_1 _840_ (.A1(net134),
    .A2(_377_),
    .B1(_379_),
    .B2(_270_),
    .X(_077_));
 sky130_fd_sc_hd__nand4_1 _841_ (.A(net132),
    .B(net134),
    .C(_343_),
    .D(_366_),
    .Y(_380_));
 sky130_fd_sc_hd__nor4_1 _842_ (.A(_263_),
    .B(_251_),
    .C(_310_),
    .D(_380_),
    .Y(_381_));
 sky130_fd_sc_hd__o21ai_0 _843_ (.A1(_240_),
    .A2(_381_),
    .B1(_270_),
    .Y(_382_));
 sky130_fd_sc_hd__nor2_1 _844_ (.A(net135),
    .B(_237_),
    .Y(_383_));
 sky130_fd_sc_hd__a22oi_1 _845_ (.A1(net64),
    .A2(_213_),
    .B1(_381_),
    .B2(_383_),
    .Y(_384_));
 sky130_fd_sc_hd__o2bb2ai_1 _846_ (.A1_N(net135),
    .A2_N(_382_),
    .B1(_384_),
    .B2(_269_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _847_ (.A(net136),
    .B(_211_),
    .Y(_385_));
 sky130_fd_sc_hd__a21o_1 _848_ (.A1(_457_),
    .A2(_461_),
    .B1(_460_),
    .X(_386_));
 sky130_fd_sc_hd__a21oi_1 _849_ (.A1(_464_),
    .A2(_386_),
    .B1(_463_),
    .Y(_387_));
 sky130_fd_sc_hd__xnor2_1 _850_ (.A(_467_),
    .B(_387_),
    .Y(_388_));
 sky130_fd_sc_hd__a221oi_1 _851_ (.A1(net65),
    .A2(_213_),
    .B1(_217_),
    .B2(_388_),
    .C1(_219_),
    .Y(_389_));
 sky130_fd_sc_hd__nor2_1 _852_ (.A(_385_),
    .B(_389_),
    .Y(_079_));
 sky130_fd_sc_hd__nor2_1 _853_ (.A(net137),
    .B(_211_),
    .Y(_390_));
 sky130_fd_sc_hd__nand2b_1 _854_ (.A_N(_463_),
    .B(_222_),
    .Y(_391_));
 sky130_fd_sc_hd__a21oi_1 _855_ (.A1(_467_),
    .A2(_391_),
    .B1(_466_),
    .Y(_392_));
 sky130_fd_sc_hd__xnor2_1 _856_ (.A(_470_),
    .B(_392_),
    .Y(_393_));
 sky130_fd_sc_hd__a221oi_1 _857_ (.A1(net66),
    .A2(_213_),
    .B1(_217_),
    .B2(_393_),
    .C1(_219_),
    .Y(_394_));
 sky130_fd_sc_hd__nor2_1 _858_ (.A(_390_),
    .B(_394_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2_1 _859_ (.A(net138),
    .B(_211_),
    .Y(_395_));
 sky130_fd_sc_hd__xor2_1 _860_ (.A(_473_),
    .B(_247_),
    .X(_396_));
 sky130_fd_sc_hd__a221oi_1 _861_ (.A1(net67),
    .A2(_213_),
    .B1(_217_),
    .B2(_396_),
    .C1(_218_),
    .Y(_397_));
 sky130_fd_sc_hd__nor2_1 _862_ (.A(_395_),
    .B(_397_),
    .Y(_081_));
 sky130_fd_sc_hd__nor2_1 _863_ (.A(net139),
    .B(_211_),
    .Y(_398_));
 sky130_fd_sc_hd__and2_0 _864_ (.A(_225_),
    .B(_228_),
    .X(_399_));
 sky130_fd_sc_hd__xnor2_1 _865_ (.A(_230_),
    .B(_399_),
    .Y(_400_));
 sky130_fd_sc_hd__a221oi_1 _866_ (.A1(net68),
    .A2(_213_),
    .B1(_217_),
    .B2(_400_),
    .C1(_218_),
    .Y(_401_));
 sky130_fd_sc_hd__nor2_1 _867_ (.A(_398_),
    .B(_401_),
    .Y(_082_));
 sky130_fd_sc_hd__nor2_1 _868_ (.A(_472_),
    .B(_475_),
    .Y(_402_));
 sky130_fd_sc_hd__o211ai_1 _869_ (.A1(_244_),
    .A2(_245_),
    .B1(_402_),
    .C1(_246_),
    .Y(_403_));
 sky130_fd_sc_hd__or3_1 _870_ (.A(_473_),
    .B(_472_),
    .C(_475_),
    .X(_404_));
 sky130_fd_sc_hd__o211ai_1 _871_ (.A1(_230_),
    .A2(_475_),
    .B1(_403_),
    .C1(_404_),
    .Y(_405_));
 sky130_fd_sc_hd__xnor2_1 _872_ (.A(_226_),
    .B(_405_),
    .Y(_406_));
 sky130_fd_sc_hd__a221oi_1 _873_ (.A1(net69),
    .A2(_266_),
    .B1(_217_),
    .B2(_406_),
    .C1(_218_),
    .Y(_407_));
 sky130_fd_sc_hd__nor2_1 _874_ (.A(net140),
    .B(_211_),
    .Y(_408_));
 sky130_fd_sc_hd__nor2_1 _875_ (.A(_407_),
    .B(_408_),
    .Y(_083_));
 sky130_fd_sc_hd__nand2_1 _876_ (.A(_227_),
    .B(_261_),
    .Y(_409_));
 sky130_fd_sc_hd__o21ai_0 _877_ (.A1(_240_),
    .A2(_409_),
    .B1(_210_),
    .Y(_410_));
 sky130_fd_sc_hd__nor2_1 _878_ (.A(net141),
    .B(_237_),
    .Y(_411_));
 sky130_fd_sc_hd__a22oi_1 _879_ (.A1(net70),
    .A2(_213_),
    .B1(_409_),
    .B2(_411_),
    .Y(_412_));
 sky130_fd_sc_hd__o2bb2ai_1 _880_ (.A1_N(net141),
    .A2_N(_410_),
    .B1(_412_),
    .B2(_269_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _881_ (.A(net142),
    .B(_237_),
    .Y(_413_));
 sky130_fd_sc_hd__a32oi_1 _882_ (.A1(net141),
    .A2(_255_),
    .A3(_413_),
    .B1(net71),
    .B2(_191_),
    .Y(_414_));
 sky130_fd_sc_hd__a21oi_1 _883_ (.A1(net141),
    .A2(_255_),
    .B1(_256_),
    .Y(_415_));
 sky130_fd_sc_hd__o21ai_0 _884_ (.A1(_219_),
    .A2(_415_),
    .B1(net142),
    .Y(_416_));
 sky130_fd_sc_hd__o21ai_0 _885_ (.A1(_221_),
    .A2(_414_),
    .B1(_416_),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_2 _886_ (.A(net184),
    .B(_130_),
    .Y(_417_));
 sky130_fd_sc_hd__clkbuf_4 _887_ (.A(_417_),
    .X(_418_));
 sky130_fd_sc_hd__mux2_1 _888_ (.A0(net185),
    .A1(net3),
    .S(_418_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _889_ (.A0(net186),
    .A1(net4),
    .S(_418_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _890_ (.A0(net187),
    .A1(net5),
    .S(_418_),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _891_ (.A0(net188),
    .A1(net6),
    .S(_418_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _892_ (.A0(net189),
    .A1(net7),
    .S(_418_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _893_ (.A0(net190),
    .A1(net8),
    .S(_418_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _894_ (.A0(net191),
    .A1(net9),
    .S(_418_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _895_ (.A0(net192),
    .A1(net10),
    .S(_418_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _896_ (.A0(net193),
    .A1(net11),
    .S(_418_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _897_ (.A0(net194),
    .A1(net12),
    .S(_418_),
    .X(_095_));
 sky130_fd_sc_hd__clkbuf_4 _898_ (.A(_417_),
    .X(_419_));
 sky130_fd_sc_hd__mux2_1 _899_ (.A0(net195),
    .A1(net13),
    .S(_419_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _900_ (.A0(net196),
    .A1(net14),
    .S(_419_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _901_ (.A0(net197),
    .A1(net15),
    .S(_419_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _902_ (.A0(net198),
    .A1(net16),
    .S(_419_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _903_ (.A0(net199),
    .A1(net17),
    .S(_419_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _904_ (.A0(net200),
    .A1(net18),
    .S(_419_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _905_ (.A0(net201),
    .A1(net19),
    .S(_419_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _906_ (.A0(net202),
    .A1(net20),
    .S(_419_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _907_ (.A0(net203),
    .A1(net21),
    .S(_419_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _908_ (.A0(net204),
    .A1(net22),
    .S(_419_),
    .X(_105_));
 sky130_fd_sc_hd__clkbuf_4 _909_ (.A(_417_),
    .X(_420_));
 sky130_fd_sc_hd__mux2_1 _910_ (.A0(net205),
    .A1(net23),
    .S(_420_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _911_ (.A0(net206),
    .A1(net24),
    .S(_420_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _912_ (.A0(net207),
    .A1(net25),
    .S(_420_),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _913_ (.A0(net208),
    .A1(net26),
    .S(_420_),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _914_ (.A0(net209),
    .A1(net27),
    .S(_420_),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _915_ (.A0(net210),
    .A1(net28),
    .S(_420_),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _916_ (.A0(net211),
    .A1(net29),
    .S(_420_),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _917_ (.A0(net212),
    .A1(net30),
    .S(_420_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _918_ (.A0(net213),
    .A1(net31),
    .S(_420_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _919_ (.A0(net214),
    .A1(net32),
    .S(_420_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _920_ (.A0(net215),
    .A1(net33),
    .S(_417_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _921_ (.A0(net216),
    .A1(net34),
    .S(_417_),
    .X(_117_));
 sky130_fd_sc_hd__xor2_1 _922_ (.A(_122_),
    .B(_125_),
    .X(_421_));
 sky130_fd_sc_hd__o22a_1 _923_ (.A1(net217),
    .A2(_143_),
    .B1(_421_),
    .B2(_123_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _924_ (.A0(net218),
    .A1(net37),
    .S(_143_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _925_ (.A0(net219),
    .A1(net38),
    .S(_143_),
    .X(_120_));
 sky130_fd_sc_hd__fa_1 _926_ (.A(_425_),
    .B(_426_),
    .CIN(_427_),
    .COUT(_428_),
    .SUM(_429_));
 sky130_fd_sc_hd__ha_1 _927_ (.A(\burst_count[7] ),
    .B(_430_),
    .COUT(_431_),
    .SUM(_432_));
 sky130_fd_sc_hd__ha_1 _928_ (.A(\burst_count[6] ),
    .B(_433_),
    .COUT(_434_),
    .SUM(_435_));
 sky130_fd_sc_hd__ha_1 _929_ (.A(\burst_count[5] ),
    .B(_436_),
    .COUT(_437_),
    .SUM(_438_));
 sky130_fd_sc_hd__ha_1 _930_ (.A(_439_),
    .B(_440_),
    .COUT(_441_),
    .SUM(_442_));
 sky130_fd_sc_hd__ha_1 _931_ (.A(\burst_count[4] ),
    .B(_442_),
    .COUT(_443_),
    .SUM(_444_));
 sky130_fd_sc_hd__ha_1 _932_ (.A(\burst_count[3] ),
    .B(_445_),
    .COUT(_446_),
    .SUM(_447_));
 sky130_fd_sc_hd__ha_1 _933_ (.A(_448_),
    .B(_449_),
    .COUT(_450_),
    .SUM(_451_));
 sky130_fd_sc_hd__ha_1 _934_ (.A(\burst_count[2] ),
    .B(_451_),
    .COUT(_452_),
    .SUM(_453_));
 sky130_fd_sc_hd__ha_1 _935_ (.A(\burst_count[1] ),
    .B(\burst_total[0] ),
    .COUT(_454_),
    .SUM(_455_));
 sky130_fd_sc_hd__ha_1 _936_ (.A(net111),
    .B(_456_),
    .COUT(_457_),
    .SUM(_458_));
 sky130_fd_sc_hd__ha_1 _937_ (.A(net122),
    .B(_459_),
    .COUT(_460_),
    .SUM(_461_));
 sky130_fd_sc_hd__ha_1 _938_ (.A(net133),
    .B(_462_),
    .COUT(_463_),
    .SUM(_464_));
 sky130_fd_sc_hd__ha_1 _939_ (.A(net136),
    .B(_465_),
    .COUT(_466_),
    .SUM(_467_));
 sky130_fd_sc_hd__ha_1 _940_ (.A(net137),
    .B(_468_),
    .COUT(_469_),
    .SUM(_470_));
 sky130_fd_sc_hd__ha_1 _941_ (.A(net138),
    .B(_471_),
    .COUT(_472_),
    .SUM(_473_));
 sky130_fd_sc_hd__ha_1 _942_ (.A(net139),
    .B(_474_),
    .COUT(_475_),
    .SUM(_476_));
 sky130_fd_sc_hd__ha_1 _943_ (.A(net140),
    .B(_477_),
    .COUT(_478_),
    .SUM(_479_));
 sky130_fd_sc_hd__ha_1 _944_ (.A(\burst_count[0] ),
    .B(\burst_count[1] ),
    .COUT(_480_),
    .SUM(_481_));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(\burst_count[0] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[1]$_DFFE_PN0P_  (.D(_001_),
    .Q(\burst_count[1] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \burst_count[2]$_DFFE_PN0P_  (.D(_002_),
    .Q(\burst_count[2] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[3]$_DFFE_PN0P_  (.D(_003_),
    .Q(\burst_count[3] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[4]$_DFFE_PN0P_  (.D(_004_),
    .Q(\burst_count[4] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[5]$_DFFE_PN0P_  (.D(_005_),
    .Q(\burst_count[5] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[6]$_DFFE_PN0P_  (.D(_006_),
    .Q(\burst_count[6] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_count[7]$_DFFE_PN0P_  (.D(_007_),
    .Q(\burst_count[7] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_total[0]$_DFFE_PN0P_  (.D(_008_),
    .Q(\burst_total[0] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_total[2]$_DFFE_PN0P_  (.D(_009_),
    .Q(\burst_total[2] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_total[3]$_DFFE_PN0P_  (.D(_010_),
    .Q(\burst_total[3] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \burst_total[4]$_DFFE_PN0P_  (.D(_011_),
    .Q(\burst_total[4] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hburst[0]$_DFFE_PN0P_  (.D(_012_),
    .Q(net143),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hburst[1]$_DFFE_PN0P_  (.D(_013_),
    .Q(net144),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hburst[2]$_DFFE_PN0P_  (.D(_014_),
    .Q(net145),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hbusreq$_DFFE_PN0P_  (.D(_015_),
    .Q(net146),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \hsize[0]$_DFFE_PN0P_  (.D(_016_),
    .Q(net147),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \hsize[1]$_DFFE_PN0P_  (.D(_017_),
    .Q(net148),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \hsize[2]$_DFFE_PN0P_  (.D(_018_),
    .Q(net149),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \htrans[0]$_DFFE_PN0P_  (.D(_019_),
    .Q(net150),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \htrans[1]$_DFFE_PN0P_  (.D(_020_),
    .Q(net151),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[0]$_DFFE_PN0P_  (.D(_021_),
    .Q(net152),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[10]$_DFFE_PN0P_  (.D(_022_),
    .Q(net153),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[11]$_DFFE_PN0P_  (.D(_023_),
    .Q(net154),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[12]$_DFFE_PN0P_  (.D(_024_),
    .Q(net155),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[13]$_DFFE_PN0P_  (.D(_025_),
    .Q(net156),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[14]$_DFFE_PN0P_  (.D(_026_),
    .Q(net157),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[15]$_DFFE_PN0P_  (.D(_027_),
    .Q(net158),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[16]$_DFFE_PN0P_  (.D(_028_),
    .Q(net159),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[17]$_DFFE_PN0P_  (.D(_029_),
    .Q(net160),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[18]$_DFFE_PN0P_  (.D(_030_),
    .Q(net161),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[19]$_DFFE_PN0P_  (.D(_031_),
    .Q(net162),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[1]$_DFFE_PN0P_  (.D(_032_),
    .Q(net163),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[20]$_DFFE_PN0P_  (.D(_033_),
    .Q(net164),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[21]$_DFFE_PN0P_  (.D(_034_),
    .Q(net165),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[22]$_DFFE_PN0P_  (.D(_035_),
    .Q(net166),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[23]$_DFFE_PN0P_  (.D(_036_),
    .Q(net167),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[24]$_DFFE_PN0P_  (.D(_037_),
    .Q(net168),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[25]$_DFFE_PN0P_  (.D(_038_),
    .Q(net169),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[26]$_DFFE_PN0P_  (.D(_039_),
    .Q(net170),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[27]$_DFFE_PN0P_  (.D(_040_),
    .Q(net171),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[28]$_DFFE_PN0P_  (.D(_041_),
    .Q(net172),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[29]$_DFFE_PN0P_  (.D(_042_),
    .Q(net173),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[2]$_DFFE_PN0P_  (.D(_043_),
    .Q(net174),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[30]$_DFFE_PN0P_  (.D(_044_),
    .Q(net175),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[31]$_DFFE_PN0P_  (.D(_045_),
    .Q(net176),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[3]$_DFFE_PN0P_  (.D(_046_),
    .Q(net177),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[4]$_DFFE_PN0P_  (.D(_047_),
    .Q(net178),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[5]$_DFFE_PN0P_  (.D(_048_),
    .Q(net179),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[6]$_DFFE_PN0P_  (.D(_049_),
    .Q(net180),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[7]$_DFFE_PN0P_  (.D(_050_),
    .Q(net181),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[8]$_DFFE_PN0P_  (.D(_051_),
    .Q(net182),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \hwdata[9]$_DFFE_PN0P_  (.D(_052_),
    .Q(net183),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \hwrite$_DFFE_PN0P_  (.D(_053_),
    .Q(net184),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[0]$_DFFE_PN0P_  (.D(_054_),
    .Q(net111),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[10]$_DFFE_PN0P_  (.D(_055_),
    .Q(net112),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[11]$_DFFE_PN0P_  (.D(_056_),
    .Q(net113),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[12]$_DFFE_PN0P_  (.D(_057_),
    .Q(net114),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[13]$_DFFE_PN0P_  (.D(_058_),
    .Q(net115),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[14]$_DFFE_PN0P_  (.D(_059_),
    .Q(net116),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[15]$_DFFE_PN0P_  (.D(_060_),
    .Q(net117),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[16]$_DFFE_PN0P_  (.D(_061_),
    .Q(net118),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[17]$_DFFE_PN0P_  (.D(_062_),
    .Q(net119),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[18]$_DFFE_PN0P_  (.D(_063_),
    .Q(net120),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[19]$_DFFE_PN0P_  (.D(_064_),
    .Q(net121),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[1]$_DFFE_PN0P_  (.D(_065_),
    .Q(net122),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[20]$_DFFE_PN0P_  (.D(_066_),
    .Q(net123),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[21]$_DFFE_PN0P_  (.D(_067_),
    .Q(net124),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[22]$_DFFE_PN0P_  (.D(_068_),
    .Q(net125),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[23]$_DFFE_PN0P_  (.D(_069_),
    .Q(net126),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[24]$_DFFE_PN0P_  (.D(_070_),
    .Q(net127),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[25]$_DFFE_PN0P_  (.D(_071_),
    .Q(net128),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[26]$_DFFE_PN0P_  (.D(_072_),
    .Q(net129),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[27]$_DFFE_PN0P_  (.D(_073_),
    .Q(net130),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[28]$_DFFE_PN0P_  (.D(_074_),
    .Q(net131),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[29]$_DFFE_PN0P_  (.D(_075_),
    .Q(net132),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[2]$_DFFE_PN0P_  (.D(_076_),
    .Q(net133),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[30]$_DFFE_PN0P_  (.D(_077_),
    .Q(net134),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[31]$_DFFE_PN0P_  (.D(_078_),
    .Q(net135),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[3]$_DFFE_PN0P_  (.D(_079_),
    .Q(net136),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[4]$_DFFE_PN0P_  (.D(_080_),
    .Q(net137),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[5]$_DFFE_PN0P_  (.D(_081_),
    .Q(net138),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[6]$_DFFE_PN0P_  (.D(_082_),
    .Q(net139),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[7]$_DFFE_PN0P_  (.D(_083_),
    .Q(net140),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \next_addr[8]$_DFFE_PN0P_  (.D(_084_),
    .Q(net141),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \next_addr[9]$_DFFE_PN0P_  (.D(_085_),
    .Q(net142),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[0]$_DFFE_PN0P_  (.D(_086_),
    .Q(net185),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[10]$_DFFE_PN0P_  (.D(_087_),
    .Q(net186),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[11]$_DFFE_PN0P_  (.D(_088_),
    .Q(net187),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[12]$_DFFE_PN0P_  (.D(_089_),
    .Q(net188),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[13]$_DFFE_PN0P_  (.D(_090_),
    .Q(net189),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[14]$_DFFE_PN0P_  (.D(_091_),
    .Q(net190),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[15]$_DFFE_PN0P_  (.D(_092_),
    .Q(net191),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[16]$_DFFE_PN0P_  (.D(_093_),
    .Q(net192),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[17]$_DFFE_PN0P_  (.D(_094_),
    .Q(net193),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[18]$_DFFE_PN0P_  (.D(_095_),
    .Q(net194),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[19]$_DFFE_PN0P_  (.D(_096_),
    .Q(net195),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[1]$_DFFE_PN0P_  (.D(_097_),
    .Q(net196),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[20]$_DFFE_PN0P_  (.D(_098_),
    .Q(net197),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[21]$_DFFE_PN0P_  (.D(_099_),
    .Q(net198),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[22]$_DFFE_PN0P_  (.D(_100_),
    .Q(net199),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[23]$_DFFE_PN0P_  (.D(_101_),
    .Q(net200),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[24]$_DFFE_PN0P_  (.D(_102_),
    .Q(net201),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[25]$_DFFE_PN0P_  (.D(_103_),
    .Q(net202),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[26]$_DFFE_PN0P_  (.D(_104_),
    .Q(net203),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[27]$_DFFE_PN0P_  (.D(_105_),
    .Q(net204),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[28]$_DFFE_PN0P_  (.D(_106_),
    .Q(net205),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[29]$_DFFE_PN0P_  (.D(_107_),
    .Q(net206),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[2]$_DFFE_PN0P_  (.D(_108_),
    .Q(net207),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[30]$_DFFE_PN0P_  (.D(_109_),
    .Q(net208),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[31]$_DFFE_PN0P_  (.D(_110_),
    .Q(net209),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[3]$_DFFE_PN0P_  (.D(_111_),
    .Q(net210),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[4]$_DFFE_PN0P_  (.D(_112_),
    .Q(net211),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[5]$_DFFE_PN0P_  (.D(_113_),
    .Q(net212),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[6]$_DFFE_PN0P_  (.D(_114_),
    .Q(net213),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[7]$_DFFE_PN0P_  (.D(_115_),
    .Q(net214),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[8]$_DFFE_PN0P_  (.D(_116_),
    .Q(net215),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[9]$_DFFE_PN0P_  (.D(_117_),
    .Q(net216),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFF_PN0_  (.D(_422_),
    .Q(\state[0] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \state[1]$_DFF_PN0_  (.D(_423_),
    .Q(\state[1] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \state[2]$_DFF_PN0_  (.D(_424_),
    .Q(\state[2] ),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \trans_done$_DFFE_PN0P_  (.D(_118_),
    .Q(net217),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \trans_resp[0]$_DFFE_PN0P_  (.D(_119_),
    .Q(net218),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \trans_resp[1]$_DFFE_PN0P_  (.D(_120_),
    .Q(net219),
    .RESET_B(net36),
    .CLK(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_139 ();
 sky130_fd_sc_hd__buf_16 input1 (.A(hclk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(hgrant),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(hrdata[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(hrdata[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(hrdata[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(hrdata[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(hrdata[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(hrdata[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(hrdata[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(hrdata[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(hrdata[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(hrdata[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(hrdata[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(hrdata[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(hrdata[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(hrdata[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(hrdata[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(hrdata[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(hrdata[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(hrdata[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(hrdata[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(hrdata[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(hrdata[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(hrdata[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(hrdata[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(hrdata[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(hrdata[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(hrdata[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(hrdata[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(hrdata[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(hrdata[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(hrdata[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(hrdata[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(hrdata[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(hready),
    .X(net35));
 sky130_fd_sc_hd__buf_16 input36 (.A(hreset),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(hresp[0]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(hresp[1]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(start_trans),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(trans_addr[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(trans_addr[10]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(trans_addr[11]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(trans_addr[12]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(trans_addr[13]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(trans_addr[14]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(trans_addr[15]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(trans_addr[16]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(trans_addr[17]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(trans_addr[18]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(trans_addr[19]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(trans_addr[1]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(trans_addr[20]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(trans_addr[21]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(trans_addr[22]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(trans_addr[23]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(trans_addr[24]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(trans_addr[25]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(trans_addr[26]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(trans_addr[27]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(trans_addr[28]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(trans_addr[29]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(trans_addr[2]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(trans_addr[30]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(trans_addr[31]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(trans_addr[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(trans_addr[4]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(trans_addr[5]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(trans_addr[6]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(trans_addr[7]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(trans_addr[8]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(trans_addr[9]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(trans_burst[0]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(trans_burst[1]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(trans_burst[2]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(trans_size[0]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(trans_size[1]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(trans_size[2]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(trans_write),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(write_data[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(write_data[10]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(write_data[11]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(write_data[12]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(write_data[13]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(write_data[14]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(write_data[15]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(write_data[16]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(write_data[17]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(write_data[18]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(write_data[19]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(write_data[1]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(write_data[20]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(write_data[21]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(write_data[22]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(write_data[23]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(write_data[24]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(write_data[25]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(write_data[26]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(write_data[27]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(write_data[28]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(write_data[29]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(write_data[2]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(write_data[30]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(write_data[31]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(write_data[3]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(write_data[4]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(write_data[5]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(write_data[6]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(write_data[7]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(write_data[8]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(write_data[9]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net111),
    .X(haddr[0]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net112),
    .X(haddr[10]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net113),
    .X(haddr[11]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net114),
    .X(haddr[12]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net115),
    .X(haddr[13]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net116),
    .X(haddr[14]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net117),
    .X(haddr[15]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net118),
    .X(haddr[16]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net119),
    .X(haddr[17]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net120),
    .X(haddr[18]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net121),
    .X(haddr[19]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net122),
    .X(haddr[1]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net123),
    .X(haddr[20]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net124),
    .X(haddr[21]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net125),
    .X(haddr[22]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net126),
    .X(haddr[23]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net127),
    .X(haddr[24]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net128),
    .X(haddr[25]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net129),
    .X(haddr[26]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net130),
    .X(haddr[27]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net131),
    .X(haddr[28]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net132),
    .X(haddr[29]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net133),
    .X(haddr[2]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net134),
    .X(haddr[30]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net135),
    .X(haddr[31]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net136),
    .X(haddr[3]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net137),
    .X(haddr[4]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net138),
    .X(haddr[5]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net139),
    .X(haddr[6]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net140),
    .X(haddr[7]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net141),
    .X(haddr[8]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net142),
    .X(haddr[9]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net143),
    .X(hburst[0]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net144),
    .X(hburst[1]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net145),
    .X(hburst[2]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net146),
    .X(hbusreq));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net147),
    .X(hsize[0]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net148),
    .X(hsize[1]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net149),
    .X(hsize[2]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(htrans[0]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net151),
    .X(htrans[1]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net152),
    .X(hwdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net153),
    .X(hwdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net154),
    .X(hwdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net155),
    .X(hwdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net156),
    .X(hwdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net157),
    .X(hwdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net158),
    .X(hwdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net159),
    .X(hwdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net160),
    .X(hwdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net161),
    .X(hwdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net162),
    .X(hwdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net163),
    .X(hwdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net164),
    .X(hwdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net165),
    .X(hwdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net166),
    .X(hwdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net167),
    .X(hwdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net168),
    .X(hwdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net169),
    .X(hwdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net170),
    .X(hwdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net171),
    .X(hwdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net172),
    .X(hwdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net173),
    .X(hwdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net174),
    .X(hwdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net175),
    .X(hwdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net176),
    .X(hwdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net177),
    .X(hwdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net178),
    .X(hwdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net179),
    .X(hwdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net180),
    .X(hwdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net181),
    .X(hwdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net182),
    .X(hwdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net183),
    .X(hwdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net184),
    .X(hwrite));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net185),
    .X(read_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net186),
    .X(read_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net187),
    .X(read_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net188),
    .X(read_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net189),
    .X(read_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net190),
    .X(read_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net191),
    .X(read_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net192),
    .X(read_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net193),
    .X(read_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net194),
    .X(read_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net195),
    .X(read_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net196),
    .X(read_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net197),
    .X(read_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net198),
    .X(read_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net199),
    .X(read_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net200),
    .X(read_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net201),
    .X(read_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net202),
    .X(read_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net203),
    .X(read_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net204),
    .X(read_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net205),
    .X(read_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net206),
    .X(read_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net207),
    .X(read_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net208),
    .X(read_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net209),
    .X(read_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net210),
    .X(read_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net211),
    .X(read_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net212),
    .X(read_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net213),
    .X(read_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net214),
    .X(read_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net215),
    .X(read_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net216),
    .X(read_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net217),
    .X(trans_done));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net218),
    .X(trans_resp[0]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net219),
    .X(trans_resp[1]));
 sky130_fd_sc_hd__fill_2 FILLER_0_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_231 ();
endmodule
