module power_domain_controller (clk,
    rst_n,
    start_transition,
    transition_done,
    domain_clock_on,
    domain_enable,
    domain_isolate,
    domain_isolation_on,
    domain_power_on,
    domain_reset_n,
    domain_status,
    domain_transition);
 input clk;
 input rst_n;
 input start_transition;
 output transition_done;
 output [3:0] domain_clock_on;
 input [3:0] domain_enable;
 input [3:0] domain_isolate;
 output [3:0] domain_isolation_on;
 output [3:0] domain_power_on;
 output [3:0] domain_reset_n;
 output [3:0] domain_status;
 output [3:0] domain_transition;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire \delay_counter[0] ;
 wire \delay_counter[1] ;
 wire \delay_counter[2] ;
 wire \delay_counter[3] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \target_status[0] ;
 wire \target_status[1] ;
 wire \target_status[2] ;
 wire \target_status[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net37;

 sky130_fd_sc_hd__inv_1 _152_ (.A(\delay_counter[0] ),
    .Y(_146_));
 sky130_fd_sc_hd__inv_1 _153_ (.A(\delay_counter[1] ),
    .Y(_147_));
 sky130_fd_sc_hd__clkbuf_4 _154_ (.A(\state[0] ),
    .X(_139_));
 sky130_fd_sc_hd__clkinvlp_4 _155_ (.A(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__and3_1 _156_ (.A(\state[2] ),
    .B(\state[1] ),
    .C(_140_),
    .X(_141_));
 sky130_fd_sc_hd__nand2_1 _157_ (.A(net35),
    .B(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__mux2_1 _158_ (.A0(\target_status[3] ),
    .A1(net31),
    .S(_142_),
    .X(_000_));
 sky130_fd_sc_hd__nand2_1 _159_ (.A(net34),
    .B(_141_),
    .Y(_143_));
 sky130_fd_sc_hd__mux2_1 _160_ (.A0(\target_status[2] ),
    .A1(net30),
    .S(_143_),
    .X(_001_));
 sky130_fd_sc_hd__nand2_1 _161_ (.A(net33),
    .B(_141_),
    .Y(_144_));
 sky130_fd_sc_hd__mux2_1 _162_ (.A0(\target_status[1] ),
    .A1(net29),
    .S(_144_),
    .X(_002_));
 sky130_fd_sc_hd__nand2_1 _163_ (.A(net32),
    .B(_141_),
    .Y(_145_));
 sky130_fd_sc_hd__mux2_1 _164_ (.A0(\target_status[0] ),
    .A1(net28),
    .S(_145_),
    .X(_003_));
 sky130_fd_sc_hd__nor2_2 _165_ (.A(\state[1] ),
    .B(\state[0] ),
    .Y(_036_));
 sky130_fd_sc_hd__and2_1 _166_ (.A(\state[2] ),
    .B(_036_),
    .X(_037_));
 sky130_fd_sc_hd__nand2_1 _167_ (.A(net35),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(\target_status[3] ),
    .A1(net15),
    .S(_038_),
    .X(_004_));
 sky130_fd_sc_hd__nand2_1 _169_ (.A(net34),
    .B(_037_),
    .Y(_039_));
 sky130_fd_sc_hd__mux2_1 _170_ (.A0(\target_status[2] ),
    .A1(net14),
    .S(_039_),
    .X(_005_));
 sky130_fd_sc_hd__nand2_1 _171_ (.A(net33),
    .B(_037_),
    .Y(_040_));
 sky130_fd_sc_hd__mux2_1 _172_ (.A0(\target_status[1] ),
    .A1(net13),
    .S(_040_),
    .X(_006_));
 sky130_fd_sc_hd__nand2_1 _173_ (.A(net32),
    .B(_037_),
    .Y(_041_));
 sky130_fd_sc_hd__mux2_1 _174_ (.A0(\target_status[0] ),
    .A1(net12),
    .S(_041_),
    .X(_007_));
 sky130_fd_sc_hd__nor3b_4 _175_ (.A(\state[2] ),
    .B(_139_),
    .C_N(\state[1] ),
    .Y(_042_));
 sky130_fd_sc_hd__nand2_1 _176_ (.A(net35),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__mux2_1 _177_ (.A0(\target_status[3] ),
    .A1(net23),
    .S(_043_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _178_ (.A(net34),
    .B(_042_),
    .Y(_044_));
 sky130_fd_sc_hd__mux2_1 _179_ (.A0(\target_status[2] ),
    .A1(net22),
    .S(_044_),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _180_ (.A(net33),
    .B(_042_),
    .Y(_045_));
 sky130_fd_sc_hd__mux2_1 _181_ (.A0(\target_status[1] ),
    .A1(net21),
    .S(_045_),
    .X(_010_));
 sky130_fd_sc_hd__nand2_1 _182_ (.A(net32),
    .B(_042_),
    .Y(_046_));
 sky130_fd_sc_hd__mux2_1 _183_ (.A0(\target_status[0] ),
    .A1(net20),
    .S(_046_),
    .X(_011_));
 sky130_fd_sc_hd__buf_2 _184_ (.A(\state[2] ),
    .X(_047_));
 sky130_fd_sc_hd__buf_2 _185_ (.A(_047_),
    .X(_048_));
 sky130_fd_sc_hd__buf_6 _186_ (.A(\delay_counter[2] ),
    .X(_049_));
 sky130_fd_sc_hd__nor3b_2 _187_ (.A(_049_),
    .B(\delay_counter[3] ),
    .C_N(_150_),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _188_ (.A(\delay_counter[0] ),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _189_ (.A(net11),
    .B(_146_),
    .Y(_052_));
 sky130_fd_sc_hd__or3b_2 _190_ (.A(\delay_counter[2] ),
    .B(\delay_counter[3] ),
    .C_N(_150_),
    .X(_053_));
 sky130_fd_sc_hd__buf_2 _191_ (.A(\state[1] ),
    .X(_054_));
 sky130_fd_sc_hd__inv_1 _192_ (.A(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__a21oi_1 _193_ (.A1(\delay_counter[0] ),
    .A2(_053_),
    .B1(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__a221oi_1 _194_ (.A1(_139_),
    .A2(_051_),
    .B1(_052_),
    .B2(_036_),
    .C1(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__o21ai_0 _195_ (.A1(_140_),
    .A2(_053_),
    .B1(_055_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2b_1 _196_ (.A(_054_),
    .B_N(\state[2] ),
    .Y(_059_));
 sky130_fd_sc_hd__a32oi_1 _197_ (.A1(_048_),
    .A2(\delay_counter[0] ),
    .A3(_058_),
    .B1(_059_),
    .B2(_051_),
    .Y(_060_));
 sky130_fd_sc_hd__xnor2_2 _198_ (.A(net5),
    .B(net31),
    .Y(_061_));
 sky130_fd_sc_hd__xnor2_2 _199_ (.A(net2),
    .B(net28),
    .Y(_062_));
 sky130_fd_sc_hd__xnor2_2 _200_ (.A(net4),
    .B(net30),
    .Y(_063_));
 sky130_fd_sc_hd__xnor2_2 _201_ (.A(net3),
    .B(net29),
    .Y(_064_));
 sky130_fd_sc_hd__nand4_1 _202_ (.A(_061_),
    .B(_062_),
    .C(_063_),
    .D(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__or3_1 _203_ (.A(\state[2] ),
    .B(\state[1] ),
    .C(\state[0] ),
    .X(_066_));
 sky130_fd_sc_hd__or3_1 _204_ (.A(_146_),
    .B(_065_),
    .C(_066_),
    .X(_067_));
 sky130_fd_sc_hd__o211ai_1 _205_ (.A1(_048_),
    .A2(_057_),
    .B1(_060_),
    .C1(_067_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _206_ (.A(_149_),
    .B(_053_),
    .Y(_068_));
 sky130_fd_sc_hd__nand3_1 _207_ (.A(_047_),
    .B(_147_),
    .C(_050_),
    .Y(_069_));
 sky130_fd_sc_hd__o21ai_0 _208_ (.A1(_047_),
    .A2(_068_),
    .B1(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__inv_1 _209_ (.A(net11),
    .Y(_071_));
 sky130_fd_sc_hd__a41oi_4 _210_ (.A1(_061_),
    .A2(_062_),
    .A3(_063_),
    .A4(_064_),
    .B1(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__nor3_1 _211_ (.A(\delay_counter[1] ),
    .B(_066_),
    .C(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__nand2_1 _212_ (.A(_047_),
    .B(_054_),
    .Y(_074_));
 sky130_fd_sc_hd__nand3_1 _213_ (.A(_149_),
    .B(_053_),
    .C(_059_),
    .Y(_075_));
 sky130_fd_sc_hd__o21ai_0 _214_ (.A1(_149_),
    .A2(_050_),
    .B1(_042_),
    .Y(_076_));
 sky130_fd_sc_hd__o211ai_1 _215_ (.A1(\delay_counter[1] ),
    .A2(_074_),
    .B1(_075_),
    .C1(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__a211oi_1 _216_ (.A1(_139_),
    .A2(_070_),
    .B1(_073_),
    .C1(_077_),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _217_ (.A(_148_),
    .B(_036_),
    .Y(_078_));
 sky130_fd_sc_hd__nand2b_1 _218_ (.A_N(_054_),
    .B(_148_),
    .Y(_079_));
 sky130_fd_sc_hd__o21ai_0 _219_ (.A1(_047_),
    .A2(_078_),
    .B1(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2b_1 _220_ (.A(\delay_counter[3] ),
    .B_N(_150_),
    .Y(_081_));
 sky130_fd_sc_hd__nand2_1 _221_ (.A(_139_),
    .B(_148_),
    .Y(_082_));
 sky130_fd_sc_hd__or3_1 _222_ (.A(_049_),
    .B(_081_),
    .C(_082_),
    .X(_083_));
 sky130_fd_sc_hd__nor3b_1 _223_ (.A(_139_),
    .B(_049_),
    .C_N(_054_),
    .Y(_084_));
 sky130_fd_sc_hd__o21ai_0 _224_ (.A1(_148_),
    .A2(_081_),
    .B1(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__nand3_1 _225_ (.A(_055_),
    .B(_140_),
    .C(_049_),
    .Y(_086_));
 sky130_fd_sc_hd__a31o_1 _226_ (.A1(_083_),
    .A2(_085_),
    .A3(_086_),
    .B1(_047_),
    .X(_087_));
 sky130_fd_sc_hd__nor3_1 _227_ (.A(_049_),
    .B(_081_),
    .C(_079_),
    .Y(_088_));
 sky130_fd_sc_hd__a21boi_0 _228_ (.A1(_148_),
    .A2(_074_),
    .B1_N(_049_),
    .Y(_089_));
 sky130_fd_sc_hd__a21oi_1 _229_ (.A1(_048_),
    .A2(_088_),
    .B1(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__a32oi_1 _230_ (.A1(_049_),
    .A2(_072_),
    .A3(_080_),
    .B1(_087_),
    .B2(_090_),
    .Y(_014_));
 sky130_fd_sc_hd__nor3_1 _231_ (.A(_150_),
    .B(\delay_counter[0] ),
    .C(\delay_counter[1] ),
    .Y(_091_));
 sky130_fd_sc_hd__a21oi_1 _232_ (.A1(_055_),
    .A2(_150_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__o31ai_1 _233_ (.A1(_049_),
    .A2(\delay_counter[0] ),
    .A3(\delay_counter[1] ),
    .B1(\delay_counter[3] ),
    .Y(_093_));
 sky130_fd_sc_hd__o31a_1 _234_ (.A1(_049_),
    .A2(\delay_counter[3] ),
    .A3(_092_),
    .B1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__nand3b_1 _235_ (.A_N(_047_),
    .B(\delay_counter[3] ),
    .C(_036_),
    .Y(_095_));
 sky130_fd_sc_hd__nor2_1 _236_ (.A(\delay_counter[3] ),
    .B(_150_),
    .Y(_096_));
 sky130_fd_sc_hd__nor4_1 _237_ (.A(\state[1] ),
    .B(_049_),
    .C(\delay_counter[0] ),
    .D(\delay_counter[1] ),
    .Y(_097_));
 sky130_fd_sc_hd__mux2_1 _238_ (.A0(\delay_counter[3] ),
    .A1(_096_),
    .S(_097_),
    .X(_098_));
 sky130_fd_sc_hd__a2bb2oi_1 _239_ (.A1_N(_072_),
    .A2_N(_095_),
    .B1(_098_),
    .B2(_048_),
    .Y(_099_));
 sky130_fd_sc_hd__o31ai_1 _240_ (.A1(_048_),
    .A2(_036_),
    .A3(_094_),
    .B1(_099_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_1 _241_ (.A(_054_),
    .B(_140_),
    .Y(_100_));
 sky130_fd_sc_hd__nand2b_1 _242_ (.A_N(\state[1] ),
    .B(_139_),
    .Y(_101_));
 sky130_fd_sc_hd__nand2_1 _243_ (.A(net32),
    .B(\target_status[0] ),
    .Y(_102_));
 sky130_fd_sc_hd__o21ai_0 _244_ (.A1(_101_),
    .A2(_102_),
    .B1(net16),
    .Y(_103_));
 sky130_fd_sc_hd__nor2b_1 _245_ (.A(\target_status[0] ),
    .B_N(net32),
    .Y(_104_));
 sky130_fd_sc_hd__nor2_1 _246_ (.A(net16),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__a21oi_1 _247_ (.A1(_048_),
    .A2(_103_),
    .B1(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__o22a_1 _248_ (.A1(net16),
    .A2(_100_),
    .B1(_106_),
    .B2(net6),
    .X(_016_));
 sky130_fd_sc_hd__nand2_1 _249_ (.A(net33),
    .B(\target_status[1] ),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _250_ (.A1(_101_),
    .A2(_107_),
    .B1(net17),
    .Y(_108_));
 sky130_fd_sc_hd__nor2b_1 _251_ (.A(\target_status[1] ),
    .B_N(net33),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _252_ (.A(net17),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__a21oi_1 _253_ (.A1(_048_),
    .A2(_108_),
    .B1(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__o22a_1 _254_ (.A1(net17),
    .A2(_100_),
    .B1(_111_),
    .B2(net7),
    .X(_017_));
 sky130_fd_sc_hd__nand2_1 _255_ (.A(net34),
    .B(\target_status[2] ),
    .Y(_112_));
 sky130_fd_sc_hd__o21ai_0 _256_ (.A1(_101_),
    .A2(_112_),
    .B1(net18),
    .Y(_113_));
 sky130_fd_sc_hd__nor2b_1 _257_ (.A(\target_status[2] ),
    .B_N(net34),
    .Y(_114_));
 sky130_fd_sc_hd__nor2_1 _258_ (.A(net18),
    .B(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__a21oi_1 _259_ (.A1(_048_),
    .A2(_113_),
    .B1(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__o22a_1 _260_ (.A1(net18),
    .A2(_100_),
    .B1(_116_),
    .B2(net8),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _261_ (.A(net35),
    .B(\target_status[3] ),
    .Y(_117_));
 sky130_fd_sc_hd__o21ai_0 _262_ (.A1(_101_),
    .A2(_117_),
    .B1(net19),
    .Y(_118_));
 sky130_fd_sc_hd__nor2b_1 _263_ (.A(\target_status[3] ),
    .B_N(net35),
    .Y(_119_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(net19),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__a21oi_1 _265_ (.A1(_048_),
    .A2(_118_),
    .B1(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__o22a_1 _266_ (.A1(net19),
    .A2(_100_),
    .B1(_121_),
    .B2(net9),
    .X(_019_));
 sky130_fd_sc_hd__and3b_1 _267_ (.A_N(\state[2] ),
    .B(\state[1] ),
    .C(_139_),
    .X(_122_));
 sky130_fd_sc_hd__and2_1 _268_ (.A(_050_),
    .B(_122_),
    .X(_123_));
 sky130_fd_sc_hd__a21oi_1 _269_ (.A1(net32),
    .A2(_123_),
    .B1(net24),
    .Y(_124_));
 sky130_fd_sc_hd__a21oi_1 _270_ (.A1(_104_),
    .A2(_122_),
    .B1(_124_),
    .Y(_020_));
 sky130_fd_sc_hd__a21oi_1 _271_ (.A1(net33),
    .A2(_123_),
    .B1(net25),
    .Y(_125_));
 sky130_fd_sc_hd__a21oi_1 _272_ (.A1(_109_),
    .A2(_122_),
    .B1(_125_),
    .Y(_021_));
 sky130_fd_sc_hd__a21oi_1 _273_ (.A1(net34),
    .A2(_123_),
    .B1(net26),
    .Y(_126_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_114_),
    .A2(_122_),
    .B1(_126_),
    .Y(_022_));
 sky130_fd_sc_hd__a21oi_1 _275_ (.A1(net35),
    .A2(_123_),
    .B1(net27),
    .Y(_127_));
 sky130_fd_sc_hd__a21oi_1 _276_ (.A1(_119_),
    .A2(_122_),
    .B1(_127_),
    .Y(_023_));
 sky130_fd_sc_hd__nand3_2 _277_ (.A(_047_),
    .B(_054_),
    .C(_140_),
    .Y(_128_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(net32),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nand2b_1 _279_ (.A_N(_066_),
    .B(_072_),
    .Y(_130_));
 sky130_fd_sc_hd__buf_6 _280_ (.A(_130_),
    .X(_131_));
 sky130_fd_sc_hd__mux2i_1 _281_ (.A0(_062_),
    .A1(_129_),
    .S(_131_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _282_ (.A(net33),
    .B(_128_),
    .Y(_132_));
 sky130_fd_sc_hd__mux2i_1 _283_ (.A0(_064_),
    .A1(_132_),
    .S(_131_),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _284_ (.A(net34),
    .B(_128_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2i_1 _285_ (.A0(_063_),
    .A1(_133_),
    .S(_131_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2_1 _286_ (.A(net35),
    .B(_128_),
    .Y(_134_));
 sky130_fd_sc_hd__mux2i_1 _287_ (.A0(_061_),
    .A1(_134_),
    .S(_131_),
    .Y(_027_));
 sky130_fd_sc_hd__o211ai_1 _288_ (.A1(_047_),
    .A2(_054_),
    .B1(_140_),
    .C1(_053_),
    .Y(_135_));
 sky130_fd_sc_hd__nand2_1 _289_ (.A(_139_),
    .B(_050_),
    .Y(_136_));
 sky130_fd_sc_hd__o2111a_1 _290_ (.A1(_066_),
    .A2(_072_),
    .B1(_135_),
    .C1(_074_),
    .D1(_136_),
    .X(_028_));
 sky130_fd_sc_hd__nand3b_1 _291_ (.A_N(_048_),
    .B(_054_),
    .C(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__o21ai_0 _292_ (.A1(_054_),
    .A2(_136_),
    .B1(_137_),
    .Y(_029_));
 sky130_fd_sc_hd__or2_0 _293_ (.A(_059_),
    .B(_123_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(net2),
    .A1(\target_status[0] ),
    .S(_131_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(net3),
    .A1(\target_status[1] ),
    .S(_131_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(net4),
    .A1(\target_status[2] ),
    .S(_131_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(net5),
    .A1(\target_status[3] ),
    .S(_131_),
    .X(_034_));
 sky130_fd_sc_hd__o21bai_1 _298_ (.A1(_139_),
    .A2(_059_),
    .B1_N(net36),
    .Y(_138_));
 sky130_fd_sc_hd__o311a_1 _299_ (.A1(_047_),
    .A2(_055_),
    .A3(net36),
    .B1(_131_),
    .C1(_138_),
    .X(_035_));
 sky130_fd_sc_hd__ha_1 _300_ (.A(_146_),
    .B(_147_),
    .COUT(_148_),
    .SUM(_149_));
 sky130_fd_sc_hd__ha_1 _301_ (.A(_146_),
    .B(_147_),
    .COUT(_150_),
    .SUM(_151_));
 sky130_fd_sc_hd__dfrtp_1 _302_ (.D(_000_),
    .Q(net31),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _303_ (.D(_001_),
    .Q(net30),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _304_ (.D(_002_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _305_ (.D(_003_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _306_ (.D(_004_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _307_ (.D(_005_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _308_ (.D(_006_),
    .Q(net13),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _309_ (.D(_007_),
    .Q(net12),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _310_ (.D(_008_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _311_ (.D(_009_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _312_ (.D(_010_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 _313_ (.D(_011_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_counter[0]$_DFFE_PN0P_  (.D(_012_),
    .Q(\delay_counter[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_counter[1]$_DFFE_PN0P_  (.D(_013_),
    .Q(\delay_counter[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_counter[2]$_DFFE_PN0P_  (.D(_014_),
    .Q(\delay_counter[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \delay_counter[3]$_DFFE_PN0P_  (.D(_015_),
    .Q(\delay_counter[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \domain_isolation_on[0]$_DFFE_PN1P_  (.D(_016_),
    .Q(net16),
    .SET_B(net10),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \domain_isolation_on[1]$_DFFE_PN1P_  (.D(_017_),
    .Q(net17),
    .SET_B(net10),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \domain_isolation_on[2]$_DFFE_PN1P_  (.D(_018_),
    .Q(net18),
    .SET_B(net10),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \domain_isolation_on[3]$_DFFE_PN1P_  (.D(_019_),
    .Q(net19),
    .SET_B(net10),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \domain_reset_n[0]$_DFFE_PN0P_  (.D(_020_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \domain_reset_n[1]$_DFFE_PN0P_  (.D(_021_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \domain_reset_n[2]$_DFFE_PN0P_  (.D(_022_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \domain_reset_n[3]$_DFFE_PN0P_  (.D(_023_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \domain_transition[0]$_DFFE_PN0P_  (.D(_024_),
    .Q(net32),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \domain_transition[1]$_DFFE_PN0P_  (.D(_025_),
    .Q(net33),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \domain_transition[2]$_DFFE_PN0P_  (.D(_026_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \domain_transition[3]$_DFFE_PN0P_  (.D(_027_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFFE_PN0P_  (.D(_028_),
    .Q(\state[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \state[1]$_DFFE_PN0P_  (.D(_029_),
    .Q(\state[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \state[2]$_DFFE_PN0P_  (.D(_030_),
    .Q(\state[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \target_status[0]$_DFFE_PN0P_  (.D(_031_),
    .Q(\target_status[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \target_status[1]$_DFFE_PN0P_  (.D(_032_),
    .Q(\target_status[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \target_status[2]$_DFFE_PN0P_  (.D(_033_),
    .Q(\target_status[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \target_status[3]$_DFFE_PN0P_  (.D(_034_),
    .Q(\target_status[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \transition_done$_DFFE_PN1P_  (.D(_035_),
    .Q(net36),
    .SET_B(net10),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net10),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_45 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(domain_enable[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(domain_enable[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(domain_enable[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(domain_enable[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(domain_isolate[0]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(domain_isolate[1]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(domain_isolate[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(domain_isolate[3]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input9 (.A(net37),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(start_transition),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net12),
    .X(domain_clock_on[0]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(domain_clock_on[1]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(domain_clock_on[2]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(domain_clock_on[3]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(domain_isolation_on[0]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(domain_isolation_on[1]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(domain_isolation_on[2]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(domain_isolation_on[3]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(domain_power_on[0]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(domain_power_on[1]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(domain_power_on[2]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(domain_power_on[3]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(domain_reset_n[0]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(domain_reset_n[1]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(domain_reset_n[2]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(domain_reset_n[3]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(domain_status[0]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(domain_status[1]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(domain_status[2]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(domain_status[3]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(domain_transition[0]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(domain_transition[1]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(domain_transition[2]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(domain_transition[3]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(transition_done));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net37));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_125 ();
endmodule
