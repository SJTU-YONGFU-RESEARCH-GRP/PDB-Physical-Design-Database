module credit_based_fifo (clk,
    credit_return,
    empty,
    full,
    ready_in,
    ready_out,
    rst_n,
    valid_in,
    valid_out,
    credits_available,
    data_in,
    data_out,
    fifo_level);
 input clk;
 input credit_return;
 output empty;
 output full;
 input ready_in;
 output ready_out;
 input rst_n;
 input valid_in;
 output valid_out;
 output [4:0] credits_available;
 input [7:0] data_in;
 output [7:0] data_out;
 output [4:0] fifo_level;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \read_ptr[0] ;
 wire \read_ptr[1] ;
 wire \read_ptr[2] ;
 wire \read_ptr[3] ;
 wire \read_ptr[4] ;
 wire \write_ptr[0] ;
 wire \write_ptr[1] ;
 wire \write_ptr[2] ;
 wire \write_ptr[3] ;
 wire \write_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 INV_X1 _0616_ (.A(_0615_),
    .ZN(net18));
 CLKBUF_X2 _0617_ (.A(_0588_),
    .Z(_0158_));
 INV_X1 _0618_ (.A(_0158_),
    .ZN(_0159_));
 BUF_X4 _0619_ (.A(_0591_),
    .Z(_0160_));
 XNOR2_X1 _0620_ (.A(_0583_),
    .B(_0160_),
    .ZN(net20));
 NAND4_X1 _0621_ (.A1(_0159_),
    .A2(net18),
    .A3(net19),
    .A4(net20),
    .ZN(_0161_));
 AOI21_X1 _0622_ (.A(_0590_),
    .B1(_0160_),
    .B2(_0594_),
    .ZN(_0162_));
 INV_X1 _0623_ (.A(_0582_),
    .ZN(_0163_));
 NAND3_X1 _0624_ (.A1(_0592_),
    .A2(_0163_),
    .A3(_0160_),
    .ZN(_0164_));
 AOI21_X1 _0625_ (.A(_0161_),
    .B1(_0162_),
    .B2(_0164_),
    .ZN(_0165_));
 AND4_X1 _0626_ (.A1(_0158_),
    .A2(net18),
    .A3(net19),
    .A4(net20),
    .ZN(_0166_));
 AND2_X1 _0627_ (.A1(_0164_),
    .A2(_0162_),
    .ZN(_0167_));
 BUF_X4 _0628_ (.A(\write_ptr[4] ),
    .Z(_0168_));
 XOR2_X2 _0629_ (.A(_0168_),
    .B(\read_ptr[4] ),
    .Z(_0169_));
 OR2_X1 _0630_ (.A1(_0587_),
    .A2(_0590_),
    .ZN(_0170_));
 INV_X1 _0631_ (.A(_0583_),
    .ZN(_0171_));
 AOI21_X1 _0632_ (.A(_0170_),
    .B1(_0160_),
    .B2(_0171_),
    .ZN(_0172_));
 NOR2_X1 _0633_ (.A1(_0158_),
    .A2(_0587_),
    .ZN(_0173_));
 OAI21_X1 _0634_ (.A(_0169_),
    .B1(_0172_),
    .B2(_0173_),
    .ZN(_0174_));
 OR3_X1 _0635_ (.A1(_0169_),
    .A2(_0172_),
    .A3(_0173_),
    .ZN(_0175_));
 AOI221_X2 _0636_ (.A(_0165_),
    .B1(_0166_),
    .B2(_0167_),
    .C1(_0174_),
    .C2(_0175_),
    .ZN(_0176_));
 BUF_X4 _0637_ (.A(_0176_),
    .Z(_0177_));
 INV_X1 _0638_ (.A(_0177_),
    .ZN(net23));
 INV_X1 _0639_ (.A(net8),
    .ZN(_0178_));
 INV_X1 _0640_ (.A(_0000_),
    .ZN(_0179_));
 NOR4_X4 _0641_ (.A1(net7),
    .A2(net6),
    .A3(net5),
    .A4(_0179_),
    .ZN(_0180_));
 NAND2_X1 _0642_ (.A1(_0178_),
    .A2(_0180_),
    .ZN(_0181_));
 BUF_X2 _0643_ (.A(_0181_),
    .Z(_0182_));
 NAND2_X1 _0644_ (.A1(net3),
    .A2(_0182_),
    .ZN(_0183_));
 NOR2_X2 _0645_ (.A1(net23),
    .A2(_0183_),
    .ZN(_0595_));
 INV_X1 _0646_ (.A(_0595_),
    .ZN(_0598_));
 XNOR2_X2 _0647_ (.A(_0168_),
    .B(\read_ptr[4] ),
    .ZN(_0184_));
 AND4_X1 _0648_ (.A1(_0592_),
    .A2(_0158_),
    .A3(_0615_),
    .A4(_0160_),
    .ZN(_0185_));
 AND2_X1 _0649_ (.A1(_0184_),
    .A2(_0185_),
    .ZN(net17));
 INV_X1 _0650_ (.A(net1),
    .ZN(_0596_));
 BUF_X2 _0651_ (.A(rst_n),
    .Z(_0186_));
 INV_X1 _0652_ (.A(net2),
    .ZN(_0187_));
 AOI22_X4 _0653_ (.A1(net25),
    .A2(_0187_),
    .B1(_0184_),
    .B2(_0185_),
    .ZN(_0188_));
 NAND2_X4 _0654_ (.A1(_0186_),
    .A2(_0188_),
    .ZN(_0189_));
 CLKBUF_X2 _0655_ (.A(\read_ptr[1] ),
    .Z(_0190_));
 BUF_X4 _0656_ (.A(_0190_),
    .Z(_0191_));
 BUF_X4 _0657_ (.A(_0191_),
    .Z(_0192_));
 MUX2_X1 _0658_ (.A(\mem[0][0] ),
    .B(\mem[2][0] ),
    .S(_0192_),
    .Z(_0193_));
 MUX2_X1 _0659_ (.A(\mem[1][0] ),
    .B(\mem[3][0] ),
    .S(_0192_),
    .Z(_0194_));
 CLKBUF_X3 _0660_ (.A(\read_ptr[0] ),
    .Z(_0195_));
 BUF_X4 _0661_ (.A(_0195_),
    .Z(_0196_));
 MUX2_X1 _0662_ (.A(_0193_),
    .B(_0194_),
    .S(_0196_),
    .Z(_0197_));
 MUX2_X1 _0663_ (.A(\mem[8][0] ),
    .B(\mem[10][0] ),
    .S(_0192_),
    .Z(_0198_));
 MUX2_X1 _0664_ (.A(\mem[9][0] ),
    .B(\mem[11][0] ),
    .S(_0192_),
    .Z(_0199_));
 MUX2_X1 _0665_ (.A(_0198_),
    .B(_0199_),
    .S(_0196_),
    .Z(_0200_));
 CLKBUF_X3 _0666_ (.A(\read_ptr[3] ),
    .Z(_0201_));
 CLKBUF_X3 _0667_ (.A(_0201_),
    .Z(_0202_));
 MUX2_X1 _0668_ (.A(_0197_),
    .B(_0200_),
    .S(_0202_),
    .Z(_0203_));
 BUF_X2 _0669_ (.A(\read_ptr[2] ),
    .Z(_0204_));
 NOR2_X4 _0670_ (.A1(_0204_),
    .A2(_0189_),
    .ZN(_0205_));
 INV_X1 _0671_ (.A(_0204_),
    .ZN(_0206_));
 NOR2_X4 _0672_ (.A1(_0206_),
    .A2(_0189_),
    .ZN(_0207_));
 MUX2_X1 _0673_ (.A(\mem[4][0] ),
    .B(\mem[6][0] ),
    .S(_0191_),
    .Z(_0208_));
 MUX2_X1 _0674_ (.A(\mem[5][0] ),
    .B(\mem[7][0] ),
    .S(_0191_),
    .Z(_0209_));
 MUX2_X1 _0675_ (.A(_0208_),
    .B(_0209_),
    .S(_0195_),
    .Z(_0210_));
 MUX2_X1 _0676_ (.A(\mem[12][0] ),
    .B(\mem[14][0] ),
    .S(_0191_),
    .Z(_0211_));
 MUX2_X1 _0677_ (.A(\mem[13][0] ),
    .B(\mem[15][0] ),
    .S(_0191_),
    .Z(_0212_));
 MUX2_X1 _0678_ (.A(_0211_),
    .B(_0212_),
    .S(_0195_),
    .Z(_0213_));
 MUX2_X1 _0679_ (.A(_0210_),
    .B(_0213_),
    .S(_0201_),
    .Z(_0214_));
 AOI222_X2 _0680_ (.A1(net9),
    .A2(_0189_),
    .B1(_0203_),
    .B2(_0205_),
    .C1(_0207_),
    .C2(_0214_),
    .ZN(_0215_));
 INV_X1 _0681_ (.A(_0215_),
    .ZN(_0011_));
 CLKBUF_X3 _0682_ (.A(_0191_),
    .Z(_0216_));
 MUX2_X1 _0683_ (.A(\mem[4][1] ),
    .B(\mem[6][1] ),
    .S(_0216_),
    .Z(_0217_));
 MUX2_X1 _0684_ (.A(\mem[5][1] ),
    .B(\mem[7][1] ),
    .S(_0216_),
    .Z(_0218_));
 BUF_X4 _0685_ (.A(_0195_),
    .Z(_0219_));
 MUX2_X1 _0686_ (.A(_0217_),
    .B(_0218_),
    .S(_0219_),
    .Z(_0220_));
 BUF_X4 _0687_ (.A(_0191_),
    .Z(_0221_));
 MUX2_X1 _0688_ (.A(\mem[12][1] ),
    .B(\mem[14][1] ),
    .S(_0221_),
    .Z(_0222_));
 MUX2_X1 _0689_ (.A(\mem[13][1] ),
    .B(\mem[15][1] ),
    .S(_0192_),
    .Z(_0223_));
 MUX2_X1 _0690_ (.A(_0222_),
    .B(_0223_),
    .S(_0196_),
    .Z(_0224_));
 MUX2_X1 _0691_ (.A(_0220_),
    .B(_0224_),
    .S(_0202_),
    .Z(_0225_));
 BUF_X4 _0692_ (.A(_0190_),
    .Z(_0226_));
 MUX2_X1 _0693_ (.A(\mem[0][1] ),
    .B(\mem[2][1] ),
    .S(_0226_),
    .Z(_0227_));
 BUF_X4 _0694_ (.A(_0190_),
    .Z(_0228_));
 MUX2_X1 _0695_ (.A(\mem[1][1] ),
    .B(\mem[3][1] ),
    .S(_0228_),
    .Z(_0229_));
 BUF_X4 _0696_ (.A(_0195_),
    .Z(_0230_));
 MUX2_X1 _0697_ (.A(_0227_),
    .B(_0229_),
    .S(_0230_),
    .Z(_0231_));
 MUX2_X1 _0698_ (.A(\mem[8][1] ),
    .B(\mem[10][1] ),
    .S(_0228_),
    .Z(_0232_));
 CLKBUF_X3 _0699_ (.A(_0191_),
    .Z(_0233_));
 MUX2_X1 _0700_ (.A(\mem[9][1] ),
    .B(\mem[11][1] ),
    .S(_0233_),
    .Z(_0234_));
 MUX2_X1 _0701_ (.A(_0232_),
    .B(_0234_),
    .S(_0219_),
    .Z(_0235_));
 MUX2_X1 _0702_ (.A(_0231_),
    .B(_0235_),
    .S(_0201_),
    .Z(_0236_));
 AOI222_X2 _0703_ (.A1(net10),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0225_),
    .C1(_0236_),
    .C2(_0205_),
    .ZN(_0237_));
 INV_X1 _0704_ (.A(_0237_),
    .ZN(_0012_));
 MUX2_X1 _0705_ (.A(\mem[4][2] ),
    .B(\mem[6][2] ),
    .S(_0216_),
    .Z(_0238_));
 MUX2_X1 _0706_ (.A(\mem[5][2] ),
    .B(\mem[7][2] ),
    .S(_0216_),
    .Z(_0239_));
 MUX2_X1 _0707_ (.A(_0238_),
    .B(_0239_),
    .S(_0219_),
    .Z(_0240_));
 MUX2_X1 _0708_ (.A(\mem[12][2] ),
    .B(\mem[14][2] ),
    .S(_0221_),
    .Z(_0241_));
 MUX2_X1 _0709_ (.A(\mem[13][2] ),
    .B(\mem[15][2] ),
    .S(_0192_),
    .Z(_0242_));
 MUX2_X1 _0710_ (.A(_0241_),
    .B(_0242_),
    .S(_0196_),
    .Z(_0243_));
 MUX2_X1 _0711_ (.A(_0240_),
    .B(_0243_),
    .S(_0202_),
    .Z(_0244_));
 MUX2_X1 _0712_ (.A(\mem[0][2] ),
    .B(\mem[2][2] ),
    .S(_0226_),
    .Z(_0245_));
 MUX2_X1 _0713_ (.A(\mem[1][2] ),
    .B(\mem[3][2] ),
    .S(_0228_),
    .Z(_0246_));
 MUX2_X1 _0714_ (.A(_0245_),
    .B(_0246_),
    .S(_0230_),
    .Z(_0247_));
 MUX2_X1 _0715_ (.A(\mem[8][2] ),
    .B(\mem[10][2] ),
    .S(_0228_),
    .Z(_0248_));
 MUX2_X1 _0716_ (.A(\mem[9][2] ),
    .B(\mem[11][2] ),
    .S(_0233_),
    .Z(_0249_));
 MUX2_X1 _0717_ (.A(_0248_),
    .B(_0249_),
    .S(_0219_),
    .Z(_0250_));
 MUX2_X1 _0718_ (.A(_0247_),
    .B(_0250_),
    .S(_0201_),
    .Z(_0251_));
 AOI222_X2 _0719_ (.A1(net11),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0244_),
    .C1(_0251_),
    .C2(_0205_),
    .ZN(_0252_));
 INV_X1 _0720_ (.A(_0252_),
    .ZN(_0013_));
 MUX2_X1 _0721_ (.A(\mem[4][3] ),
    .B(\mem[6][3] ),
    .S(_0216_),
    .Z(_0253_));
 MUX2_X1 _0722_ (.A(\mem[5][3] ),
    .B(\mem[7][3] ),
    .S(_0216_),
    .Z(_0254_));
 MUX2_X1 _0723_ (.A(_0253_),
    .B(_0254_),
    .S(_0219_),
    .Z(_0255_));
 MUX2_X1 _0724_ (.A(\mem[12][3] ),
    .B(\mem[14][3] ),
    .S(_0221_),
    .Z(_0256_));
 MUX2_X1 _0725_ (.A(\mem[13][3] ),
    .B(\mem[15][3] ),
    .S(_0192_),
    .Z(_0257_));
 MUX2_X1 _0726_ (.A(_0256_),
    .B(_0257_),
    .S(_0196_),
    .Z(_0258_));
 MUX2_X1 _0727_ (.A(_0255_),
    .B(_0258_),
    .S(_0202_),
    .Z(_0259_));
 MUX2_X1 _0728_ (.A(\mem[0][3] ),
    .B(\mem[2][3] ),
    .S(_0226_),
    .Z(_0260_));
 MUX2_X1 _0729_ (.A(\mem[1][3] ),
    .B(\mem[3][3] ),
    .S(_0226_),
    .Z(_0261_));
 MUX2_X1 _0730_ (.A(_0260_),
    .B(_0261_),
    .S(_0230_),
    .Z(_0262_));
 MUX2_X1 _0731_ (.A(\mem[8][3] ),
    .B(\mem[10][3] ),
    .S(_0228_),
    .Z(_0263_));
 MUX2_X1 _0732_ (.A(\mem[9][3] ),
    .B(\mem[11][3] ),
    .S(_0233_),
    .Z(_0264_));
 MUX2_X1 _0733_ (.A(_0263_),
    .B(_0264_),
    .S(_0230_),
    .Z(_0265_));
 MUX2_X1 _0734_ (.A(_0262_),
    .B(_0265_),
    .S(_0201_),
    .Z(_0266_));
 AOI222_X2 _0735_ (.A1(net12),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0259_),
    .C1(_0266_),
    .C2(_0205_),
    .ZN(_0267_));
 INV_X1 _0736_ (.A(_0267_),
    .ZN(_0014_));
 MUX2_X1 _0737_ (.A(\mem[4][4] ),
    .B(\mem[6][4] ),
    .S(_0233_),
    .Z(_0268_));
 MUX2_X1 _0738_ (.A(\mem[5][4] ),
    .B(\mem[7][4] ),
    .S(_0216_),
    .Z(_0269_));
 MUX2_X1 _0739_ (.A(_0268_),
    .B(_0269_),
    .S(_0219_),
    .Z(_0270_));
 MUX2_X1 _0740_ (.A(\mem[12][4] ),
    .B(\mem[14][4] ),
    .S(_0221_),
    .Z(_0271_));
 MUX2_X1 _0741_ (.A(\mem[13][4] ),
    .B(\mem[15][4] ),
    .S(_0192_),
    .Z(_0272_));
 MUX2_X1 _0742_ (.A(_0271_),
    .B(_0272_),
    .S(_0196_),
    .Z(_0273_));
 MUX2_X1 _0743_ (.A(_0270_),
    .B(_0273_),
    .S(_0202_),
    .Z(_0274_));
 MUX2_X1 _0744_ (.A(\mem[0][4] ),
    .B(\mem[2][4] ),
    .S(_0226_),
    .Z(_0275_));
 MUX2_X1 _0745_ (.A(\mem[1][4] ),
    .B(\mem[3][4] ),
    .S(_0226_),
    .Z(_0276_));
 MUX2_X1 _0746_ (.A(_0275_),
    .B(_0276_),
    .S(_0230_),
    .Z(_0277_));
 MUX2_X1 _0747_ (.A(\mem[8][4] ),
    .B(\mem[10][4] ),
    .S(_0228_),
    .Z(_0278_));
 MUX2_X1 _0748_ (.A(\mem[9][4] ),
    .B(\mem[11][4] ),
    .S(_0233_),
    .Z(_0279_));
 MUX2_X1 _0749_ (.A(_0278_),
    .B(_0279_),
    .S(_0230_),
    .Z(_0280_));
 MUX2_X1 _0750_ (.A(_0277_),
    .B(_0280_),
    .S(_0201_),
    .Z(_0281_));
 AOI222_X2 _0751_ (.A1(net13),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0274_),
    .C1(_0281_),
    .C2(_0205_),
    .ZN(_0282_));
 INV_X1 _0752_ (.A(_0282_),
    .ZN(_0015_));
 MUX2_X1 _0753_ (.A(\mem[4][5] ),
    .B(\mem[6][5] ),
    .S(_0233_),
    .Z(_0283_));
 MUX2_X1 _0754_ (.A(\mem[5][5] ),
    .B(\mem[7][5] ),
    .S(_0216_),
    .Z(_0284_));
 MUX2_X1 _0755_ (.A(_0283_),
    .B(_0284_),
    .S(_0219_),
    .Z(_0285_));
 MUX2_X1 _0756_ (.A(\mem[12][5] ),
    .B(\mem[14][5] ),
    .S(_0221_),
    .Z(_0286_));
 MUX2_X1 _0757_ (.A(\mem[13][5] ),
    .B(\mem[15][5] ),
    .S(_0221_),
    .Z(_0287_));
 MUX2_X1 _0758_ (.A(_0286_),
    .B(_0287_),
    .S(_0196_),
    .Z(_0288_));
 MUX2_X1 _0759_ (.A(_0285_),
    .B(_0288_),
    .S(_0202_),
    .Z(_0289_));
 MUX2_X1 _0760_ (.A(\mem[0][5] ),
    .B(\mem[2][5] ),
    .S(_0226_),
    .Z(_0290_));
 MUX2_X1 _0761_ (.A(\mem[1][5] ),
    .B(\mem[3][5] ),
    .S(_0226_),
    .Z(_0291_));
 MUX2_X1 _0762_ (.A(_0290_),
    .B(_0291_),
    .S(_0230_),
    .Z(_0292_));
 MUX2_X1 _0763_ (.A(\mem[8][5] ),
    .B(\mem[10][5] ),
    .S(_0228_),
    .Z(_0293_));
 MUX2_X1 _0764_ (.A(\mem[9][5] ),
    .B(\mem[11][5] ),
    .S(_0233_),
    .Z(_0294_));
 MUX2_X1 _0765_ (.A(_0293_),
    .B(_0294_),
    .S(_0230_),
    .Z(_0295_));
 MUX2_X1 _0766_ (.A(_0292_),
    .B(_0295_),
    .S(_0201_),
    .Z(_0296_));
 AOI222_X2 _0767_ (.A1(net14),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0289_),
    .C1(_0296_),
    .C2(_0205_),
    .ZN(_0297_));
 INV_X1 _0768_ (.A(_0297_),
    .ZN(_0016_));
 MUX2_X1 _0769_ (.A(\mem[4][6] ),
    .B(\mem[6][6] ),
    .S(_0233_),
    .Z(_0298_));
 MUX2_X1 _0770_ (.A(\mem[5][6] ),
    .B(\mem[7][6] ),
    .S(_0216_),
    .Z(_0299_));
 MUX2_X1 _0771_ (.A(_0298_),
    .B(_0299_),
    .S(_0219_),
    .Z(_0300_));
 MUX2_X1 _0772_ (.A(\mem[12][6] ),
    .B(\mem[14][6] ),
    .S(_0221_),
    .Z(_0301_));
 MUX2_X1 _0773_ (.A(\mem[13][6] ),
    .B(\mem[15][6] ),
    .S(_0221_),
    .Z(_0302_));
 MUX2_X1 _0774_ (.A(_0301_),
    .B(_0302_),
    .S(_0196_),
    .Z(_0303_));
 MUX2_X1 _0775_ (.A(_0300_),
    .B(_0303_),
    .S(_0202_),
    .Z(_0304_));
 MUX2_X1 _0776_ (.A(\mem[0][6] ),
    .B(\mem[2][6] ),
    .S(_0191_),
    .Z(_0305_));
 MUX2_X1 _0777_ (.A(\mem[1][6] ),
    .B(\mem[3][6] ),
    .S(_0226_),
    .Z(_0306_));
 MUX2_X1 _0778_ (.A(_0305_),
    .B(_0306_),
    .S(_0195_),
    .Z(_0307_));
 MUX2_X1 _0779_ (.A(\mem[8][6] ),
    .B(\mem[10][6] ),
    .S(_0228_),
    .Z(_0308_));
 MUX2_X1 _0780_ (.A(\mem[9][6] ),
    .B(\mem[11][6] ),
    .S(_0233_),
    .Z(_0309_));
 MUX2_X1 _0781_ (.A(_0308_),
    .B(_0309_),
    .S(_0230_),
    .Z(_0310_));
 MUX2_X1 _0782_ (.A(_0307_),
    .B(_0310_),
    .S(_0201_),
    .Z(_0311_));
 AOI222_X2 _0783_ (.A1(net15),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0304_),
    .C1(_0311_),
    .C2(_0205_),
    .ZN(_0312_));
 INV_X1 _0784_ (.A(_0312_),
    .ZN(_0017_));
 MUX2_X1 _0785_ (.A(\mem[4][7] ),
    .B(\mem[6][7] ),
    .S(_0233_),
    .Z(_0313_));
 MUX2_X1 _0786_ (.A(\mem[5][7] ),
    .B(\mem[7][7] ),
    .S(_0216_),
    .Z(_0314_));
 MUX2_X1 _0787_ (.A(_0313_),
    .B(_0314_),
    .S(_0219_),
    .Z(_0315_));
 MUX2_X1 _0788_ (.A(\mem[12][7] ),
    .B(\mem[14][7] ),
    .S(_0221_),
    .Z(_0316_));
 MUX2_X1 _0789_ (.A(\mem[13][7] ),
    .B(\mem[15][7] ),
    .S(_0221_),
    .Z(_0317_));
 MUX2_X1 _0790_ (.A(_0316_),
    .B(_0317_),
    .S(_0219_),
    .Z(_0318_));
 MUX2_X1 _0791_ (.A(_0315_),
    .B(_0318_),
    .S(_0202_),
    .Z(_0319_));
 MUX2_X1 _0792_ (.A(\mem[0][7] ),
    .B(\mem[2][7] ),
    .S(_0191_),
    .Z(_0320_));
 MUX2_X1 _0793_ (.A(\mem[1][7] ),
    .B(\mem[3][7] ),
    .S(_0226_),
    .Z(_0321_));
 MUX2_X1 _0794_ (.A(_0320_),
    .B(_0321_),
    .S(_0195_),
    .Z(_0322_));
 MUX2_X1 _0795_ (.A(\mem[8][7] ),
    .B(\mem[10][7] ),
    .S(_0228_),
    .Z(_0323_));
 MUX2_X1 _0796_ (.A(\mem[9][7] ),
    .B(\mem[11][7] ),
    .S(_0228_),
    .Z(_0324_));
 MUX2_X1 _0797_ (.A(_0323_),
    .B(_0324_),
    .S(_0230_),
    .Z(_0325_));
 MUX2_X1 _0798_ (.A(_0322_),
    .B(_0325_),
    .S(_0201_),
    .Z(_0326_));
 AOI222_X2 _0799_ (.A1(net16),
    .A2(_0189_),
    .B1(_0207_),
    .B2(_0319_),
    .C1(_0326_),
    .C2(_0205_),
    .ZN(_0327_));
 INV_X1 _0800_ (.A(_0327_),
    .ZN(_0018_));
 CLKBUF_X2 _0801_ (.A(data_in[0]),
    .Z(_0328_));
 BUF_X2 _0802_ (.A(_0328_),
    .Z(_0329_));
 INV_X2 _0803_ (.A(_0186_),
    .ZN(_0330_));
 BUF_X1 _0804_ (.A(\write_ptr[2] ),
    .Z(_0331_));
 BUF_X1 _0805_ (.A(\write_ptr[3] ),
    .Z(_0332_));
 NOR3_X1 _0806_ (.A1(_0330_),
    .A2(_0331_),
    .A3(_0332_),
    .ZN(_0333_));
 AND2_X1 _0807_ (.A1(net3),
    .A2(_0602_),
    .ZN(_0334_));
 AND4_X1 _0808_ (.A1(_0177_),
    .A2(_0182_),
    .A3(_0333_),
    .A4(_0334_),
    .ZN(_0335_));
 BUF_X4 _0809_ (.A(_0335_),
    .Z(_0336_));
 MUX2_X1 _0810_ (.A(\mem[0][0] ),
    .B(_0329_),
    .S(_0336_),
    .Z(_0019_));
 CLKBUF_X2 _0811_ (.A(data_in[1]),
    .Z(_0337_));
 CLKBUF_X2 _0812_ (.A(_0337_),
    .Z(_0338_));
 MUX2_X1 _0813_ (.A(\mem[0][1] ),
    .B(_0338_),
    .S(_0336_),
    .Z(_0020_));
 CLKBUF_X2 _0814_ (.A(data_in[2]),
    .Z(_0339_));
 BUF_X2 _0815_ (.A(_0339_),
    .Z(_0340_));
 MUX2_X1 _0816_ (.A(\mem[0][2] ),
    .B(_0340_),
    .S(_0336_),
    .Z(_0021_));
 BUF_X1 _0817_ (.A(data_in[3]),
    .Z(_0341_));
 BUF_X2 _0818_ (.A(_0341_),
    .Z(_0342_));
 MUX2_X1 _0819_ (.A(\mem[0][3] ),
    .B(_0342_),
    .S(_0336_),
    .Z(_0022_));
 BUF_X1 _0820_ (.A(data_in[4]),
    .Z(_0343_));
 BUF_X2 _0821_ (.A(_0343_),
    .Z(_0344_));
 MUX2_X1 _0822_ (.A(\mem[0][4] ),
    .B(_0344_),
    .S(_0336_),
    .Z(_0023_));
 BUF_X1 _0823_ (.A(data_in[5]),
    .Z(_0345_));
 BUF_X2 _0824_ (.A(_0345_),
    .Z(_0346_));
 MUX2_X1 _0825_ (.A(\mem[0][5] ),
    .B(_0346_),
    .S(_0336_),
    .Z(_0024_));
 BUF_X1 _0826_ (.A(data_in[6]),
    .Z(_0347_));
 BUF_X2 _0827_ (.A(_0347_),
    .Z(_0348_));
 MUX2_X1 _0828_ (.A(\mem[0][6] ),
    .B(_0348_),
    .S(_0336_),
    .Z(_0025_));
 BUF_X1 _0829_ (.A(data_in[7]),
    .Z(_0349_));
 BUF_X2 _0830_ (.A(_0349_),
    .Z(_0350_));
 MUX2_X1 _0831_ (.A(\mem[0][7] ),
    .B(_0350_),
    .S(_0336_),
    .Z(_0026_));
 NOR2_X1 _0832_ (.A1(_0330_),
    .A2(_0331_),
    .ZN(_0351_));
 AND2_X1 _0833_ (.A1(_0332_),
    .A2(_0351_),
    .ZN(_0352_));
 AND2_X1 _0834_ (.A1(net3),
    .A2(_0603_),
    .ZN(_0353_));
 AND4_X1 _0835_ (.A1(_0177_),
    .A2(_0182_),
    .A3(_0352_),
    .A4(_0353_),
    .ZN(_0354_));
 BUF_X4 _0836_ (.A(_0354_),
    .Z(_0355_));
 MUX2_X1 _0837_ (.A(\mem[10][0] ),
    .B(_0329_),
    .S(_0355_),
    .Z(_0027_));
 MUX2_X1 _0838_ (.A(\mem[10][1] ),
    .B(_0338_),
    .S(_0355_),
    .Z(_0028_));
 MUX2_X1 _0839_ (.A(\mem[10][2] ),
    .B(_0340_),
    .S(_0355_),
    .Z(_0029_));
 MUX2_X1 _0840_ (.A(\mem[10][3] ),
    .B(_0342_),
    .S(_0355_),
    .Z(_0030_));
 MUX2_X1 _0841_ (.A(\mem[10][4] ),
    .B(_0344_),
    .S(_0355_),
    .Z(_0031_));
 MUX2_X1 _0842_ (.A(\mem[10][5] ),
    .B(_0346_),
    .S(_0355_),
    .Z(_0032_));
 MUX2_X1 _0843_ (.A(\mem[10][6] ),
    .B(_0348_),
    .S(_0355_),
    .Z(_0033_));
 MUX2_X1 _0844_ (.A(\mem[10][7] ),
    .B(_0350_),
    .S(_0355_),
    .Z(_0034_));
 AND3_X1 _0845_ (.A1(net3),
    .A2(_0607_),
    .A3(_0181_),
    .ZN(_0356_));
 AND3_X1 _0846_ (.A1(_0177_),
    .A2(_0352_),
    .A3(_0356_),
    .ZN(_0357_));
 BUF_X4 _0847_ (.A(_0357_),
    .Z(_0358_));
 MUX2_X1 _0848_ (.A(\mem[11][0] ),
    .B(_0329_),
    .S(_0358_),
    .Z(_0035_));
 MUX2_X1 _0849_ (.A(\mem[11][1] ),
    .B(_0338_),
    .S(_0358_),
    .Z(_0036_));
 MUX2_X1 _0850_ (.A(\mem[11][2] ),
    .B(_0340_),
    .S(_0358_),
    .Z(_0037_));
 MUX2_X1 _0851_ (.A(\mem[11][3] ),
    .B(_0342_),
    .S(_0358_),
    .Z(_0038_));
 MUX2_X1 _0852_ (.A(\mem[11][4] ),
    .B(_0344_),
    .S(_0358_),
    .Z(_0039_));
 MUX2_X1 _0853_ (.A(\mem[11][5] ),
    .B(_0346_),
    .S(_0358_),
    .Z(_0040_));
 MUX2_X1 _0854_ (.A(\mem[11][6] ),
    .B(_0348_),
    .S(_0358_),
    .Z(_0041_));
 MUX2_X1 _0855_ (.A(\mem[11][7] ),
    .B(_0350_),
    .S(_0358_),
    .Z(_0042_));
 BUF_X4 _0856_ (.A(_0176_),
    .Z(_0359_));
 AND2_X1 _0857_ (.A1(_0186_),
    .A2(_0331_),
    .ZN(_0360_));
 AND2_X1 _0858_ (.A1(_0332_),
    .A2(_0360_),
    .ZN(_0361_));
 AND4_X1 _0859_ (.A1(_0359_),
    .A2(_0182_),
    .A3(_0334_),
    .A4(_0361_),
    .ZN(_0362_));
 BUF_X8 _0860_ (.A(_0362_),
    .Z(_0363_));
 MUX2_X1 _0861_ (.A(\mem[12][0] ),
    .B(_0329_),
    .S(_0363_),
    .Z(_0043_));
 MUX2_X1 _0862_ (.A(\mem[12][1] ),
    .B(_0338_),
    .S(_0363_),
    .Z(_0044_));
 MUX2_X1 _0863_ (.A(\mem[12][2] ),
    .B(_0340_),
    .S(_0363_),
    .Z(_0045_));
 MUX2_X1 _0864_ (.A(\mem[12][3] ),
    .B(_0342_),
    .S(_0363_),
    .Z(_0046_));
 MUX2_X1 _0865_ (.A(\mem[12][4] ),
    .B(_0344_),
    .S(_0363_),
    .Z(_0047_));
 MUX2_X1 _0866_ (.A(\mem[12][5] ),
    .B(_0346_),
    .S(_0363_),
    .Z(_0048_));
 MUX2_X1 _0867_ (.A(\mem[12][6] ),
    .B(_0348_),
    .S(_0363_),
    .Z(_0049_));
 MUX2_X1 _0868_ (.A(\mem[12][7] ),
    .B(_0350_),
    .S(_0363_),
    .Z(_0050_));
 AND2_X1 _0869_ (.A1(net3),
    .A2(_0605_),
    .ZN(_0364_));
 AND4_X1 _0870_ (.A1(_0359_),
    .A2(_0182_),
    .A3(_0361_),
    .A4(_0364_),
    .ZN(_0365_));
 BUF_X8 _0871_ (.A(_0365_),
    .Z(_0366_));
 MUX2_X1 _0872_ (.A(\mem[13][0] ),
    .B(_0329_),
    .S(_0366_),
    .Z(_0051_));
 MUX2_X1 _0873_ (.A(\mem[13][1] ),
    .B(_0338_),
    .S(_0366_),
    .Z(_0052_));
 MUX2_X1 _0874_ (.A(\mem[13][2] ),
    .B(_0340_),
    .S(_0366_),
    .Z(_0053_));
 MUX2_X1 _0875_ (.A(\mem[13][3] ),
    .B(_0342_),
    .S(_0366_),
    .Z(_0054_));
 MUX2_X1 _0876_ (.A(\mem[13][4] ),
    .B(_0344_),
    .S(_0366_),
    .Z(_0055_));
 MUX2_X1 _0877_ (.A(\mem[13][5] ),
    .B(_0346_),
    .S(_0366_),
    .Z(_0056_));
 MUX2_X1 _0878_ (.A(\mem[13][6] ),
    .B(_0348_),
    .S(_0366_),
    .Z(_0057_));
 MUX2_X1 _0879_ (.A(\mem[13][7] ),
    .B(_0350_),
    .S(_0366_),
    .Z(_0058_));
 AND4_X1 _0880_ (.A1(_0359_),
    .A2(_0182_),
    .A3(_0353_),
    .A4(_0361_),
    .ZN(_0367_));
 BUF_X8 _0881_ (.A(_0367_),
    .Z(_0368_));
 MUX2_X1 _0882_ (.A(\mem[14][0] ),
    .B(_0329_),
    .S(_0368_),
    .Z(_0059_));
 MUX2_X1 _0883_ (.A(\mem[14][1] ),
    .B(_0338_),
    .S(_0368_),
    .Z(_0060_));
 MUX2_X1 _0884_ (.A(\mem[14][2] ),
    .B(_0340_),
    .S(_0368_),
    .Z(_0061_));
 MUX2_X1 _0885_ (.A(\mem[14][3] ),
    .B(_0342_),
    .S(_0368_),
    .Z(_0062_));
 MUX2_X1 _0886_ (.A(\mem[14][4] ),
    .B(_0344_),
    .S(_0368_),
    .Z(_0063_));
 MUX2_X1 _0887_ (.A(\mem[14][5] ),
    .B(_0346_),
    .S(_0368_),
    .Z(_0064_));
 MUX2_X1 _0888_ (.A(\mem[14][6] ),
    .B(_0348_),
    .S(_0368_),
    .Z(_0065_));
 MUX2_X1 _0889_ (.A(\mem[14][7] ),
    .B(_0350_),
    .S(_0368_),
    .Z(_0066_));
 AND3_X1 _0890_ (.A1(_0177_),
    .A2(_0356_),
    .A3(_0361_),
    .ZN(_0369_));
 BUF_X4 _0891_ (.A(_0369_),
    .Z(_0370_));
 MUX2_X1 _0892_ (.A(\mem[15][0] ),
    .B(_0329_),
    .S(_0370_),
    .Z(_0067_));
 MUX2_X1 _0893_ (.A(\mem[15][1] ),
    .B(_0338_),
    .S(_0370_),
    .Z(_0068_));
 MUX2_X1 _0894_ (.A(\mem[15][2] ),
    .B(_0340_),
    .S(_0370_),
    .Z(_0069_));
 MUX2_X1 _0895_ (.A(\mem[15][3] ),
    .B(_0342_),
    .S(_0370_),
    .Z(_0070_));
 MUX2_X1 _0896_ (.A(\mem[15][4] ),
    .B(_0344_),
    .S(_0370_),
    .Z(_0071_));
 MUX2_X1 _0897_ (.A(\mem[15][5] ),
    .B(_0346_),
    .S(_0370_),
    .Z(_0072_));
 MUX2_X1 _0898_ (.A(\mem[15][6] ),
    .B(_0348_),
    .S(_0370_),
    .Z(_0073_));
 MUX2_X1 _0899_ (.A(\mem[15][7] ),
    .B(_0350_),
    .S(_0370_),
    .Z(_0074_));
 AND4_X1 _0900_ (.A1(_0359_),
    .A2(_0182_),
    .A3(_0333_),
    .A4(_0364_),
    .ZN(_0371_));
 BUF_X8 _0901_ (.A(_0371_),
    .Z(_0372_));
 MUX2_X1 _0902_ (.A(\mem[1][0] ),
    .B(_0329_),
    .S(_0372_),
    .Z(_0075_));
 MUX2_X1 _0903_ (.A(\mem[1][1] ),
    .B(_0338_),
    .S(_0372_),
    .Z(_0076_));
 MUX2_X1 _0904_ (.A(\mem[1][2] ),
    .B(_0340_),
    .S(_0372_),
    .Z(_0077_));
 MUX2_X1 _0905_ (.A(\mem[1][3] ),
    .B(_0342_),
    .S(_0372_),
    .Z(_0078_));
 MUX2_X1 _0906_ (.A(\mem[1][4] ),
    .B(_0344_),
    .S(_0372_),
    .Z(_0079_));
 MUX2_X1 _0907_ (.A(\mem[1][5] ),
    .B(_0346_),
    .S(_0372_),
    .Z(_0080_));
 MUX2_X1 _0908_ (.A(\mem[1][6] ),
    .B(_0348_),
    .S(_0372_),
    .Z(_0081_));
 MUX2_X1 _0909_ (.A(\mem[1][7] ),
    .B(_0350_),
    .S(_0372_),
    .Z(_0082_));
 AND4_X1 _0910_ (.A1(_0359_),
    .A2(_0182_),
    .A3(_0333_),
    .A4(_0353_),
    .ZN(_0373_));
 BUF_X8 _0911_ (.A(_0373_),
    .Z(_0374_));
 MUX2_X1 _0912_ (.A(\mem[2][0] ),
    .B(_0329_),
    .S(_0374_),
    .Z(_0083_));
 MUX2_X1 _0913_ (.A(\mem[2][1] ),
    .B(_0338_),
    .S(_0374_),
    .Z(_0084_));
 MUX2_X1 _0914_ (.A(\mem[2][2] ),
    .B(_0340_),
    .S(_0374_),
    .Z(_0085_));
 MUX2_X1 _0915_ (.A(\mem[2][3] ),
    .B(_0342_),
    .S(_0374_),
    .Z(_0086_));
 MUX2_X1 _0916_ (.A(\mem[2][4] ),
    .B(_0344_),
    .S(_0374_),
    .Z(_0087_));
 MUX2_X1 _0917_ (.A(\mem[2][5] ),
    .B(_0346_),
    .S(_0374_),
    .Z(_0088_));
 MUX2_X1 _0918_ (.A(\mem[2][6] ),
    .B(_0348_),
    .S(_0374_),
    .Z(_0089_));
 MUX2_X1 _0919_ (.A(\mem[2][7] ),
    .B(_0350_),
    .S(_0374_),
    .Z(_0090_));
 AND3_X1 _0920_ (.A1(_0177_),
    .A2(_0333_),
    .A3(_0356_),
    .ZN(_0375_));
 BUF_X4 _0921_ (.A(_0375_),
    .Z(_0376_));
 MUX2_X1 _0922_ (.A(\mem[3][0] ),
    .B(_0329_),
    .S(_0376_),
    .Z(_0091_));
 MUX2_X1 _0923_ (.A(\mem[3][1] ),
    .B(_0338_),
    .S(_0376_),
    .Z(_0092_));
 MUX2_X1 _0924_ (.A(\mem[3][2] ),
    .B(_0340_),
    .S(_0376_),
    .Z(_0093_));
 MUX2_X1 _0925_ (.A(\mem[3][3] ),
    .B(_0342_),
    .S(_0376_),
    .Z(_0094_));
 MUX2_X1 _0926_ (.A(\mem[3][4] ),
    .B(_0344_),
    .S(_0376_),
    .Z(_0095_));
 MUX2_X1 _0927_ (.A(\mem[3][5] ),
    .B(_0346_),
    .S(_0376_),
    .Z(_0096_));
 MUX2_X1 _0928_ (.A(\mem[3][6] ),
    .B(_0348_),
    .S(_0376_),
    .Z(_0097_));
 MUX2_X1 _0929_ (.A(\mem[3][7] ),
    .B(_0350_),
    .S(_0376_),
    .Z(_0098_));
 NOR2_X1 _0930_ (.A1(_0330_),
    .A2(_0332_),
    .ZN(_0377_));
 AND2_X1 _0931_ (.A1(_0331_),
    .A2(_0377_),
    .ZN(_0378_));
 AND4_X1 _0932_ (.A1(_0359_),
    .A2(_0182_),
    .A3(_0334_),
    .A4(_0378_),
    .ZN(_0379_));
 BUF_X8 _0933_ (.A(_0379_),
    .Z(_0380_));
 MUX2_X1 _0934_ (.A(\mem[4][0] ),
    .B(_0328_),
    .S(_0380_),
    .Z(_0099_));
 MUX2_X1 _0935_ (.A(\mem[4][1] ),
    .B(_0337_),
    .S(_0380_),
    .Z(_0100_));
 MUX2_X1 _0936_ (.A(\mem[4][2] ),
    .B(_0339_),
    .S(_0380_),
    .Z(_0101_));
 MUX2_X1 _0937_ (.A(\mem[4][3] ),
    .B(_0341_),
    .S(_0380_),
    .Z(_0102_));
 MUX2_X1 _0938_ (.A(\mem[4][4] ),
    .B(_0343_),
    .S(_0380_),
    .Z(_0103_));
 MUX2_X1 _0939_ (.A(\mem[4][5] ),
    .B(_0345_),
    .S(_0380_),
    .Z(_0104_));
 MUX2_X1 _0940_ (.A(\mem[4][6] ),
    .B(_0347_),
    .S(_0380_),
    .Z(_0105_));
 MUX2_X1 _0941_ (.A(\mem[4][7] ),
    .B(_0349_),
    .S(_0380_),
    .Z(_0106_));
 AND4_X1 _0942_ (.A1(_0359_),
    .A2(_0181_),
    .A3(_0364_),
    .A4(_0378_),
    .ZN(_0381_));
 BUF_X8 _0943_ (.A(_0381_),
    .Z(_0382_));
 MUX2_X1 _0944_ (.A(\mem[5][0] ),
    .B(_0328_),
    .S(_0382_),
    .Z(_0107_));
 MUX2_X1 _0945_ (.A(\mem[5][1] ),
    .B(_0337_),
    .S(_0382_),
    .Z(_0108_));
 MUX2_X1 _0946_ (.A(\mem[5][2] ),
    .B(_0339_),
    .S(_0382_),
    .Z(_0109_));
 MUX2_X1 _0947_ (.A(\mem[5][3] ),
    .B(_0341_),
    .S(_0382_),
    .Z(_0110_));
 MUX2_X1 _0948_ (.A(\mem[5][4] ),
    .B(_0343_),
    .S(_0382_),
    .Z(_0111_));
 MUX2_X1 _0949_ (.A(\mem[5][5] ),
    .B(_0345_),
    .S(_0382_),
    .Z(_0112_));
 MUX2_X1 _0950_ (.A(\mem[5][6] ),
    .B(_0347_),
    .S(_0382_),
    .Z(_0113_));
 MUX2_X1 _0951_ (.A(\mem[5][7] ),
    .B(_0349_),
    .S(_0382_),
    .Z(_0114_));
 AND4_X1 _0952_ (.A1(_0359_),
    .A2(_0181_),
    .A3(_0353_),
    .A4(_0378_),
    .ZN(_0383_));
 BUF_X8 _0953_ (.A(_0383_),
    .Z(_0384_));
 MUX2_X1 _0954_ (.A(\mem[6][0] ),
    .B(_0328_),
    .S(_0384_),
    .Z(_0115_));
 MUX2_X1 _0955_ (.A(\mem[6][1] ),
    .B(_0337_),
    .S(_0384_),
    .Z(_0116_));
 MUX2_X1 _0956_ (.A(\mem[6][2] ),
    .B(_0339_),
    .S(_0384_),
    .Z(_0117_));
 MUX2_X1 _0957_ (.A(\mem[6][3] ),
    .B(_0341_),
    .S(_0384_),
    .Z(_0118_));
 MUX2_X1 _0958_ (.A(\mem[6][4] ),
    .B(_0343_),
    .S(_0384_),
    .Z(_0119_));
 MUX2_X1 _0959_ (.A(\mem[6][5] ),
    .B(_0345_),
    .S(_0384_),
    .Z(_0120_));
 MUX2_X1 _0960_ (.A(\mem[6][6] ),
    .B(_0347_),
    .S(_0384_),
    .Z(_0121_));
 MUX2_X1 _0961_ (.A(\mem[6][7] ),
    .B(_0349_),
    .S(_0384_),
    .Z(_0122_));
 AND3_X1 _0962_ (.A1(_0177_),
    .A2(_0356_),
    .A3(_0378_),
    .ZN(_0385_));
 BUF_X4 _0963_ (.A(_0385_),
    .Z(_0386_));
 MUX2_X1 _0964_ (.A(\mem[7][0] ),
    .B(_0328_),
    .S(_0386_),
    .Z(_0123_));
 MUX2_X1 _0965_ (.A(\mem[7][1] ),
    .B(_0337_),
    .S(_0386_),
    .Z(_0124_));
 MUX2_X1 _0966_ (.A(\mem[7][2] ),
    .B(_0339_),
    .S(_0386_),
    .Z(_0125_));
 MUX2_X1 _0967_ (.A(\mem[7][3] ),
    .B(_0341_),
    .S(_0386_),
    .Z(_0126_));
 MUX2_X1 _0968_ (.A(\mem[7][4] ),
    .B(_0343_),
    .S(_0386_),
    .Z(_0127_));
 MUX2_X1 _0969_ (.A(\mem[7][5] ),
    .B(_0345_),
    .S(_0386_),
    .Z(_0128_));
 MUX2_X1 _0970_ (.A(\mem[7][6] ),
    .B(_0347_),
    .S(_0386_),
    .Z(_0129_));
 MUX2_X1 _0971_ (.A(\mem[7][7] ),
    .B(_0349_),
    .S(_0386_),
    .Z(_0130_));
 AND4_X1 _0972_ (.A1(_0359_),
    .A2(_0181_),
    .A3(_0334_),
    .A4(_0352_),
    .ZN(_0387_));
 BUF_X8 _0973_ (.A(_0387_),
    .Z(_0388_));
 MUX2_X1 _0974_ (.A(\mem[8][0] ),
    .B(_0328_),
    .S(_0388_),
    .Z(_0131_));
 MUX2_X1 _0975_ (.A(\mem[8][1] ),
    .B(_0337_),
    .S(_0388_),
    .Z(_0132_));
 MUX2_X1 _0976_ (.A(\mem[8][2] ),
    .B(_0339_),
    .S(_0388_),
    .Z(_0133_));
 MUX2_X1 _0977_ (.A(\mem[8][3] ),
    .B(_0341_),
    .S(_0388_),
    .Z(_0134_));
 MUX2_X1 _0978_ (.A(\mem[8][4] ),
    .B(_0343_),
    .S(_0388_),
    .Z(_0135_));
 MUX2_X1 _0979_ (.A(\mem[8][5] ),
    .B(_0345_),
    .S(_0388_),
    .Z(_0136_));
 MUX2_X1 _0980_ (.A(\mem[8][6] ),
    .B(_0347_),
    .S(_0388_),
    .Z(_0137_));
 MUX2_X1 _0981_ (.A(\mem[8][7] ),
    .B(_0349_),
    .S(_0388_),
    .Z(_0138_));
 AND4_X1 _0982_ (.A1(_0359_),
    .A2(_0181_),
    .A3(_0352_),
    .A4(_0364_),
    .ZN(_0389_));
 BUF_X8 _0983_ (.A(_0389_),
    .Z(_0390_));
 MUX2_X1 _0984_ (.A(\mem[9][0] ),
    .B(_0328_),
    .S(_0390_),
    .Z(_0139_));
 MUX2_X1 _0985_ (.A(\mem[9][1] ),
    .B(_0337_),
    .S(_0390_),
    .Z(_0140_));
 MUX2_X1 _0986_ (.A(\mem[9][2] ),
    .B(_0339_),
    .S(_0390_),
    .Z(_0141_));
 MUX2_X1 _0987_ (.A(\mem[9][3] ),
    .B(_0341_),
    .S(_0390_),
    .Z(_0142_));
 MUX2_X1 _0988_ (.A(\mem[9][4] ),
    .B(_0343_),
    .S(_0390_),
    .Z(_0143_));
 MUX2_X1 _0989_ (.A(\mem[9][5] ),
    .B(_0345_),
    .S(_0390_),
    .Z(_0144_));
 MUX2_X1 _0990_ (.A(\mem[9][6] ),
    .B(_0347_),
    .S(_0390_),
    .Z(_0145_));
 MUX2_X1 _0991_ (.A(\mem[9][7] ),
    .B(_0349_),
    .S(_0390_),
    .Z(_0146_));
 BUF_X2 _0992_ (.A(_0186_),
    .Z(_0391_));
 AND2_X1 _0993_ (.A1(_0178_),
    .A2(_0584_),
    .ZN(_0392_));
 INV_X1 _0994_ (.A(_0599_),
    .ZN(_0393_));
 AOI21_X1 _0995_ (.A(_0393_),
    .B1(_0180_),
    .B2(net4),
    .ZN(_0394_));
 AOI221_X2 _0996_ (.A(_0597_),
    .B1(_0180_),
    .B2(_0392_),
    .C1(_0394_),
    .C2(net8),
    .ZN(_0395_));
 MUX2_X1 _0997_ (.A(net4),
    .B(_0000_),
    .S(_0395_),
    .Z(_0396_));
 AND2_X1 _0998_ (.A1(_0391_),
    .A2(_0396_),
    .ZN(_0006_));
 MUX2_X1 _0999_ (.A(net5),
    .B(_0005_),
    .S(_0395_),
    .Z(_0397_));
 AND2_X1 _1000_ (.A1(_0391_),
    .A2(_0397_),
    .ZN(_0007_));
 XOR2_X1 _1001_ (.A(_0585_),
    .B(_0612_),
    .Z(_0398_));
 MUX2_X1 _1002_ (.A(net6),
    .B(_0398_),
    .S(_0395_),
    .Z(_0399_));
 AND2_X1 _1003_ (.A1(_0391_),
    .A2(_0399_),
    .ZN(_0008_));
 AOI21_X1 _1004_ (.A(_0609_),
    .B1(_0610_),
    .B2(net4),
    .ZN(_0400_));
 INV_X1 _1005_ (.A(_0400_),
    .ZN(_0401_));
 AOI21_X1 _1006_ (.A(_0611_),
    .B1(_0401_),
    .B2(_0612_),
    .ZN(_0402_));
 XNOR2_X1 _1007_ (.A(_0614_),
    .B(_0402_),
    .ZN(_0403_));
 MUX2_X1 _1008_ (.A(net7),
    .B(_0403_),
    .S(_0395_),
    .Z(_0404_));
 AND2_X1 _1009_ (.A1(_0391_),
    .A2(_0404_),
    .ZN(_0009_));
 AOI21_X1 _1010_ (.A(_0611_),
    .B1(_0612_),
    .B2(_0585_),
    .ZN(_0405_));
 INV_X1 _1011_ (.A(_0405_),
    .ZN(_0406_));
 AOI21_X1 _1012_ (.A(_0613_),
    .B1(_0406_),
    .B2(_0614_),
    .ZN(_0407_));
 XNOR2_X1 _1013_ (.A(_0584_),
    .B(_0407_),
    .ZN(_0408_));
 AOI21_X1 _1014_ (.A(net8),
    .B1(_0395_),
    .B2(_0408_),
    .ZN(_0409_));
 AND3_X1 _1015_ (.A1(net8),
    .A2(_0395_),
    .A3(_0408_),
    .ZN(_0410_));
 OAI21_X1 _1016_ (.A(_0391_),
    .B1(_0409_),
    .B2(_0410_),
    .ZN(_0010_));
 MUX2_X1 _1017_ (.A(_0196_),
    .B(_0003_),
    .S(_0188_),
    .Z(_0411_));
 AND2_X1 _1018_ (.A1(_0391_),
    .A2(_0411_),
    .ZN(_0147_));
 MUX2_X1 _1019_ (.A(_0192_),
    .B(_0004_),
    .S(_0188_),
    .Z(_0412_));
 AND2_X1 _1020_ (.A1(_0391_),
    .A2(_0412_),
    .ZN(_0148_));
 NAND2_X1 _1021_ (.A1(_0601_),
    .A2(_0188_),
    .ZN(_0413_));
 XNOR2_X1 _1022_ (.A(_0206_),
    .B(_0413_),
    .ZN(_0414_));
 NOR2_X1 _1023_ (.A1(_0330_),
    .A2(_0414_),
    .ZN(_0149_));
 NAND4_X1 _1024_ (.A1(_0196_),
    .A2(_0192_),
    .A3(_0204_),
    .A4(_0188_),
    .ZN(_0415_));
 XOR2_X1 _1025_ (.A(_0202_),
    .B(_0415_),
    .Z(_0416_));
 NOR2_X1 _1026_ (.A1(_0330_),
    .A2(_0416_),
    .ZN(_0150_));
 NAND4_X1 _1027_ (.A1(_0204_),
    .A2(_0202_),
    .A3(_0601_),
    .A4(_0188_),
    .ZN(_0417_));
 XOR2_X1 _1028_ (.A(\read_ptr[4] ),
    .B(_0417_),
    .Z(_0418_));
 NOR2_X1 _1029_ (.A1(_0330_),
    .A2(_0418_),
    .ZN(_0151_));
 NAND2_X1 _1030_ (.A1(net25),
    .A2(_0187_),
    .ZN(_0419_));
 AOI21_X1 _1031_ (.A(_0330_),
    .B1(net17),
    .B2(_0419_),
    .ZN(_0152_));
 AND2_X1 _1032_ (.A1(_0186_),
    .A2(\write_ptr[0] ),
    .ZN(_0420_));
 AND2_X1 _1033_ (.A1(_0391_),
    .A2(_0001_),
    .ZN(_0421_));
 MUX2_X1 _1034_ (.A(_0420_),
    .B(_0421_),
    .S(_0595_),
    .Z(_0153_));
 AND2_X1 _1035_ (.A1(_0186_),
    .A2(\write_ptr[1] ),
    .ZN(_0422_));
 AND2_X1 _1036_ (.A1(_0391_),
    .A2(_0002_),
    .ZN(_0423_));
 MUX2_X1 _1037_ (.A(_0422_),
    .B(_0423_),
    .S(_0595_),
    .Z(_0154_));
 NAND2_X1 _1038_ (.A1(_0177_),
    .A2(_0356_),
    .ZN(_0424_));
 MUX2_X1 _1039_ (.A(_0351_),
    .B(_0360_),
    .S(_0424_),
    .Z(_0155_));
 AND2_X1 _1040_ (.A1(_0391_),
    .A2(_0332_),
    .ZN(_0425_));
 NAND3_X1 _1041_ (.A1(_0331_),
    .A2(\write_ptr[1] ),
    .A3(\write_ptr[0] ),
    .ZN(_0426_));
 NOR3_X1 _1042_ (.A1(net23),
    .A2(_0183_),
    .A3(_0426_),
    .ZN(_0427_));
 MUX2_X1 _1043_ (.A(_0425_),
    .B(_0377_),
    .S(_0427_),
    .Z(_0156_));
 AND2_X1 _1044_ (.A1(_0168_),
    .A2(_0186_),
    .ZN(_0428_));
 NOR2_X1 _1045_ (.A1(_0168_),
    .A2(_0330_),
    .ZN(_0429_));
 AND4_X1 _1046_ (.A1(_0331_),
    .A2(_0332_),
    .A3(_0177_),
    .A4(_0356_),
    .ZN(_0430_));
 MUX2_X1 _1047_ (.A(_0428_),
    .B(_0429_),
    .S(_0430_),
    .Z(_0157_));
 XNOR2_X1 _1048_ (.A(_0158_),
    .B(_0167_),
    .ZN(net21));
 NOR3_X1 _1049_ (.A1(_0169_),
    .A2(_0172_),
    .A3(_0173_),
    .ZN(_0431_));
 INV_X1 _1050_ (.A(_0590_),
    .ZN(_0432_));
 INV_X1 _1051_ (.A(_0160_),
    .ZN(_0433_));
 OAI21_X1 _1052_ (.A(_0432_),
    .B1(_0433_),
    .B2(_0583_),
    .ZN(_0434_));
 AOI211_X2 _1053_ (.A(_0587_),
    .B(_0184_),
    .C1(_0434_),
    .C2(_0158_),
    .ZN(_0435_));
 NOR2_X1 _1054_ (.A1(_0431_),
    .A2(_0435_),
    .ZN(net22));
 AND2_X1 _1055_ (.A1(_0177_),
    .A2(_0182_),
    .ZN(net24));
 FA_X1 _1056_ (.A(\read_ptr[1] ),
    .B(_0581_),
    .CI(_0582_),
    .CO(_0583_),
    .S(net19));
 FA_X1 _1057_ (.A(net4),
    .B(net5),
    .CI(_0584_),
    .CO(_0585_),
    .S(_0005_));
 HA_X1 _1058_ (.A(_0586_),
    .B(\write_ptr[3] ),
    .CO(_0587_),
    .S(_0588_));
 HA_X1 _1059_ (.A(_0589_),
    .B(\write_ptr[2] ),
    .CO(_0590_),
    .S(_0591_));
 HA_X1 _1060_ (.A(_0593_),
    .B(\write_ptr[1] ),
    .CO(_0594_),
    .S(_0592_));
 HA_X1 _1061_ (.A(_0595_),
    .B(_0596_),
    .CO(_0584_),
    .S(_0597_));
 HA_X1 _1062_ (.A(_0598_),
    .B(net1),
    .CO(_0599_),
    .S(_0600_));
 HA_X1 _1063_ (.A(\read_ptr[0] ),
    .B(\read_ptr[1] ),
    .CO(_0601_),
    .S(_0004_));
 HA_X1 _1064_ (.A(_0001_),
    .B(_0581_),
    .CO(_0602_),
    .S(_0002_));
 HA_X1 _1065_ (.A(_0001_),
    .B(\write_ptr[1] ),
    .CO(_0603_),
    .S(_0604_));
 HA_X1 _1066_ (.A(\write_ptr[0] ),
    .B(_0581_),
    .CO(_0605_),
    .S(_0606_));
 HA_X1 _1067_ (.A(\write_ptr[0] ),
    .B(\write_ptr[1] ),
    .CO(_0607_),
    .S(_0608_));
 HA_X1 _1068_ (.A(net5),
    .B(_0584_),
    .CO(_0609_),
    .S(_0610_));
 HA_X1 _1069_ (.A(net6),
    .B(_0584_),
    .CO(_0611_),
    .S(_0612_));
 HA_X1 _1070_ (.A(net7),
    .B(_0584_),
    .CO(_0613_),
    .S(_0614_));
 HA_X1 _1071_ (.A(\read_ptr[0] ),
    .B(_0001_),
    .CO(_0582_),
    .S(_0615_));
 DFF_X2 \credit_count[0]$_SDFFE_PN0P_  (.D(_0006_),
    .CK(clknet_4_5_0_clk),
    .Q(net4),
    .QN(_0000_));
 DFF_X2 \credit_count[1]$_SDFFE_PN0P_  (.D(_0007_),
    .CK(clknet_4_5_0_clk),
    .Q(net5),
    .QN(_0580_));
 DFF_X2 \credit_count[2]$_SDFFE_PN0P_  (.D(_0008_),
    .CK(clknet_4_5_0_clk),
    .Q(net6),
    .QN(_0579_));
 DFF_X2 \credit_count[3]$_SDFFE_PN0P_  (.D(_0009_),
    .CK(clknet_4_5_0_clk),
    .Q(net7),
    .QN(_0578_));
 DFF_X2 \credit_count[4]$_SDFFE_PN1P_  (.D(_0010_),
    .CK(clknet_4_5_0_clk),
    .Q(net8),
    .QN(_0577_));
 DFF_X1 \data_out[0]$_DFFE_PP_  (.D(_0011_),
    .CK(clknet_4_13_0_clk),
    .Q(net9),
    .QN(_0576_));
 DFF_X1 \data_out[1]$_DFFE_PP_  (.D(_0012_),
    .CK(clknet_4_8_0_clk),
    .Q(net10),
    .QN(_0575_));
 DFF_X1 \data_out[2]$_DFFE_PP_  (.D(_0013_),
    .CK(clknet_4_10_0_clk),
    .Q(net11),
    .QN(_0574_));
 DFF_X1 \data_out[3]$_DFFE_PP_  (.D(_0014_),
    .CK(clknet_4_15_0_clk),
    .Q(net12),
    .QN(_0573_));
 DFF_X1 \data_out[4]$_DFFE_PP_  (.D(_0015_),
    .CK(clknet_4_11_0_clk),
    .Q(net13),
    .QN(_0572_));
 DFF_X1 \data_out[5]$_DFFE_PP_  (.D(_0016_),
    .CK(clknet_4_10_0_clk),
    .Q(net14),
    .QN(_0571_));
 DFF_X1 \data_out[6]$_DFFE_PP_  (.D(_0017_),
    .CK(clknet_4_14_0_clk),
    .Q(net15),
    .QN(_0570_));
 DFF_X1 \data_out[7]$_DFFE_PP_  (.D(_0018_),
    .CK(clknet_4_9_0_clk),
    .Q(net16),
    .QN(_0569_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0019_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[0][0] ),
    .QN(_0568_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0020_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[0][1] ),
    .QN(_0567_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0021_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[0][2] ),
    .QN(_0566_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0022_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[0][3] ),
    .QN(_0565_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0023_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[0][4] ),
    .QN(_0564_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0024_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[0][5] ),
    .QN(_0563_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0025_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[0][6] ),
    .QN(_0562_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0026_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[0][7] ),
    .QN(_0561_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0027_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[10][0] ),
    .QN(_0560_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0028_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][1] ),
    .QN(_0559_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0029_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][2] ),
    .QN(_0558_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0030_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[10][3] ),
    .QN(_0557_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0031_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[10][4] ),
    .QN(_0556_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0032_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[10][5] ),
    .QN(_0555_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0033_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[10][6] ),
    .QN(_0554_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0034_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[10][7] ),
    .QN(_0553_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0035_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[11][0] ),
    .QN(_0552_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0036_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][1] ),
    .QN(_0551_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0037_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][2] ),
    .QN(_0550_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0038_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[11][3] ),
    .QN(_0549_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0039_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[11][4] ),
    .QN(_0548_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0040_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[11][5] ),
    .QN(_0547_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0041_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[11][6] ),
    .QN(_0546_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0042_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[11][7] ),
    .QN(_0545_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0043_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[12][0] ),
    .QN(_0544_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0044_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[12][1] ),
    .QN(_0543_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0045_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[12][2] ),
    .QN(_0542_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[12][3] ),
    .QN(_0541_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[12][4] ),
    .QN(_0540_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[12][5] ),
    .QN(_0539_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[12][6] ),
    .QN(_0538_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[12][7] ),
    .QN(_0537_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[13][0] ),
    .QN(_0536_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[13][1] ),
    .QN(_0535_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[13][2] ),
    .QN(_0534_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[13][3] ),
    .QN(_0533_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[13][4] ),
    .QN(_0532_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[13][5] ),
    .QN(_0531_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[13][6] ),
    .QN(_0530_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[13][7] ),
    .QN(_0529_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_4_13_0_clk),
    .Q(\mem[14][0] ),
    .QN(_0528_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0060_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[14][1] ),
    .QN(_0527_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0061_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[14][2] ),
    .QN(_0526_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0062_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[14][3] ),
    .QN(_0525_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0063_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[14][4] ),
    .QN(_0524_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[14][5] ),
    .QN(_0523_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[14][6] ),
    .QN(_0522_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[14][7] ),
    .QN(_0521_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[15][0] ),
    .QN(_0520_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[15][1] ),
    .QN(_0519_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[15][2] ),
    .QN(_0518_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[15][3] ),
    .QN(_0517_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[15][4] ),
    .QN(_0516_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_4_11_0_clk),
    .Q(\mem[15][5] ),
    .QN(_0515_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[15][6] ),
    .QN(_0514_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_4_9_0_clk),
    .Q(\mem[15][7] ),
    .QN(_0513_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[1][0] ),
    .QN(_0512_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[1][1] ),
    .QN(_0511_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[1][2] ),
    .QN(_0510_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[1][3] ),
    .QN(_0509_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[1][4] ),
    .QN(_0508_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[1][5] ),
    .QN(_0507_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[1][6] ),
    .QN(_0506_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[1][7] ),
    .QN(_0505_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[2][0] ),
    .QN(_0504_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[2][1] ),
    .QN(_0503_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[2][2] ),
    .QN(_0502_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[2][3] ),
    .QN(_0501_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[2][4] ),
    .QN(_0500_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[2][5] ),
    .QN(_0499_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[2][6] ),
    .QN(_0498_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[2][7] ),
    .QN(_0497_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_4_15_0_clk),
    .Q(\mem[3][0] ),
    .QN(_0496_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[3][1] ),
    .QN(_0495_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_4_8_0_clk),
    .Q(\mem[3][2] ),
    .QN(_0494_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[3][3] ),
    .QN(_0493_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[3][4] ),
    .QN(_0492_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_4_10_0_clk),
    .Q(\mem[3][5] ),
    .QN(_0491_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_4_14_0_clk),
    .Q(\mem[3][6] ),
    .QN(_0490_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_4_12_0_clk),
    .Q(\mem[3][7] ),
    .QN(_0489_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[4][0] ),
    .QN(_0488_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[4][1] ),
    .QN(_0487_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[4][2] ),
    .QN(_0486_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[4][3] ),
    .QN(_0485_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[4][4] ),
    .QN(_0484_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[4][5] ),
    .QN(_0483_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[4][6] ),
    .QN(_0482_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[4][7] ),
    .QN(_0481_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[5][0] ),
    .QN(_0480_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[5][1] ),
    .QN(_0479_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[5][2] ),
    .QN(_0478_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[5][3] ),
    .QN(_0477_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[5][4] ),
    .QN(_0476_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[5][5] ),
    .QN(_0475_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[5][6] ),
    .QN(_0474_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[5][7] ),
    .QN(_0473_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[6][0] ),
    .QN(_0472_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[6][1] ),
    .QN(_0471_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[6][2] ),
    .QN(_0470_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[6][3] ),
    .QN(_0469_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[6][4] ),
    .QN(_0468_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[6][5] ),
    .QN(_0467_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[6][6] ),
    .QN(_0466_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[6][7] ),
    .QN(_0465_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_4_5_0_clk),
    .Q(\mem[7][0] ),
    .QN(_0464_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_4_0_0_clk),
    .Q(\mem[7][1] ),
    .QN(_0463_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[7][2] ),
    .QN(_0462_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[7][3] ),
    .QN(_0461_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[7][4] ),
    .QN(_0460_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[7][5] ),
    .QN(_0459_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[7][6] ),
    .QN(_0458_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_4_1_0_clk),
    .Q(\mem[7][7] ),
    .QN(_0457_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[8][0] ),
    .QN(_0456_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[8][1] ),
    .QN(_0455_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[8][2] ),
    .QN(_0454_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[8][3] ),
    .QN(_0453_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[8][4] ),
    .QN(_0452_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[8][5] ),
    .QN(_0451_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_4_4_0_clk),
    .Q(\mem[8][6] ),
    .QN(_0450_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[8][7] ),
    .QN(_0449_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[9][0] ),
    .QN(_0448_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[9][1] ),
    .QN(_0447_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[9][2] ),
    .QN(_0446_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_4_7_0_clk),
    .Q(\mem[9][3] ),
    .QN(_0445_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[9][4] ),
    .QN(_0444_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_4_2_0_clk),
    .Q(\mem[9][5] ),
    .QN(_0443_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_4_6_0_clk),
    .Q(\mem[9][6] ),
    .QN(_0442_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_4_3_0_clk),
    .Q(\mem[9][7] ),
    .QN(_0441_));
 DFF_X2 \read_ptr[0]$_SDFFE_PN0P_  (.D(_0147_),
    .CK(clknet_4_13_0_clk),
    .Q(\read_ptr[0] ),
    .QN(_0003_));
 DFF_X2 \read_ptr[1]$_SDFFE_PN0P_  (.D(_0148_),
    .CK(clknet_4_13_0_clk),
    .Q(\read_ptr[1] ),
    .QN(_0593_));
 DFF_X1 \read_ptr[2]$_SDFFE_PN0P_  (.D(_0149_),
    .CK(clknet_4_13_0_clk),
    .Q(\read_ptr[2] ),
    .QN(_0589_));
 DFF_X1 \read_ptr[3]$_SDFFE_PN0P_  (.D(_0150_),
    .CK(clknet_4_13_0_clk),
    .Q(\read_ptr[3] ),
    .QN(_0586_));
 DFF_X2 \read_ptr[4]$_SDFFE_PN0P_  (.D(_0151_),
    .CK(clknet_4_15_0_clk),
    .Q(\read_ptr[4] ),
    .QN(_0440_));
 DFF_X2 \valid_out$_SDFFE_PN0P_  (.D(_0152_),
    .CK(clknet_4_15_0_clk),
    .Q(net25),
    .QN(_0439_));
 DFF_X2 \write_ptr[0]$_SDFFE_PN0N_  (.D(_0153_),
    .CK(clknet_4_5_0_clk),
    .Q(\write_ptr[0] ),
    .QN(_0001_));
 DFF_X2 \write_ptr[1]$_SDFFE_PN0N_  (.D(_0154_),
    .CK(clknet_4_7_0_clk),
    .Q(\write_ptr[1] ),
    .QN(_0581_));
 DFF_X1 \write_ptr[2]$_SDFFE_PN0N_  (.D(_0155_),
    .CK(clknet_4_7_0_clk),
    .Q(\write_ptr[2] ),
    .QN(_0438_));
 DFF_X1 \write_ptr[3]$_SDFFE_PN0N_  (.D(_0156_),
    .CK(clknet_4_7_0_clk),
    .Q(\write_ptr[3] ),
    .QN(_0437_));
 DFF_X1 \write_ptr[4]$_SDFFE_PN0N_  (.D(_0157_),
    .CK(clknet_4_15_0_clk),
    .Q(\write_ptr[4] ),
    .QN(_0436_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_75 ();
 BUF_X1 input1 (.A(credit_return),
    .Z(net1));
 BUF_X1 input2 (.A(ready_in),
    .Z(net2));
 BUF_X1 input3 (.A(valid_in),
    .Z(net3));
 BUF_X1 output4 (.A(net4),
    .Z(credits_available[0]));
 BUF_X1 output5 (.A(net5),
    .Z(credits_available[1]));
 BUF_X1 output6 (.A(net6),
    .Z(credits_available[2]));
 BUF_X1 output7 (.A(net7),
    .Z(credits_available[3]));
 BUF_X1 output8 (.A(net8),
    .Z(credits_available[4]));
 BUF_X1 output9 (.A(net9),
    .Z(data_out[0]));
 BUF_X1 output10 (.A(net10),
    .Z(data_out[1]));
 BUF_X1 output11 (.A(net11),
    .Z(data_out[2]));
 BUF_X1 output12 (.A(net12),
    .Z(data_out[3]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[4]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[5]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[6]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[7]));
 BUF_X1 output17 (.A(net17),
    .Z(empty));
 BUF_X1 output18 (.A(net18),
    .Z(fifo_level[0]));
 BUF_X1 output19 (.A(net19),
    .Z(fifo_level[1]));
 BUF_X1 output20 (.A(net20),
    .Z(fifo_level[2]));
 BUF_X1 output21 (.A(net21),
    .Z(fifo_level[3]));
 BUF_X1 output22 (.A(net22),
    .Z(fifo_level[4]));
 BUF_X1 output23 (.A(net23),
    .Z(full));
 BUF_X1 output24 (.A(net24),
    .Z(ready_out));
 BUF_X1 output25 (.A(net25),
    .Z(valid_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X2 clkload0 (.A(clknet_4_0_0_clk));
 INV_X2 clkload1 (.A(clknet_4_1_0_clk));
 INV_X1 clkload2 (.A(clknet_4_3_0_clk));
 INV_X2 clkload3 (.A(clknet_4_4_0_clk));
 CLKBUF_X1 clkload4 (.A(clknet_4_5_0_clk));
 INV_X2 clkload5 (.A(clknet_4_6_0_clk));
 INV_X4 clkload6 (.A(clknet_4_7_0_clk));
 INV_X2 clkload7 (.A(clknet_4_8_0_clk));
 INV_X2 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_10_0_clk));
 INV_X2 clkload10 (.A(clknet_4_11_0_clk));
 INV_X4 clkload11 (.A(clknet_4_12_0_clk));
 INV_X2 clkload12 (.A(clknet_4_13_0_clk));
 INV_X2 clkload13 (.A(clknet_4_14_0_clk));
 CLKBUF_X1 clkload14 (.A(clknet_4_15_0_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_73 ();
 FILLCELL_X1 FILLER_0_77 ();
 FILLCELL_X32 FILLER_0_89 ();
 FILLCELL_X32 FILLER_0_121 ();
 FILLCELL_X16 FILLER_0_153 ();
 FILLCELL_X8 FILLER_0_169 ();
 FILLCELL_X4 FILLER_0_180 ();
 FILLCELL_X8 FILLER_0_187 ();
 FILLCELL_X1 FILLER_0_195 ();
 FILLCELL_X32 FILLER_0_216 ();
 FILLCELL_X32 FILLER_0_248 ();
 FILLCELL_X2 FILLER_0_280 ();
 FILLCELL_X1 FILLER_0_282 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X8 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_73 ();
 FILLCELL_X1 FILLER_1_77 ();
 FILLCELL_X2 FILLER_1_85 ();
 FILLCELL_X1 FILLER_1_87 ();
 FILLCELL_X1 FILLER_1_105 ();
 FILLCELL_X2 FILLER_1_113 ();
 FILLCELL_X1 FILLER_1_132 ();
 FILLCELL_X2 FILLER_1_140 ();
 FILLCELL_X1 FILLER_1_142 ();
 FILLCELL_X2 FILLER_1_167 ();
 FILLCELL_X1 FILLER_1_176 ();
 FILLCELL_X1 FILLER_1_194 ();
 FILLCELL_X32 FILLER_1_215 ();
 FILLCELL_X32 FILLER_1_247 ();
 FILLCELL_X4 FILLER_1_279 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_65 ();
 FILLCELL_X1 FILLER_2_73 ();
 FILLCELL_X2 FILLER_2_91 ();
 FILLCELL_X2 FILLER_2_100 ();
 FILLCELL_X1 FILLER_2_102 ();
 FILLCELL_X1 FILLER_2_120 ();
 FILLCELL_X4 FILLER_2_138 ();
 FILLCELL_X1 FILLER_2_142 ();
 FILLCELL_X1 FILLER_2_177 ();
 FILLCELL_X16 FILLER_2_195 ();
 FILLCELL_X8 FILLER_2_211 ();
 FILLCELL_X4 FILLER_2_219 ();
 FILLCELL_X2 FILLER_2_223 ();
 FILLCELL_X32 FILLER_2_242 ();
 FILLCELL_X8 FILLER_2_274 ();
 FILLCELL_X1 FILLER_2_282 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_73 ();
 FILLCELL_X2 FILLER_3_77 ();
 FILLCELL_X1 FILLER_3_79 ();
 FILLCELL_X4 FILLER_3_104 ();
 FILLCELL_X2 FILLER_3_115 ();
 FILLCELL_X1 FILLER_3_124 ();
 FILLCELL_X8 FILLER_3_136 ();
 FILLCELL_X4 FILLER_3_144 ();
 FILLCELL_X1 FILLER_3_148 ();
 FILLCELL_X2 FILLER_3_170 ();
 FILLCELL_X2 FILLER_3_179 ();
 FILLCELL_X4 FILLER_3_202 ();
 FILLCELL_X2 FILLER_3_208 ();
 FILLCELL_X1 FILLER_3_210 ();
 FILLCELL_X32 FILLER_3_242 ();
 FILLCELL_X8 FILLER_3_274 ();
 FILLCELL_X1 FILLER_3_282 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_25 ();
 FILLCELL_X2 FILLER_4_29 ();
 FILLCELL_X32 FILLER_4_48 ();
 FILLCELL_X8 FILLER_4_80 ();
 FILLCELL_X8 FILLER_4_95 ();
 FILLCELL_X4 FILLER_4_103 ();
 FILLCELL_X1 FILLER_4_107 ();
 FILLCELL_X32 FILLER_4_112 ();
 FILLCELL_X16 FILLER_4_144 ();
 FILLCELL_X8 FILLER_4_160 ();
 FILLCELL_X4 FILLER_4_168 ();
 FILLCELL_X16 FILLER_4_186 ();
 FILLCELL_X8 FILLER_4_202 ();
 FILLCELL_X4 FILLER_4_210 ();
 FILLCELL_X2 FILLER_4_214 ();
 FILLCELL_X8 FILLER_4_223 ();
 FILLCELL_X16 FILLER_4_255 ();
 FILLCELL_X8 FILLER_4_271 ();
 FILLCELL_X4 FILLER_4_279 ();
 FILLCELL_X2 FILLER_5_1 ();
 FILLCELL_X1 FILLER_5_3 ();
 FILLCELL_X1 FILLER_5_38 ();
 FILLCELL_X1 FILLER_5_46 ();
 FILLCELL_X4 FILLER_5_64 ();
 FILLCELL_X2 FILLER_5_68 ();
 FILLCELL_X1 FILLER_5_70 ();
 FILLCELL_X2 FILLER_5_88 ();
 FILLCELL_X1 FILLER_5_90 ();
 FILLCELL_X8 FILLER_5_95 ();
 FILLCELL_X4 FILLER_5_103 ();
 FILLCELL_X2 FILLER_5_107 ();
 FILLCELL_X1 FILLER_5_109 ();
 FILLCELL_X8 FILLER_5_134 ();
 FILLCELL_X2 FILLER_5_142 ();
 FILLCELL_X1 FILLER_5_144 ();
 FILLCELL_X2 FILLER_5_169 ();
 FILLCELL_X8 FILLER_5_195 ();
 FILLCELL_X4 FILLER_5_203 ();
 FILLCELL_X32 FILLER_5_238 ();
 FILLCELL_X8 FILLER_5_270 ();
 FILLCELL_X4 FILLER_5_278 ();
 FILLCELL_X1 FILLER_5_282 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_47 ();
 FILLCELL_X1 FILLER_6_55 ();
 FILLCELL_X8 FILLER_6_77 ();
 FILLCELL_X4 FILLER_6_85 ();
 FILLCELL_X1 FILLER_6_89 ();
 FILLCELL_X4 FILLER_6_104 ();
 FILLCELL_X1 FILLER_6_108 ();
 FILLCELL_X1 FILLER_6_133 ();
 FILLCELL_X4 FILLER_6_141 ();
 FILLCELL_X1 FILLER_6_145 ();
 FILLCELL_X4 FILLER_6_153 ();
 FILLCELL_X1 FILLER_6_157 ();
 FILLCELL_X1 FILLER_6_165 ();
 FILLCELL_X1 FILLER_6_173 ();
 FILLCELL_X1 FILLER_6_188 ();
 FILLCELL_X1 FILLER_6_203 ();
 FILLCELL_X2 FILLER_6_211 ();
 FILLCELL_X1 FILLER_6_213 ();
 FILLCELL_X4 FILLER_6_221 ();
 FILLCELL_X2 FILLER_6_225 ();
 FILLCELL_X8 FILLER_6_232 ();
 FILLCELL_X2 FILLER_6_240 ();
 FILLCELL_X16 FILLER_6_259 ();
 FILLCELL_X8 FILLER_6_275 ();
 FILLCELL_X8 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_9 ();
 FILLCELL_X2 FILLER_7_13 ();
 FILLCELL_X8 FILLER_7_29 ();
 FILLCELL_X4 FILLER_7_37 ();
 FILLCELL_X2 FILLER_7_41 ();
 FILLCELL_X1 FILLER_7_43 ();
 FILLCELL_X16 FILLER_7_51 ();
 FILLCELL_X2 FILLER_7_67 ();
 FILLCELL_X2 FILLER_7_100 ();
 FILLCELL_X1 FILLER_7_102 ();
 FILLCELL_X8 FILLER_7_117 ();
 FILLCELL_X2 FILLER_7_125 ();
 FILLCELL_X1 FILLER_7_127 ();
 FILLCELL_X2 FILLER_7_135 ();
 FILLCELL_X1 FILLER_7_137 ();
 FILLCELL_X16 FILLER_7_162 ();
 FILLCELL_X8 FILLER_7_192 ();
 FILLCELL_X2 FILLER_7_200 ();
 FILLCELL_X4 FILLER_7_216 ();
 FILLCELL_X4 FILLER_7_227 ();
 FILLCELL_X16 FILLER_7_255 ();
 FILLCELL_X8 FILLER_7_271 ();
 FILLCELL_X4 FILLER_7_279 ();
 FILLCELL_X2 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_3 ();
 FILLCELL_X8 FILLER_8_21 ();
 FILLCELL_X4 FILLER_8_29 ();
 FILLCELL_X1 FILLER_8_54 ();
 FILLCELL_X8 FILLER_8_72 ();
 FILLCELL_X1 FILLER_8_80 ();
 FILLCELL_X2 FILLER_8_88 ();
 FILLCELL_X16 FILLER_8_138 ();
 FILLCELL_X8 FILLER_8_154 ();
 FILLCELL_X2 FILLER_8_162 ();
 FILLCELL_X8 FILLER_8_171 ();
 FILLCELL_X4 FILLER_8_179 ();
 FILLCELL_X2 FILLER_8_183 ();
 FILLCELL_X1 FILLER_8_185 ();
 FILLCELL_X8 FILLER_8_193 ();
 FILLCELL_X2 FILLER_8_201 ();
 FILLCELL_X2 FILLER_8_210 ();
 FILLCELL_X1 FILLER_8_232 ();
 FILLCELL_X4 FILLER_8_240 ();
 FILLCELL_X4 FILLER_8_251 ();
 FILLCELL_X8 FILLER_8_272 ();
 FILLCELL_X2 FILLER_8_280 ();
 FILLCELL_X1 FILLER_8_282 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_16 ();
 FILLCELL_X1 FILLER_9_18 ();
 FILLCELL_X2 FILLER_9_26 ();
 FILLCELL_X1 FILLER_9_28 ();
 FILLCELL_X2 FILLER_9_60 ();
 FILLCELL_X1 FILLER_9_62 ();
 FILLCELL_X2 FILLER_9_77 ();
 FILLCELL_X4 FILLER_9_96 ();
 FILLCELL_X2 FILLER_9_100 ();
 FILLCELL_X1 FILLER_9_102 ();
 FILLCELL_X32 FILLER_9_108 ();
 FILLCELL_X16 FILLER_9_140 ();
 FILLCELL_X8 FILLER_9_156 ();
 FILLCELL_X4 FILLER_9_164 ();
 FILLCELL_X2 FILLER_9_168 ();
 FILLCELL_X4 FILLER_9_183 ();
 FILLCELL_X1 FILLER_9_187 ();
 FILLCELL_X16 FILLER_9_195 ();
 FILLCELL_X4 FILLER_9_211 ();
 FILLCELL_X4 FILLER_9_239 ();
 FILLCELL_X8 FILLER_9_248 ();
 FILLCELL_X8 FILLER_9_270 ();
 FILLCELL_X4 FILLER_9_278 ();
 FILLCELL_X1 FILLER_9_282 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_27 ();
 FILLCELL_X1 FILLER_10_29 ();
 FILLCELL_X8 FILLER_10_47 ();
 FILLCELL_X4 FILLER_10_55 ();
 FILLCELL_X2 FILLER_10_59 ();
 FILLCELL_X16 FILLER_10_78 ();
 FILLCELL_X8 FILLER_10_94 ();
 FILLCELL_X1 FILLER_10_102 ();
 FILLCELL_X1 FILLER_10_163 ();
 FILLCELL_X2 FILLER_10_181 ();
 FILLCELL_X2 FILLER_10_190 ();
 FILLCELL_X2 FILLER_10_199 ();
 FILLCELL_X1 FILLER_10_201 ();
 FILLCELL_X4 FILLER_10_209 ();
 FILLCELL_X1 FILLER_10_213 ();
 FILLCELL_X4 FILLER_10_221 ();
 FILLCELL_X1 FILLER_10_225 ();
 FILLCELL_X4 FILLER_10_233 ();
 FILLCELL_X1 FILLER_10_247 ();
 FILLCELL_X8 FILLER_10_269 ();
 FILLCELL_X4 FILLER_10_277 ();
 FILLCELL_X2 FILLER_10_281 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_33 ();
 FILLCELL_X1 FILLER_11_35 ();
 FILLCELL_X32 FILLER_11_49 ();
 FILLCELL_X8 FILLER_11_122 ();
 FILLCELL_X2 FILLER_11_130 ();
 FILLCELL_X1 FILLER_11_132 ();
 FILLCELL_X4 FILLER_11_140 ();
 FILLCELL_X1 FILLER_11_144 ();
 FILLCELL_X1 FILLER_11_189 ();
 FILLCELL_X2 FILLER_11_197 ();
 FILLCELL_X1 FILLER_11_199 ();
 FILLCELL_X8 FILLER_11_224 ();
 FILLCELL_X2 FILLER_11_232 ();
 FILLCELL_X1 FILLER_11_234 ();
 FILLCELL_X4 FILLER_11_259 ();
 FILLCELL_X2 FILLER_11_263 ();
 FILLCELL_X1 FILLER_11_265 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_5 ();
 FILLCELL_X2 FILLER_12_9 ();
 FILLCELL_X1 FILLER_12_11 ();
 FILLCELL_X1 FILLER_12_49 ();
 FILLCELL_X8 FILLER_12_74 ();
 FILLCELL_X4 FILLER_12_82 ();
 FILLCELL_X2 FILLER_12_93 ();
 FILLCELL_X1 FILLER_12_95 ();
 FILLCELL_X1 FILLER_12_115 ();
 FILLCELL_X1 FILLER_12_147 ();
 FILLCELL_X2 FILLER_12_155 ();
 FILLCELL_X1 FILLER_12_157 ();
 FILLCELL_X2 FILLER_12_165 ();
 FILLCELL_X4 FILLER_12_174 ();
 FILLCELL_X4 FILLER_12_185 ();
 FILLCELL_X4 FILLER_12_206 ();
 FILLCELL_X16 FILLER_12_226 ();
 FILLCELL_X4 FILLER_12_242 ();
 FILLCELL_X2 FILLER_12_246 ();
 FILLCELL_X1 FILLER_12_248 ();
 FILLCELL_X2 FILLER_12_266 ();
 FILLCELL_X1 FILLER_12_268 ();
 FILLCELL_X8 FILLER_12_272 ();
 FILLCELL_X2 FILLER_12_280 ();
 FILLCELL_X1 FILLER_12_282 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_9 ();
 FILLCELL_X1 FILLER_13_13 ();
 FILLCELL_X2 FILLER_13_31 ();
 FILLCELL_X1 FILLER_13_33 ();
 FILLCELL_X8 FILLER_13_41 ();
 FILLCELL_X4 FILLER_13_49 ();
 FILLCELL_X2 FILLER_13_53 ();
 FILLCELL_X1 FILLER_13_55 ();
 FILLCELL_X2 FILLER_13_63 ();
 FILLCELL_X1 FILLER_13_65 ();
 FILLCELL_X8 FILLER_13_73 ();
 FILLCELL_X4 FILLER_13_81 ();
 FILLCELL_X8 FILLER_13_92 ();
 FILLCELL_X32 FILLER_13_114 ();
 FILLCELL_X32 FILLER_13_146 ();
 FILLCELL_X16 FILLER_13_178 ();
 FILLCELL_X8 FILLER_13_194 ();
 FILLCELL_X4 FILLER_13_202 ();
 FILLCELL_X2 FILLER_13_206 ();
 FILLCELL_X1 FILLER_13_208 ();
 FILLCELL_X4 FILLER_13_226 ();
 FILLCELL_X8 FILLER_13_271 ();
 FILLCELL_X4 FILLER_13_279 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_5 ();
 FILLCELL_X4 FILLER_14_30 ();
 FILLCELL_X2 FILLER_14_34 ();
 FILLCELL_X2 FILLER_14_53 ();
 FILLCELL_X4 FILLER_14_72 ();
 FILLCELL_X1 FILLER_14_76 ();
 FILLCELL_X4 FILLER_14_105 ();
 FILLCELL_X16 FILLER_14_127 ();
 FILLCELL_X1 FILLER_14_143 ();
 FILLCELL_X2 FILLER_14_161 ();
 FILLCELL_X1 FILLER_14_163 ();
 FILLCELL_X2 FILLER_14_171 ();
 FILLCELL_X1 FILLER_14_173 ();
 FILLCELL_X16 FILLER_14_191 ();
 FILLCELL_X4 FILLER_14_207 ();
 FILLCELL_X4 FILLER_14_218 ();
 FILLCELL_X2 FILLER_14_229 ();
 FILLCELL_X2 FILLER_14_238 ();
 FILLCELL_X1 FILLER_14_240 ();
 FILLCELL_X2 FILLER_14_248 ();
 FILLCELL_X1 FILLER_14_250 ();
 FILLCELL_X2 FILLER_14_258 ();
 FILLCELL_X16 FILLER_14_267 ();
 FILLCELL_X1 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_19 ();
 FILLCELL_X1 FILLER_15_28 ();
 FILLCELL_X4 FILLER_15_43 ();
 FILLCELL_X2 FILLER_15_47 ();
 FILLCELL_X32 FILLER_15_70 ();
 FILLCELL_X2 FILLER_15_102 ();
 FILLCELL_X1 FILLER_15_104 ();
 FILLCELL_X8 FILLER_15_122 ();
 FILLCELL_X1 FILLER_15_130 ();
 FILLCELL_X2 FILLER_15_138 ();
 FILLCELL_X4 FILLER_15_164 ();
 FILLCELL_X1 FILLER_15_168 ();
 FILLCELL_X32 FILLER_15_183 ();
 FILLCELL_X16 FILLER_15_215 ();
 FILLCELL_X1 FILLER_15_231 ();
 FILLCELL_X8 FILLER_15_273 ();
 FILLCELL_X2 FILLER_15_281 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X1 FILLER_16_49 ();
 FILLCELL_X4 FILLER_16_67 ();
 FILLCELL_X2 FILLER_16_71 ();
 FILLCELL_X1 FILLER_16_73 ();
 FILLCELL_X4 FILLER_16_98 ();
 FILLCELL_X2 FILLER_16_102 ();
 FILLCELL_X8 FILLER_16_138 ();
 FILLCELL_X4 FILLER_16_146 ();
 FILLCELL_X2 FILLER_16_150 ();
 FILLCELL_X2 FILLER_16_173 ();
 FILLCELL_X1 FILLER_16_175 ();
 FILLCELL_X8 FILLER_16_202 ();
 FILLCELL_X2 FILLER_16_210 ();
 FILLCELL_X32 FILLER_16_231 ();
 FILLCELL_X8 FILLER_16_263 ();
 FILLCELL_X8 FILLER_16_274 ();
 FILLCELL_X1 FILLER_16_282 ();
 FILLCELL_X32 FILLER_17_4 ();
 FILLCELL_X32 FILLER_17_36 ();
 FILLCELL_X16 FILLER_17_68 ();
 FILLCELL_X4 FILLER_17_84 ();
 FILLCELL_X2 FILLER_17_88 ();
 FILLCELL_X1 FILLER_17_90 ();
 FILLCELL_X16 FILLER_17_98 ();
 FILLCELL_X8 FILLER_17_114 ();
 FILLCELL_X2 FILLER_17_122 ();
 FILLCELL_X16 FILLER_17_145 ();
 FILLCELL_X2 FILLER_17_161 ();
 FILLCELL_X1 FILLER_17_163 ();
 FILLCELL_X8 FILLER_17_171 ();
 FILLCELL_X2 FILLER_17_210 ();
 FILLCELL_X32 FILLER_17_226 ();
 FILLCELL_X4 FILLER_17_258 ();
 FILLCELL_X8 FILLER_17_269 ();
 FILLCELL_X4 FILLER_17_277 ();
 FILLCELL_X2 FILLER_17_281 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_9 ();
 FILLCELL_X1 FILLER_18_13 ();
 FILLCELL_X4 FILLER_18_31 ();
 FILLCELL_X2 FILLER_18_35 ();
 FILLCELL_X4 FILLER_18_85 ();
 FILLCELL_X1 FILLER_18_89 ();
 FILLCELL_X4 FILLER_18_111 ();
 FILLCELL_X8 FILLER_18_139 ();
 FILLCELL_X1 FILLER_18_147 ();
 FILLCELL_X4 FILLER_18_155 ();
 FILLCELL_X16 FILLER_18_166 ();
 FILLCELL_X8 FILLER_18_182 ();
 FILLCELL_X4 FILLER_18_197 ();
 FILLCELL_X4 FILLER_18_208 ();
 FILLCELL_X1 FILLER_18_229 ();
 FILLCELL_X2 FILLER_18_244 ();
 FILLCELL_X2 FILLER_18_280 ();
 FILLCELL_X1 FILLER_18_282 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X4 FILLER_19_20 ();
 FILLCELL_X2 FILLER_19_24 ();
 FILLCELL_X1 FILLER_19_26 ();
 FILLCELL_X2 FILLER_19_65 ();
 FILLCELL_X2 FILLER_19_91 ();
 FILLCELL_X16 FILLER_19_110 ();
 FILLCELL_X8 FILLER_19_126 ();
 FILLCELL_X2 FILLER_19_134 ();
 FILLCELL_X4 FILLER_19_158 ();
 FILLCELL_X2 FILLER_19_162 ();
 FILLCELL_X1 FILLER_19_219 ();
 FILLCELL_X4 FILLER_19_244 ();
 FILLCELL_X2 FILLER_19_255 ();
 FILLCELL_X8 FILLER_19_271 ();
 FILLCELL_X4 FILLER_19_279 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_17 ();
 FILLCELL_X2 FILLER_20_21 ();
 FILLCELL_X2 FILLER_20_47 ();
 FILLCELL_X1 FILLER_20_49 ();
 FILLCELL_X4 FILLER_20_57 ();
 FILLCELL_X2 FILLER_20_61 ();
 FILLCELL_X1 FILLER_20_63 ();
 FILLCELL_X4 FILLER_20_69 ();
 FILLCELL_X2 FILLER_20_73 ();
 FILLCELL_X4 FILLER_20_82 ();
 FILLCELL_X2 FILLER_20_86 ();
 FILLCELL_X1 FILLER_20_88 ();
 FILLCELL_X16 FILLER_20_110 ();
 FILLCELL_X4 FILLER_20_126 ();
 FILLCELL_X1 FILLER_20_147 ();
 FILLCELL_X1 FILLER_20_155 ();
 FILLCELL_X8 FILLER_20_177 ();
 FILLCELL_X1 FILLER_20_185 ();
 FILLCELL_X8 FILLER_20_210 ();
 FILLCELL_X4 FILLER_20_218 ();
 FILLCELL_X2 FILLER_20_222 ();
 FILLCELL_X1 FILLER_20_224 ();
 FILLCELL_X8 FILLER_20_232 ();
 FILLCELL_X4 FILLER_20_240 ();
 FILLCELL_X2 FILLER_20_244 ();
 FILLCELL_X4 FILLER_20_277 ();
 FILLCELL_X2 FILLER_20_281 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_9 ();
 FILLCELL_X1 FILLER_21_13 ();
 FILLCELL_X16 FILLER_21_31 ();
 FILLCELL_X16 FILLER_21_59 ();
 FILLCELL_X8 FILLER_21_75 ();
 FILLCELL_X1 FILLER_21_83 ();
 FILLCELL_X2 FILLER_21_88 ();
 FILLCELL_X32 FILLER_21_104 ();
 FILLCELL_X2 FILLER_21_136 ();
 FILLCELL_X16 FILLER_21_145 ();
 FILLCELL_X1 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_186 ();
 FILLCELL_X16 FILLER_21_197 ();
 FILLCELL_X1 FILLER_21_213 ();
 FILLCELL_X2 FILLER_21_221 ();
 FILLCELL_X16 FILLER_21_230 ();
 FILLCELL_X4 FILLER_21_246 ();
 FILLCELL_X1 FILLER_21_250 ();
 FILLCELL_X8 FILLER_21_268 ();
 FILLCELL_X4 FILLER_21_276 ();
 FILLCELL_X2 FILLER_21_280 ();
 FILLCELL_X1 FILLER_21_282 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_5 ();
 FILLCELL_X2 FILLER_22_9 ();
 FILLCELL_X1 FILLER_22_35 ();
 FILLCELL_X2 FILLER_22_53 ();
 FILLCELL_X2 FILLER_22_62 ();
 FILLCELL_X1 FILLER_22_64 ();
 FILLCELL_X1 FILLER_22_99 ();
 FILLCELL_X2 FILLER_22_107 ();
 FILLCELL_X8 FILLER_22_150 ();
 FILLCELL_X2 FILLER_22_158 ();
 FILLCELL_X1 FILLER_22_160 ();
 FILLCELL_X8 FILLER_22_175 ();
 FILLCELL_X4 FILLER_22_183 ();
 FILLCELL_X4 FILLER_22_197 ();
 FILLCELL_X2 FILLER_22_201 ();
 FILLCELL_X1 FILLER_22_227 ();
 FILLCELL_X1 FILLER_22_249 ();
 FILLCELL_X8 FILLER_22_274 ();
 FILLCELL_X1 FILLER_22_282 ();
 FILLCELL_X8 FILLER_23_5 ();
 FILLCELL_X2 FILLER_23_13 ();
 FILLCELL_X4 FILLER_23_29 ();
 FILLCELL_X2 FILLER_23_33 ();
 FILLCELL_X4 FILLER_23_52 ();
 FILLCELL_X1 FILLER_23_56 ();
 FILLCELL_X1 FILLER_23_88 ();
 FILLCELL_X4 FILLER_23_103 ();
 FILLCELL_X2 FILLER_23_107 ();
 FILLCELL_X16 FILLER_23_155 ();
 FILLCELL_X8 FILLER_23_171 ();
 FILLCELL_X4 FILLER_23_179 ();
 FILLCELL_X16 FILLER_23_190 ();
 FILLCELL_X4 FILLER_23_206 ();
 FILLCELL_X4 FILLER_23_217 ();
 FILLCELL_X2 FILLER_23_221 ();
 FILLCELL_X1 FILLER_23_230 ();
 FILLCELL_X16 FILLER_23_256 ();
 FILLCELL_X8 FILLER_23_272 ();
 FILLCELL_X2 FILLER_23_280 ();
 FILLCELL_X1 FILLER_23_282 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X4 FILLER_24_33 ();
 FILLCELL_X8 FILLER_24_64 ();
 FILLCELL_X4 FILLER_24_72 ();
 FILLCELL_X16 FILLER_24_126 ();
 FILLCELL_X4 FILLER_24_149 ();
 FILLCELL_X4 FILLER_24_160 ();
 FILLCELL_X2 FILLER_24_164 ();
 FILLCELL_X2 FILLER_24_207 ();
 FILLCELL_X1 FILLER_24_209 ();
 FILLCELL_X2 FILLER_24_227 ();
 FILLCELL_X4 FILLER_24_231 ();
 FILLCELL_X1 FILLER_24_235 ();
 FILLCELL_X16 FILLER_24_260 ();
 FILLCELL_X4 FILLER_24_276 ();
 FILLCELL_X2 FILLER_24_280 ();
 FILLCELL_X1 FILLER_24_282 ();
 FILLCELL_X16 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_17 ();
 FILLCELL_X16 FILLER_25_52 ();
 FILLCELL_X4 FILLER_25_68 ();
 FILLCELL_X2 FILLER_25_72 ();
 FILLCELL_X1 FILLER_25_74 ();
 FILLCELL_X8 FILLER_25_88 ();
 FILLCELL_X1 FILLER_25_96 ();
 FILLCELL_X4 FILLER_25_114 ();
 FILLCELL_X2 FILLER_25_118 ();
 FILLCELL_X16 FILLER_25_124 ();
 FILLCELL_X16 FILLER_25_153 ();
 FILLCELL_X4 FILLER_25_169 ();
 FILLCELL_X2 FILLER_25_173 ();
 FILLCELL_X4 FILLER_25_204 ();
 FILLCELL_X2 FILLER_26_1 ();
 FILLCELL_X1 FILLER_26_41 ();
 FILLCELL_X4 FILLER_26_63 ();
 FILLCELL_X4 FILLER_26_87 ();
 FILLCELL_X2 FILLER_26_91 ();
 FILLCELL_X1 FILLER_26_93 ();
 FILLCELL_X8 FILLER_26_101 ();
 FILLCELL_X4 FILLER_26_109 ();
 FILLCELL_X2 FILLER_26_113 ();
 FILLCELL_X1 FILLER_26_115 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X8 FILLER_26_161 ();
 FILLCELL_X2 FILLER_26_169 ();
 FILLCELL_X8 FILLER_26_223 ();
 FILLCELL_X4 FILLER_26_231 ();
 FILLCELL_X16 FILLER_26_240 ();
 FILLCELL_X1 FILLER_26_256 ();
 FILLCELL_X16 FILLER_26_264 ();
 FILLCELL_X2 FILLER_26_280 ();
 FILLCELL_X1 FILLER_26_282 ();
 FILLCELL_X2 FILLER_27_1 ();
 FILLCELL_X8 FILLER_27_20 ();
 FILLCELL_X4 FILLER_27_28 ();
 FILLCELL_X2 FILLER_27_32 ();
 FILLCELL_X1 FILLER_27_34 ();
 FILLCELL_X16 FILLER_27_52 ();
 FILLCELL_X8 FILLER_27_68 ();
 FILLCELL_X4 FILLER_27_76 ();
 FILLCELL_X1 FILLER_27_80 ();
 FILLCELL_X16 FILLER_27_87 ();
 FILLCELL_X4 FILLER_27_103 ();
 FILLCELL_X1 FILLER_27_107 ();
 FILLCELL_X4 FILLER_27_120 ();
 FILLCELL_X32 FILLER_27_137 ();
 FILLCELL_X4 FILLER_27_169 ();
 FILLCELL_X32 FILLER_27_190 ();
 FILLCELL_X8 FILLER_27_229 ();
 FILLCELL_X2 FILLER_27_237 ();
 FILLCELL_X16 FILLER_27_263 ();
 FILLCELL_X4 FILLER_27_279 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X4 FILLER_28_65 ();
 FILLCELL_X1 FILLER_28_69 ();
 FILLCELL_X8 FILLER_28_99 ();
 FILLCELL_X2 FILLER_28_107 ();
 FILLCELL_X1 FILLER_28_121 ();
 FILLCELL_X8 FILLER_28_134 ();
 FILLCELL_X4 FILLER_28_142 ();
 FILLCELL_X4 FILLER_28_164 ();
 FILLCELL_X2 FILLER_28_189 ();
 FILLCELL_X1 FILLER_28_191 ();
 FILLCELL_X8 FILLER_28_201 ();
 FILLCELL_X1 FILLER_28_209 ();
 FILLCELL_X2 FILLER_28_217 ();
 FILLCELL_X8 FILLER_28_236 ();
 FILLCELL_X2 FILLER_28_244 ();
 FILLCELL_X2 FILLER_28_253 ();
 FILLCELL_X1 FILLER_28_255 ();
 FILLCELL_X2 FILLER_28_263 ();
 FILLCELL_X1 FILLER_28_282 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_9 ();
 FILLCELL_X16 FILLER_29_29 ();
 FILLCELL_X8 FILLER_29_45 ();
 FILLCELL_X4 FILLER_29_53 ();
 FILLCELL_X1 FILLER_29_57 ();
 FILLCELL_X1 FILLER_29_71 ();
 FILLCELL_X8 FILLER_29_78 ();
 FILLCELL_X16 FILLER_29_91 ();
 FILLCELL_X1 FILLER_29_119 ();
 FILLCELL_X2 FILLER_29_125 ();
 FILLCELL_X1 FILLER_29_127 ();
 FILLCELL_X4 FILLER_29_135 ();
 FILLCELL_X2 FILLER_29_139 ();
 FILLCELL_X1 FILLER_29_141 ();
 FILLCELL_X16 FILLER_29_162 ();
 FILLCELL_X1 FILLER_29_208 ();
 FILLCELL_X16 FILLER_29_264 ();
 FILLCELL_X2 FILLER_29_280 ();
 FILLCELL_X1 FILLER_29_282 ();
 FILLCELL_X4 FILLER_30_4 ();
 FILLCELL_X2 FILLER_30_8 ();
 FILLCELL_X2 FILLER_30_24 ();
 FILLCELL_X1 FILLER_30_26 ();
 FILLCELL_X4 FILLER_30_37 ();
 FILLCELL_X1 FILLER_30_41 ();
 FILLCELL_X32 FILLER_30_61 ();
 FILLCELL_X32 FILLER_30_93 ();
 FILLCELL_X8 FILLER_30_125 ();
 FILLCELL_X4 FILLER_30_133 ();
 FILLCELL_X2 FILLER_30_137 ();
 FILLCELL_X1 FILLER_30_139 ();
 FILLCELL_X8 FILLER_30_170 ();
 FILLCELL_X2 FILLER_30_178 ();
 FILLCELL_X1 FILLER_30_191 ();
 FILLCELL_X4 FILLER_30_203 ();
 FILLCELL_X8 FILLER_30_212 ();
 FILLCELL_X32 FILLER_30_251 ();
 FILLCELL_X1 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_30 ();
 FILLCELL_X2 FILLER_31_38 ();
 FILLCELL_X2 FILLER_31_53 ();
 FILLCELL_X16 FILLER_31_57 ();
 FILLCELL_X4 FILLER_31_73 ();
 FILLCELL_X2 FILLER_31_77 ();
 FILLCELL_X1 FILLER_31_79 ();
 FILLCELL_X1 FILLER_31_84 ();
 FILLCELL_X1 FILLER_31_90 ();
 FILLCELL_X32 FILLER_31_99 ();
 FILLCELL_X16 FILLER_31_131 ();
 FILLCELL_X1 FILLER_31_147 ();
 FILLCELL_X2 FILLER_31_186 ();
 FILLCELL_X4 FILLER_31_191 ();
 FILLCELL_X2 FILLER_31_195 ();
 FILLCELL_X1 FILLER_31_197 ();
 FILLCELL_X1 FILLER_31_209 ();
 FILLCELL_X32 FILLER_31_214 ();
 FILLCELL_X32 FILLER_31_246 ();
 FILLCELL_X4 FILLER_31_278 ();
 FILLCELL_X1 FILLER_31_282 ();
 FILLCELL_X1 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_6 ();
 FILLCELL_X2 FILLER_32_13 ();
 FILLCELL_X1 FILLER_32_19 ();
 FILLCELL_X4 FILLER_32_36 ();
 FILLCELL_X16 FILLER_32_62 ();
 FILLCELL_X4 FILLER_32_78 ();
 FILLCELL_X1 FILLER_32_96 ();
 FILLCELL_X2 FILLER_32_105 ();
 FILLCELL_X2 FILLER_32_110 ();
 FILLCELL_X1 FILLER_32_112 ();
 FILLCELL_X2 FILLER_32_117 ();
 FILLCELL_X8 FILLER_32_123 ();
 FILLCELL_X4 FILLER_32_131 ();
 FILLCELL_X1 FILLER_32_135 ();
 FILLCELL_X1 FILLER_32_140 ();
 FILLCELL_X32 FILLER_32_151 ();
 FILLCELL_X2 FILLER_32_183 ();
 FILLCELL_X1 FILLER_32_185 ();
 FILLCELL_X32 FILLER_32_221 ();
 FILLCELL_X16 FILLER_32_253 ();
 FILLCELL_X8 FILLER_32_269 ();
 FILLCELL_X4 FILLER_32_277 ();
 FILLCELL_X2 FILLER_32_281 ();
 FILLCELL_X4 FILLER_33_21 ();
 FILLCELL_X2 FILLER_33_45 ();
 FILLCELL_X1 FILLER_33_47 ();
 FILLCELL_X16 FILLER_33_58 ();
 FILLCELL_X1 FILLER_33_107 ();
 FILLCELL_X1 FILLER_33_115 ();
 FILLCELL_X2 FILLER_33_120 ();
 FILLCELL_X4 FILLER_33_128 ();
 FILLCELL_X2 FILLER_33_154 ();
 FILLCELL_X4 FILLER_33_158 ();
 FILLCELL_X16 FILLER_33_179 ();
 FILLCELL_X4 FILLER_33_195 ();
 FILLCELL_X2 FILLER_33_199 ();
 FILLCELL_X8 FILLER_33_204 ();
 FILLCELL_X32 FILLER_33_231 ();
 FILLCELL_X16 FILLER_33_263 ();
 FILLCELL_X4 FILLER_33_279 ();
 FILLCELL_X8 FILLER_34_34 ();
 FILLCELL_X4 FILLER_34_42 ();
 FILLCELL_X1 FILLER_34_46 ();
 FILLCELL_X4 FILLER_34_91 ();
 FILLCELL_X4 FILLER_34_99 ();
 FILLCELL_X2 FILLER_34_103 ();
 FILLCELL_X8 FILLER_34_109 ();
 FILLCELL_X1 FILLER_34_117 ();
 FILLCELL_X4 FILLER_34_135 ();
 FILLCELL_X1 FILLER_34_139 ();
 FILLCELL_X2 FILLER_34_166 ();
 FILLCELL_X2 FILLER_34_176 ();
 FILLCELL_X4 FILLER_34_195 ();
 FILLCELL_X2 FILLER_34_199 ();
 FILLCELL_X1 FILLER_34_201 ();
 FILLCELL_X32 FILLER_34_240 ();
 FILLCELL_X8 FILLER_34_272 ();
 FILLCELL_X2 FILLER_34_280 ();
 FILLCELL_X1 FILLER_34_282 ();
 FILLCELL_X1 FILLER_35_11 ();
 FILLCELL_X2 FILLER_35_16 ();
 FILLCELL_X16 FILLER_35_39 ();
 FILLCELL_X8 FILLER_35_55 ();
 FILLCELL_X4 FILLER_35_63 ();
 FILLCELL_X2 FILLER_35_67 ();
 FILLCELL_X1 FILLER_35_69 ();
 FILLCELL_X1 FILLER_35_116 ();
 FILLCELL_X8 FILLER_35_131 ();
 FILLCELL_X2 FILLER_35_139 ();
 FILLCELL_X1 FILLER_35_141 ();
 FILLCELL_X4 FILLER_35_168 ();
 FILLCELL_X1 FILLER_35_178 ();
 FILLCELL_X4 FILLER_35_189 ();
 FILLCELL_X2 FILLER_35_193 ();
 FILLCELL_X1 FILLER_35_199 ();
 FILLCELL_X1 FILLER_35_227 ();
 FILLCELL_X32 FILLER_35_237 ();
 FILLCELL_X8 FILLER_35_269 ();
 FILLCELL_X4 FILLER_35_277 ();
 FILLCELL_X2 FILLER_35_281 ();
 FILLCELL_X8 FILLER_36_1 ();
 FILLCELL_X2 FILLER_36_9 ();
 FILLCELL_X1 FILLER_36_11 ();
 FILLCELL_X8 FILLER_36_35 ();
 FILLCELL_X4 FILLER_36_43 ();
 FILLCELL_X2 FILLER_36_47 ();
 FILLCELL_X1 FILLER_36_49 ();
 FILLCELL_X16 FILLER_36_53 ();
 FILLCELL_X8 FILLER_36_69 ();
 FILLCELL_X4 FILLER_36_77 ();
 FILLCELL_X1 FILLER_36_81 ();
 FILLCELL_X1 FILLER_36_102 ();
 FILLCELL_X1 FILLER_36_110 ();
 FILLCELL_X16 FILLER_36_128 ();
 FILLCELL_X4 FILLER_36_144 ();
 FILLCELL_X8 FILLER_36_191 ();
 FILLCELL_X2 FILLER_36_199 ();
 FILLCELL_X1 FILLER_36_201 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X16 FILLER_36_257 ();
 FILLCELL_X8 FILLER_36_273 ();
 FILLCELL_X2 FILLER_36_281 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X8 FILLER_37_65 ();
 FILLCELL_X4 FILLER_37_73 ();
 FILLCELL_X32 FILLER_37_90 ();
 FILLCELL_X16 FILLER_37_122 ();
 FILLCELL_X8 FILLER_37_138 ();
 FILLCELL_X2 FILLER_37_146 ();
 FILLCELL_X2 FILLER_37_167 ();
 FILLCELL_X16 FILLER_37_172 ();
 FILLCELL_X1 FILLER_37_188 ();
 FILLCELL_X2 FILLER_37_195 ();
 FILLCELL_X1 FILLER_37_197 ();
 FILLCELL_X4 FILLER_37_201 ();
 FILLCELL_X1 FILLER_37_210 ();
 FILLCELL_X2 FILLER_37_214 ();
 FILLCELL_X32 FILLER_37_219 ();
 FILLCELL_X32 FILLER_37_251 ();
endmodule
